* NGSPICE file created from BundleParser.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

.subckt BundleParser vdd gnd clock_i enable_i bundle_i[127] bundle_i[126] bundle_i[125]
+ bundle_i[124] bundle_i[123] bundle_i[122] bundle_i[121] bundle_i[120] bundle_i[119]
+ bundle_i[118] bundle_i[117] bundle_i[116] bundle_i[115] bundle_i[114] bundle_i[113]
+ bundle_i[112] bundle_i[111] bundle_i[110] bundle_i[109] bundle_i[108] bundle_i[107]
+ bundle_i[106] bundle_i[105] bundle_i[104] bundle_i[103] bundle_i[102] bundle_i[101]
+ bundle_i[100] bundle_i[99] bundle_i[98] bundle_i[97] bundle_i[96] bundle_i[95] bundle_i[94]
+ bundle_i[93] bundle_i[92] bundle_i[91] bundle_i[90] bundle_i[89] bundle_i[88] bundle_i[87]
+ bundle_i[86] bundle_i[85] bundle_i[84] bundle_i[83] bundle_i[82] bundle_i[81] bundle_i[80]
+ bundle_i[79] bundle_i[78] bundle_i[77] bundle_i[76] bundle_i[75] bundle_i[74] bundle_i[73]
+ bundle_i[72] bundle_i[71] bundle_i[70] bundle_i[69] bundle_i[68] bundle_i[67] bundle_i[66]
+ bundle_i[65] bundle_i[64] bundle_i[63] bundle_i[62] bundle_i[61] bundle_i[60] bundle_i[59]
+ bundle_i[58] bundle_i[57] bundle_i[56] bundle_i[55] bundle_i[54] bundle_i[53] bundle_i[52]
+ bundle_i[51] bundle_i[50] bundle_i[49] bundle_i[48] bundle_i[47] bundle_i[46] bundle_i[45]
+ bundle_i[44] bundle_i[43] bundle_i[42] bundle_i[41] bundle_i[40] bundle_i[39] bundle_i[38]
+ bundle_i[37] bundle_i[36] bundle_i[35] bundle_i[34] bundle_i[33] bundle_i[32] bundle_i[31]
+ bundle_i[30] bundle_i[29] bundle_i[28] bundle_i[27] bundle_i[26] bundle_i[25] bundle_i[24]
+ bundle_i[23] bundle_i[22] bundle_i[21] bundle_i[20] bundle_i[19] bundle_i[18] bundle_i[17]
+ bundle_i[16] bundle_i[15] bundle_i[14] bundle_i[13] bundle_i[12] bundle_i[11] bundle_i[10]
+ bundle_i[9] bundle_i[8] bundle_i[7] bundle_i[6] bundle_i[5] bundle_i[4] bundle_i[3]
+ bundle_i[2] bundle_i[1] bundle_i[0] bundleAddress_i[63] bundleAddress_i[62] bundleAddress_i[61]
+ bundleAddress_i[60] bundleAddress_i[59] bundleAddress_i[58] bundleAddress_i[57]
+ bundleAddress_i[56] bundleAddress_i[55] bundleAddress_i[54] bundleAddress_i[53]
+ bundleAddress_i[52] bundleAddress_i[51] bundleAddress_i[50] bundleAddress_i[49]
+ bundleAddress_i[48] bundleAddress_i[47] bundleAddress_i[46] bundleAddress_i[45]
+ bundleAddress_i[44] bundleAddress_i[43] bundleAddress_i[42] bundleAddress_i[41]
+ bundleAddress_i[40] bundleAddress_i[39] bundleAddress_i[38] bundleAddress_i[37]
+ bundleAddress_i[36] bundleAddress_i[35] bundleAddress_i[34] bundleAddress_i[33]
+ bundleAddress_i[32] bundleAddress_i[31] bundleAddress_i[30] bundleAddress_i[29]
+ bundleAddress_i[28] bundleAddress_i[27] bundleAddress_i[26] bundleAddress_i[25]
+ bundleAddress_i[24] bundleAddress_i[23] bundleAddress_i[22] bundleAddress_i[21]
+ bundleAddress_i[20] bundleAddress_i[19] bundleAddress_i[18] bundleAddress_i[17]
+ bundleAddress_i[16] bundleAddress_i[15] bundleAddress_i[14] bundleAddress_i[13]
+ bundleAddress_i[12] bundleAddress_i[11] bundleAddress_i[10] bundleAddress_i[9] bundleAddress_i[8]
+ bundleAddress_i[7] bundleAddress_i[6] bundleAddress_i[5] bundleAddress_i[4] bundleAddress_i[3]
+ bundleAddress_i[2] bundleAddress_i[1] bundleAddress_i[0] bundleLen_i[1] bundleLen_i[0]
+ is64Bit_i bundlePid_i[31] bundlePid_i[30] bundlePid_i[29] bundlePid_i[28] bundlePid_i[27]
+ bundlePid_i[26] bundlePid_i[25] bundlePid_i[24] bundlePid_i[23] bundlePid_i[22]
+ bundlePid_i[21] bundlePid_i[20] bundlePid_i[19] bundlePid_i[18] bundlePid_i[17]
+ bundlePid_i[16] bundlePid_i[15] bundlePid_i[14] bundlePid_i[13] bundlePid_i[12]
+ bundlePid_i[11] bundlePid_i[10] bundlePid_i[9] bundlePid_i[8] bundlePid_i[7] bundlePid_i[6]
+ bundlePid_i[5] bundlePid_i[4] bundlePid_i[3] bundlePid_i[2] bundlePid_i[1] bundlePid_i[0]
+ bundleTid_i[63] bundleTid_i[62] bundleTid_i[61] bundleTid_i[60] bundleTid_i[59]
+ bundleTid_i[58] bundleTid_i[57] bundleTid_i[56] bundleTid_i[55] bundleTid_i[54]
+ bundleTid_i[53] bundleTid_i[52] bundleTid_i[51] bundleTid_i[50] bundleTid_i[49]
+ bundleTid_i[48] bundleTid_i[47] bundleTid_i[46] bundleTid_i[45] bundleTid_i[44]
+ bundleTid_i[43] bundleTid_i[42] bundleTid_i[41] bundleTid_i[40] bundleTid_i[39]
+ bundleTid_i[38] bundleTid_i[37] bundleTid_i[36] bundleTid_i[35] bundleTid_i[34]
+ bundleTid_i[33] bundleTid_i[32] bundleTid_i[31] bundleTid_i[30] bundleTid_i[29]
+ bundleTid_i[28] bundleTid_i[27] bundleTid_i[26] bundleTid_i[25] bundleTid_i[24]
+ bundleTid_i[23] bundleTid_i[22] bundleTid_i[21] bundleTid_i[20] bundleTid_i[19]
+ bundleTid_i[18] bundleTid_i[17] bundleTid_i[16] bundleTid_i[15] bundleTid_i[14]
+ bundleTid_i[13] bundleTid_i[12] bundleTid_i[11] bundleTid_i[10] bundleTid_i[9] bundleTid_i[8]
+ bundleTid_i[7] bundleTid_i[6] bundleTid_i[5] bundleTid_i[4] bundleTid_i[3] bundleTid_i[2]
+ bundleTid_i[1] bundleTid_i[0] bundleStartMajId_i[63] bundleStartMajId_i[62] bundleStartMajId_i[61]
+ bundleStartMajId_i[60] bundleStartMajId_i[59] bundleStartMajId_i[58] bundleStartMajId_i[57]
+ bundleStartMajId_i[56] bundleStartMajId_i[55] bundleStartMajId_i[54] bundleStartMajId_i[53]
+ bundleStartMajId_i[52] bundleStartMajId_i[51] bundleStartMajId_i[50] bundleStartMajId_i[49]
+ bundleStartMajId_i[48] bundleStartMajId_i[47] bundleStartMajId_i[46] bundleStartMajId_i[45]
+ bundleStartMajId_i[44] bundleStartMajId_i[43] bundleStartMajId_i[42] bundleStartMajId_i[41]
+ bundleStartMajId_i[40] bundleStartMajId_i[39] bundleStartMajId_i[38] bundleStartMajId_i[37]
+ bundleStartMajId_i[36] bundleStartMajId_i[35] bundleStartMajId_i[34] bundleStartMajId_i[33]
+ bundleStartMajId_i[32] bundleStartMajId_i[31] bundleStartMajId_i[30] bundleStartMajId_i[29]
+ bundleStartMajId_i[28] bundleStartMajId_i[27] bundleStartMajId_i[26] bundleStartMajId_i[25]
+ bundleStartMajId_i[24] bundleStartMajId_i[23] bundleStartMajId_i[22] bundleStartMajId_i[21]
+ bundleStartMajId_i[20] bundleStartMajId_i[19] bundleStartMajId_i[18] bundleStartMajId_i[17]
+ bundleStartMajId_i[16] bundleStartMajId_i[15] bundleStartMajId_i[14] bundleStartMajId_i[13]
+ bundleStartMajId_i[12] bundleStartMajId_i[11] bundleStartMajId_i[10] bundleStartMajId_i[9]
+ bundleStartMajId_i[8] bundleStartMajId_i[7] bundleStartMajId_i[6] bundleStartMajId_i[5]
+ bundleStartMajId_i[4] bundleStartMajId_i[3] bundleStartMajId_i[2] bundleStartMajId_i[1]
+ bundleStartMajId_i[0] enable1_i enable2_i enable3_i enable4_i enable1_o enable2_o
+ enable3_o enable4_o instr1_o[31] instr1_o[30] instr1_o[29] instr1_o[28] instr1_o[27]
+ instr1_o[26] instr1_o[25] instr1_o[24] instr1_o[23] instr1_o[22] instr1_o[21] instr1_o[20]
+ instr1_o[19] instr1_o[18] instr1_o[17] instr1_o[16] instr1_o[15] instr1_o[14] instr1_o[13]
+ instr1_o[12] instr1_o[11] instr1_o[10] instr1_o[9] instr1_o[8] instr1_o[7] instr1_o[6]
+ instr1_o[5] instr1_o[4] instr1_o[3] instr1_o[2] instr1_o[1] instr1_o[0] instr2_o[31]
+ instr2_o[30] instr2_o[29] instr2_o[28] instr2_o[27] instr2_o[26] instr2_o[25] instr2_o[24]
+ instr2_o[23] instr2_o[22] instr2_o[21] instr2_o[20] instr2_o[19] instr2_o[18] instr2_o[17]
+ instr2_o[16] instr2_o[15] instr2_o[14] instr2_o[13] instr2_o[12] instr2_o[11] instr2_o[10]
+ instr2_o[9] instr2_o[8] instr2_o[7] instr2_o[6] instr2_o[5] instr2_o[4] instr2_o[3]
+ instr2_o[2] instr2_o[1] instr2_o[0] instr3_o[31] instr3_o[30] instr3_o[29] instr3_o[28]
+ instr3_o[27] instr3_o[26] instr3_o[25] instr3_o[24] instr3_o[23] instr3_o[22] instr3_o[21]
+ instr3_o[20] instr3_o[19] instr3_o[18] instr3_o[17] instr3_o[16] instr3_o[15] instr3_o[14]
+ instr3_o[13] instr3_o[12] instr3_o[11] instr3_o[10] instr3_o[9] instr3_o[8] instr3_o[7]
+ instr3_o[6] instr3_o[5] instr3_o[4] instr3_o[3] instr3_o[2] instr3_o[1] instr3_o[0]
+ instr4_o[31] instr4_o[30] instr4_o[29] instr4_o[28] instr4_o[27] instr4_o[26] instr4_o[25]
+ instr4_o[24] instr4_o[23] instr4_o[22] instr4_o[21] instr4_o[20] instr4_o[19] instr4_o[18]
+ instr4_o[17] instr4_o[16] instr4_o[15] instr4_o[14] instr4_o[13] instr4_o[12] instr4_o[11]
+ instr4_o[10] instr4_o[9] instr4_o[8] instr4_o[7] instr4_o[6] instr4_o[5] instr4_o[4]
+ instr4_o[3] instr4_o[2] instr4_o[1] instr4_o[0] addr1_o[63] addr1_o[62] addr1_o[61]
+ addr1_o[60] addr1_o[59] addr1_o[58] addr1_o[57] addr1_o[56] addr1_o[55] addr1_o[54]
+ addr1_o[53] addr1_o[52] addr1_o[51] addr1_o[50] addr1_o[49] addr1_o[48] addr1_o[47]
+ addr1_o[46] addr1_o[45] addr1_o[44] addr1_o[43] addr1_o[42] addr1_o[41] addr1_o[40]
+ addr1_o[39] addr1_o[38] addr1_o[37] addr1_o[36] addr1_o[35] addr1_o[34] addr1_o[33]
+ addr1_o[32] addr1_o[31] addr1_o[30] addr1_o[29] addr1_o[28] addr1_o[27] addr1_o[26]
+ addr1_o[25] addr1_o[24] addr1_o[23] addr1_o[22] addr1_o[21] addr1_o[20] addr1_o[19]
+ addr1_o[18] addr1_o[17] addr1_o[16] addr1_o[15] addr1_o[14] addr1_o[13] addr1_o[12]
+ addr1_o[11] addr1_o[10] addr1_o[9] addr1_o[8] addr1_o[7] addr1_o[6] addr1_o[5] addr1_o[4]
+ addr1_o[3] addr1_o[2] addr1_o[1] addr1_o[0] addr2_o[63] addr2_o[62] addr2_o[61]
+ addr2_o[60] addr2_o[59] addr2_o[58] addr2_o[57] addr2_o[56] addr2_o[55] addr2_o[54]
+ addr2_o[53] addr2_o[52] addr2_o[51] addr2_o[50] addr2_o[49] addr2_o[48] addr2_o[47]
+ addr2_o[46] addr2_o[45] addr2_o[44] addr2_o[43] addr2_o[42] addr2_o[41] addr2_o[40]
+ addr2_o[39] addr2_o[38] addr2_o[37] addr2_o[36] addr2_o[35] addr2_o[34] addr2_o[33]
+ addr2_o[32] addr2_o[31] addr2_o[30] addr2_o[29] addr2_o[28] addr2_o[27] addr2_o[26]
+ addr2_o[25] addr2_o[24] addr2_o[23] addr2_o[22] addr2_o[21] addr2_o[20] addr2_o[19]
+ addr2_o[18] addr2_o[17] addr2_o[16] addr2_o[15] addr2_o[14] addr2_o[13] addr2_o[12]
+ addr2_o[11] addr2_o[10] addr2_o[9] addr2_o[8] addr2_o[7] addr2_o[6] addr2_o[5] addr2_o[4]
+ addr2_o[3] addr2_o[2] addr2_o[1] addr2_o[0] addr3_o[63] addr3_o[62] addr3_o[61]
+ addr3_o[60] addr3_o[59] addr3_o[58] addr3_o[57] addr3_o[56] addr3_o[55] addr3_o[54]
+ addr3_o[53] addr3_o[52] addr3_o[51] addr3_o[50] addr3_o[49] addr3_o[48] addr3_o[47]
+ addr3_o[46] addr3_o[45] addr3_o[44] addr3_o[43] addr3_o[42] addr3_o[41] addr3_o[40]
+ addr3_o[39] addr3_o[38] addr3_o[37] addr3_o[36] addr3_o[35] addr3_o[34] addr3_o[33]
+ addr3_o[32] addr3_o[31] addr3_o[30] addr3_o[29] addr3_o[28] addr3_o[27] addr3_o[26]
+ addr3_o[25] addr3_o[24] addr3_o[23] addr3_o[22] addr3_o[21] addr3_o[20] addr3_o[19]
+ addr3_o[18] addr3_o[17] addr3_o[16] addr3_o[15] addr3_o[14] addr3_o[13] addr3_o[12]
+ addr3_o[11] addr3_o[10] addr3_o[9] addr3_o[8] addr3_o[7] addr3_o[6] addr3_o[5] addr3_o[4]
+ addr3_o[3] addr3_o[2] addr3_o[1] addr3_o[0] addr4_o[63] addr4_o[62] addr4_o[61]
+ addr4_o[60] addr4_o[59] addr4_o[58] addr4_o[57] addr4_o[56] addr4_o[55] addr4_o[54]
+ addr4_o[53] addr4_o[52] addr4_o[51] addr4_o[50] addr4_o[49] addr4_o[48] addr4_o[47]
+ addr4_o[46] addr4_o[45] addr4_o[44] addr4_o[43] addr4_o[42] addr4_o[41] addr4_o[40]
+ addr4_o[39] addr4_o[38] addr4_o[37] addr4_o[36] addr4_o[35] addr4_o[34] addr4_o[33]
+ addr4_o[32] addr4_o[31] addr4_o[30] addr4_o[29] addr4_o[28] addr4_o[27] addr4_o[26]
+ addr4_o[25] addr4_o[24] addr4_o[23] addr4_o[22] addr4_o[21] addr4_o[20] addr4_o[19]
+ addr4_o[18] addr4_o[17] addr4_o[16] addr4_o[15] addr4_o[14] addr4_o[13] addr4_o[12]
+ addr4_o[11] addr4_o[10] addr4_o[9] addr4_o[8] addr4_o[7] addr4_o[6] addr4_o[5] addr4_o[4]
+ addr4_o[3] addr4_o[2] addr4_o[1] addr4_o[0] is64b1_o is64b2_o is64b3_o is64b4_o
+ pid1_o[31] pid1_o[30] pid1_o[29] pid1_o[28] pid1_o[27] pid1_o[26] pid1_o[25] pid1_o[24]
+ pid1_o[23] pid1_o[22] pid1_o[21] pid1_o[20] pid1_o[19] pid1_o[18] pid1_o[17] pid1_o[16]
+ pid1_o[15] pid1_o[14] pid1_o[13] pid1_o[12] pid1_o[11] pid1_o[10] pid1_o[9] pid1_o[8]
+ pid1_o[7] pid1_o[6] pid1_o[5] pid1_o[4] pid1_o[3] pid1_o[2] pid1_o[1] pid1_o[0]
+ pid2_o[31] pid2_o[30] pid2_o[29] pid2_o[28] pid2_o[27] pid2_o[26] pid2_o[25] pid2_o[24]
+ pid2_o[23] pid2_o[22] pid2_o[21] pid2_o[20] pid2_o[19] pid2_o[18] pid2_o[17] pid2_o[16]
+ pid2_o[15] pid2_o[14] pid2_o[13] pid2_o[12] pid2_o[11] pid2_o[10] pid2_o[9] pid2_o[8]
+ pid2_o[7] pid2_o[6] pid2_o[5] pid2_o[4] pid2_o[3] pid2_o[2] pid2_o[1] pid2_o[0]
+ pid3_o[31] pid3_o[30] pid3_o[29] pid3_o[28] pid3_o[27] pid3_o[26] pid3_o[25] pid3_o[24]
+ pid3_o[23] pid3_o[22] pid3_o[21] pid3_o[20] pid3_o[19] pid3_o[18] pid3_o[17] pid3_o[16]
+ pid3_o[15] pid3_o[14] pid3_o[13] pid3_o[12] pid3_o[11] pid3_o[10] pid3_o[9] pid3_o[8]
+ pid3_o[7] pid3_o[6] pid3_o[5] pid3_o[4] pid3_o[3] pid3_o[2] pid3_o[1] pid3_o[0]
+ pid4_o[31] pid4_o[30] pid4_o[29] pid4_o[28] pid4_o[27] pid4_o[26] pid4_o[25] pid4_o[24]
+ pid4_o[23] pid4_o[22] pid4_o[21] pid4_o[20] pid4_o[19] pid4_o[18] pid4_o[17] pid4_o[16]
+ pid4_o[15] pid4_o[14] pid4_o[13] pid4_o[12] pid4_o[11] pid4_o[10] pid4_o[9] pid4_o[8]
+ pid4_o[7] pid4_o[6] pid4_o[5] pid4_o[4] pid4_o[3] pid4_o[2] pid4_o[1] pid4_o[0]
+ tid1_o[63] tid1_o[62] tid1_o[61] tid1_o[60] tid1_o[59] tid1_o[58] tid1_o[57] tid1_o[56]
+ tid1_o[55] tid1_o[54] tid1_o[53] tid1_o[52] tid1_o[51] tid1_o[50] tid1_o[49] tid1_o[48]
+ tid1_o[47] tid1_o[46] tid1_o[45] tid1_o[44] tid1_o[43] tid1_o[42] tid1_o[41] tid1_o[40]
+ tid1_o[39] tid1_o[38] tid1_o[37] tid1_o[36] tid1_o[35] tid1_o[34] tid1_o[33] tid1_o[32]
+ tid1_o[31] tid1_o[30] tid1_o[29] tid1_o[28] tid1_o[27] tid1_o[26] tid1_o[25] tid1_o[24]
+ tid1_o[23] tid1_o[22] tid1_o[21] tid1_o[20] tid1_o[19] tid1_o[18] tid1_o[17] tid1_o[16]
+ tid1_o[15] tid1_o[14] tid1_o[13] tid1_o[12] tid1_o[11] tid1_o[10] tid1_o[9] tid1_o[8]
+ tid1_o[7] tid1_o[6] tid1_o[5] tid1_o[4] tid1_o[3] tid1_o[2] tid1_o[1] tid1_o[0]
+ tid2_o[63] tid2_o[62] tid2_o[61] tid2_o[60] tid2_o[59] tid2_o[58] tid2_o[57] tid2_o[56]
+ tid2_o[55] tid2_o[54] tid2_o[53] tid2_o[52] tid2_o[51] tid2_o[50] tid2_o[49] tid2_o[48]
+ tid2_o[47] tid2_o[46] tid2_o[45] tid2_o[44] tid2_o[43] tid2_o[42] tid2_o[41] tid2_o[40]
+ tid2_o[39] tid2_o[38] tid2_o[37] tid2_o[36] tid2_o[35] tid2_o[34] tid2_o[33] tid2_o[32]
+ tid2_o[31] tid2_o[30] tid2_o[29] tid2_o[28] tid2_o[27] tid2_o[26] tid2_o[25] tid2_o[24]
+ tid2_o[23] tid2_o[22] tid2_o[21] tid2_o[20] tid2_o[19] tid2_o[18] tid2_o[17] tid2_o[16]
+ tid2_o[15] tid2_o[14] tid2_o[13] tid2_o[12] tid2_o[11] tid2_o[10] tid2_o[9] tid2_o[8]
+ tid2_o[7] tid2_o[6] tid2_o[5] tid2_o[4] tid2_o[3] tid2_o[2] tid2_o[1] tid2_o[0]
+ tid3_o[63] tid3_o[62] tid3_o[61] tid3_o[60] tid3_o[59] tid3_o[58] tid3_o[57] tid3_o[56]
+ tid3_o[55] tid3_o[54] tid3_o[53] tid3_o[52] tid3_o[51] tid3_o[50] tid3_o[49] tid3_o[48]
+ tid3_o[47] tid3_o[46] tid3_o[45] tid3_o[44] tid3_o[43] tid3_o[42] tid3_o[41] tid3_o[40]
+ tid3_o[39] tid3_o[38] tid3_o[37] tid3_o[36] tid3_o[35] tid3_o[34] tid3_o[33] tid3_o[32]
+ tid3_o[31] tid3_o[30] tid3_o[29] tid3_o[28] tid3_o[27] tid3_o[26] tid3_o[25] tid3_o[24]
+ tid3_o[23] tid3_o[22] tid3_o[21] tid3_o[20] tid3_o[19] tid3_o[18] tid3_o[17] tid3_o[16]
+ tid3_o[15] tid3_o[14] tid3_o[13] tid3_o[12] tid3_o[11] tid3_o[10] tid3_o[9] tid3_o[8]
+ tid3_o[7] tid3_o[6] tid3_o[5] tid3_o[4] tid3_o[3] tid3_o[2] tid3_o[1] tid3_o[0]
+ tid4_o[63] tid4_o[62] tid4_o[61] tid4_o[60] tid4_o[59] tid4_o[58] tid4_o[57] tid4_o[56]
+ tid4_o[55] tid4_o[54] tid4_o[53] tid4_o[52] tid4_o[51] tid4_o[50] tid4_o[49] tid4_o[48]
+ tid4_o[47] tid4_o[46] tid4_o[45] tid4_o[44] tid4_o[43] tid4_o[42] tid4_o[41] tid4_o[40]
+ tid4_o[39] tid4_o[38] tid4_o[37] tid4_o[36] tid4_o[35] tid4_o[34] tid4_o[33] tid4_o[32]
+ tid4_o[31] tid4_o[30] tid4_o[29] tid4_o[28] tid4_o[27] tid4_o[26] tid4_o[25] tid4_o[24]
+ tid4_o[23] tid4_o[22] tid4_o[21] tid4_o[20] tid4_o[19] tid4_o[18] tid4_o[17] tid4_o[16]
+ tid4_o[15] tid4_o[14] tid4_o[13] tid4_o[12] tid4_o[11] tid4_o[10] tid4_o[9] tid4_o[8]
+ tid4_o[7] tid4_o[6] tid4_o[5] tid4_o[4] tid4_o[3] tid4_o[2] tid4_o[1] tid4_o[0]
+ majID1_o[63] majID1_o[62] majID1_o[61] majID1_o[60] majID1_o[59] majID1_o[58] majID1_o[57]
+ majID1_o[56] majID1_o[55] majID1_o[54] majID1_o[53] majID1_o[52] majID1_o[51] majID1_o[50]
+ majID1_o[49] majID1_o[48] majID1_o[47] majID1_o[46] majID1_o[45] majID1_o[44] majID1_o[43]
+ majID1_o[42] majID1_o[41] majID1_o[40] majID1_o[39] majID1_o[38] majID1_o[37] majID1_o[36]
+ majID1_o[35] majID1_o[34] majID1_o[33] majID1_o[32] majID1_o[31] majID1_o[30] majID1_o[29]
+ majID1_o[28] majID1_o[27] majID1_o[26] majID1_o[25] majID1_o[24] majID1_o[23] majID1_o[22]
+ majID1_o[21] majID1_o[20] majID1_o[19] majID1_o[18] majID1_o[17] majID1_o[16] majID1_o[15]
+ majID1_o[14] majID1_o[13] majID1_o[12] majID1_o[11] majID1_o[10] majID1_o[9] majID1_o[8]
+ majID1_o[7] majID1_o[6] majID1_o[5] majID1_o[4] majID1_o[3] majID1_o[2] majID1_o[1]
+ majID1_o[0] majID2_o[63] majID2_o[62] majID2_o[61] majID2_o[60] majID2_o[59] majID2_o[58]
+ majID2_o[57] majID2_o[56] majID2_o[55] majID2_o[54] majID2_o[53] majID2_o[52] majID2_o[51]
+ majID2_o[50] majID2_o[49] majID2_o[48] majID2_o[47] majID2_o[46] majID2_o[45] majID2_o[44]
+ majID2_o[43] majID2_o[42] majID2_o[41] majID2_o[40] majID2_o[39] majID2_o[38] majID2_o[37]
+ majID2_o[36] majID2_o[35] majID2_o[34] majID2_o[33] majID2_o[32] majID2_o[31] majID2_o[30]
+ majID2_o[29] majID2_o[28] majID2_o[27] majID2_o[26] majID2_o[25] majID2_o[24] majID2_o[23]
+ majID2_o[22] majID2_o[21] majID2_o[20] majID2_o[19] majID2_o[18] majID2_o[17] majID2_o[16]
+ majID2_o[15] majID2_o[14] majID2_o[13] majID2_o[12] majID2_o[11] majID2_o[10] majID2_o[9]
+ majID2_o[8] majID2_o[7] majID2_o[6] majID2_o[5] majID2_o[4] majID2_o[3] majID2_o[2]
+ majID2_o[1] majID2_o[0] majID3_o[63] majID3_o[62] majID3_o[61] majID3_o[60] majID3_o[59]
+ majID3_o[58] majID3_o[57] majID3_o[56] majID3_o[55] majID3_o[54] majID3_o[53] majID3_o[52]
+ majID3_o[51] majID3_o[50] majID3_o[49] majID3_o[48] majID3_o[47] majID3_o[46] majID3_o[45]
+ majID3_o[44] majID3_o[43] majID3_o[42] majID3_o[41] majID3_o[40] majID3_o[39] majID3_o[38]
+ majID3_o[37] majID3_o[36] majID3_o[35] majID3_o[34] majID3_o[33] majID3_o[32] majID3_o[31]
+ majID3_o[30] majID3_o[29] majID3_o[28] majID3_o[27] majID3_o[26] majID3_o[25] majID3_o[24]
+ majID3_o[23] majID3_o[22] majID3_o[21] majID3_o[20] majID3_o[19] majID3_o[18] majID3_o[17]
+ majID3_o[16] majID3_o[15] majID3_o[14] majID3_o[13] majID3_o[12] majID3_o[11] majID3_o[10]
+ majID3_o[9] majID3_o[8] majID3_o[7] majID3_o[6] majID3_o[5] majID3_o[4] majID3_o[3]
+ majID3_o[2] majID3_o[1] majID3_o[0] majID4_o[63] majID4_o[62] majID4_o[61] majID4_o[60]
+ majID4_o[59] majID4_o[58] majID4_o[57] majID4_o[56] majID4_o[55] majID4_o[54] majID4_o[53]
+ majID4_o[52] majID4_o[51] majID4_o[50] majID4_o[49] majID4_o[48] majID4_o[47] majID4_o[46]
+ majID4_o[45] majID4_o[44] majID4_o[43] majID4_o[42] majID4_o[41] majID4_o[40] majID4_o[39]
+ majID4_o[38] majID4_o[37] majID4_o[36] majID4_o[35] majID4_o[34] majID4_o[33] majID4_o[32]
+ majID4_o[31] majID4_o[30] majID4_o[29] majID4_o[28] majID4_o[27] majID4_o[26] majID4_o[25]
+ majID4_o[24] majID4_o[23] majID4_o[22] majID4_o[21] majID4_o[20] majID4_o[19] majID4_o[18]
+ majID4_o[17] majID4_o[16] majID4_o[15] majID4_o[14] majID4_o[13] majID4_o[12] majID4_o[11]
+ majID4_o[10] majID4_o[9] majID4_o[8] majID4_o[7] majID4_o[6] majID4_o[5] majID4_o[4]
+ majID4_o[3] majID4_o[2] majID4_o[1] majID4_o[0]
XFILL_6_DFFPOSX1_728 gnd vdd FILL
XFILL_6_DFFPOSX1_739 gnd vdd FILL
XFILL_9_6_0 gnd vdd FILL
XFILL_2_OAI21X1_240 gnd vdd FILL
XFILL_5_DFFPOSX1_9 gnd vdd FILL
XNAND2X1_580 bundleAddress_i[6] INVX2_104/A gnd INVX1_197/A vdd NAND2X1
XNAND2X1_591 INVX1_183/A NAND2X1_591/B gnd NAND2X1_591/Y vdd NAND2X1
XFILL_0_NAND2X1_309 gnd vdd FILL
XFILL_17_5_0 gnd vdd FILL
XFILL_1_DFFPOSX1_1004 gnd vdd FILL
XFILL_1_DFFPOSX1_1026 gnd vdd FILL
XFILL_5_DFFPOSX1_318 gnd vdd FILL
XFILL_5_DFFPOSX1_307 gnd vdd FILL
XFILL_1_DFFPOSX1_1015 gnd vdd FILL
XFILL_5_DFFPOSX1_329 gnd vdd FILL
XOAI21X1_1804 BUFX4_336/Y INVX2_176/Y NAND2X1_745/Y gnd OAI21X1_1804/Y vdd OAI21X1
XFILL_22_11_1 gnd vdd FILL
XOAI21X1_1815 BUFX4_364/Y INVX2_187/Y NAND2X1_756/Y gnd OAI21X1_1815/Y vdd OAI21X1
XOAI21X1_1826 OAI21X1_2/A INVX2_198/Y NAND2X1_767/Y gnd OAI21X1_1826/Y vdd OAI21X1
XFILL_3_DFFPOSX1_791 gnd vdd FILL
XFILL_0_OAI21X1_804 gnd vdd FILL
XFILL_3_DFFPOSX1_780 gnd vdd FILL
XFILL_0_OAI21X1_837 gnd vdd FILL
XFILL_0_OAI21X1_826 gnd vdd FILL
XFILL_3_CLKBUF1_90 gnd vdd FILL
XFILL_0_OAI21X1_815 gnd vdd FILL
XFILL_0_OAI21X1_848 gnd vdd FILL
XFILL_0_OAI21X1_859 gnd vdd FILL
XFILL_2_DFFPOSX1_18 gnd vdd FILL
XFILL_2_DFFPOSX1_29 gnd vdd FILL
XFILL_0_OAI21X1_1614 gnd vdd FILL
XFILL_0_OAI21X1_1603 gnd vdd FILL
XFILL_0_OAI21X1_1625 gnd vdd FILL
XBUFX2_490 BUFX2_490/A gnd majID2_o[24] vdd BUFX2
XFILL_0_OAI21X1_1647 gnd vdd FILL
XFILL_0_OAI21X1_1636 gnd vdd FILL
XFILL_2_DFFPOSX1_392 gnd vdd FILL
XFILL_2_DFFPOSX1_381 gnd vdd FILL
XFILL_2_DFFPOSX1_370 gnd vdd FILL
XFILL_0_OAI21X1_1658 gnd vdd FILL
XFILL_0_OAI21X1_1669 gnd vdd FILL
XFILL_27_10_1 gnd vdd FILL
XFILL_5_DFFPOSX1_830 gnd vdd FILL
XFILL_5_DFFPOSX1_841 gnd vdd FILL
XFILL_5_DFFPOSX1_852 gnd vdd FILL
XFILL_5_DFFPOSX1_863 gnd vdd FILL
XFILL_5_DFFPOSX1_874 gnd vdd FILL
XFILL_5_DFFPOSX1_885 gnd vdd FILL
XFILL_5_DFFPOSX1_896 gnd vdd FILL
XFILL_1_XNOR2X1_31 gnd vdd FILL
XFILL_1_XNOR2X1_20 gnd vdd FILL
XFILL_1_XNOR2X1_64 gnd vdd FILL
XFILL_1_XNOR2X1_53 gnd vdd FILL
XFILL_1_XNOR2X1_42 gnd vdd FILL
XFILL_4_DFFPOSX1_1019 gnd vdd FILL
XFILL_1_XNOR2X1_75 gnd vdd FILL
XFILL_1_XNOR2X1_97 gnd vdd FILL
XFILL_4_DFFPOSX1_1008 gnd vdd FILL
XFILL_1_XNOR2X1_86 gnd vdd FILL
XFILL_4_DFFPOSX1_420 gnd vdd FILL
XFILL_4_DFFPOSX1_431 gnd vdd FILL
XFILL_4_DFFPOSX1_442 gnd vdd FILL
XFILL_4_DFFPOSX1_453 gnd vdd FILL
XFILL_4_DFFPOSX1_464 gnd vdd FILL
XFILL_0_INVX2_109 gnd vdd FILL
XFILL_4_DFFPOSX1_486 gnd vdd FILL
XFILL_4_DFFPOSX1_497 gnd vdd FILL
XFILL_4_DFFPOSX1_475 gnd vdd FILL
XFILL_2_11_1 gnd vdd FILL
XFILL_29_18_0 gnd vdd FILL
XFILL_1_BUFX2_310 gnd vdd FILL
XFILL_1_BUFX2_354 gnd vdd FILL
XFILL_1_BUFX2_343 gnd vdd FILL
XFILL_1_BUFX2_387 gnd vdd FILL
XOAI21X1_371 BUFX4_325/Y INVX4_21/Y OAI21X1_371/C gnd OAI21X1_371/Y vdd OAI21X1
XOAI21X1_360 BUFX4_346/Y OR2X2_15/B OAI21X1_360/C gnd OAI21X1_360/Y vdd OAI21X1
XOAI21X1_382 BUFX4_346/Y INVX1_3/Y OAI21X1_382/C gnd OAI21X1_382/Y vdd OAI21X1
XAND2X2_5 bundleStartMajId_i[42] bundleStartMajId_i[41] gnd AND2X2_5/Y vdd AND2X2
XFILL_1_BUFX2_398 gnd vdd FILL
XFILL_1_OAI21X1_1309 gnd vdd FILL
XOAI21X1_393 INVX1_6/Y BUFX4_244/Y OAI21X1_393/C gnd OAI21X1_393/Y vdd OAI21X1
XFILL_6_DFFPOSX1_525 gnd vdd FILL
XFILL_6_DFFPOSX1_536 gnd vdd FILL
XFILL_6_DFFPOSX1_503 gnd vdd FILL
XFILL_6_DFFPOSX1_514 gnd vdd FILL
XFILL_7_10_1 gnd vdd FILL
XFILL_0_NAND2X1_106 gnd vdd FILL
XFILL_0_INVX1_120 gnd vdd FILL
XFILL_0_INVX1_131 gnd vdd FILL
XFILL_0_NAND2X1_128 gnd vdd FILL
XFILL_0_NAND2X1_139 gnd vdd FILL
XFILL_0_NAND2X1_117 gnd vdd FILL
XFILL_0_INVX1_142 gnd vdd FILL
XFILL_0_INVX1_164 gnd vdd FILL
XFILL_1_AOI21X1_20 gnd vdd FILL
XFILL_1_AOI21X1_31 gnd vdd FILL
XFILL_0_INVX1_153 gnd vdd FILL
XFILL_1_AOI21X1_42 gnd vdd FILL
XFILL_33_8_1 gnd vdd FILL
XFILL_32_3_0 gnd vdd FILL
XFILL_0_INVX1_186 gnd vdd FILL
XFILL_1_AOI21X1_53 gnd vdd FILL
XFILL_0_INVX1_197 gnd vdd FILL
XFILL_0_INVX1_175 gnd vdd FILL
XFILL_1_AOI21X1_64 gnd vdd FILL
XFILL_5_DFFPOSX1_104 gnd vdd FILL
XFILL_5_DFFPOSX1_126 gnd vdd FILL
XFILL_5_DFFPOSX1_115 gnd vdd FILL
XFILL_5_DFFPOSX1_137 gnd vdd FILL
XFILL_5_DFFPOSX1_148 gnd vdd FILL
XFILL_5_DFFPOSX1_159 gnd vdd FILL
XOAI21X1_1623 INVX2_126/Y BUFX4_218/Y NAND2X1_691/Y gnd DFFPOSX1_13/D vdd OAI21X1
XOAI21X1_1601 BUFX4_339/Y INVX2_137/Y NAND2X1_670/Y gnd OAI21X1_1601/Y vdd OAI21X1
XOAI21X1_1612 BUFX4_320/Y INVX2_116/Y NAND2X1_681/Y gnd DFFPOSX1_3/D vdd OAI21X1
XFILL_1_OAI21X1_1821 gnd vdd FILL
XFILL_1_OAI21X1_1810 gnd vdd FILL
XOAI21X1_1634 INVX2_137/Y BUFX4_219/Y NAND2X1_702/Y gnd DFFPOSX1_24/D vdd OAI21X1
XOAI21X1_1656 BUFX4_1/A OAI21X1_7/A BUFX2_740/A gnd OAI21X1_1657/C vdd OAI21X1
XOAI21X1_1645 INVX2_116/Y BUFX4_217/Y NAND2X1_713/Y gnd DFFPOSX1_35/D vdd OAI21X1
XOAI21X1_1678 BUFX4_2/Y BUFX4_368/Y BUFX2_721/A gnd OAI21X1_1679/C vdd OAI21X1
XOAI21X1_1689 BUFX4_136/Y INVX2_138/Y OAI21X1_1689/C gnd DFFPOSX1_57/D vdd OAI21X1
XOAI21X1_1667 BUFX4_140/Y INVX2_127/Y OAI21X1_1667/C gnd DFFPOSX1_46/D vdd OAI21X1
XFILL_0_OAI21X1_612 gnd vdd FILL
XFILL_0_OAI21X1_623 gnd vdd FILL
XFILL_0_OAI21X1_601 gnd vdd FILL
XFILL_0_OAI21X1_656 gnd vdd FILL
XFILL_0_OAI21X1_645 gnd vdd FILL
XFILL_0_OAI21X1_634 gnd vdd FILL
XFILL_1_OAI21X1_827 gnd vdd FILL
XFILL_1_OAI21X1_805 gnd vdd FILL
XFILL_1_OAI21X1_816 gnd vdd FILL
XFILL_1_OAI21X1_838 gnd vdd FILL
XFILL_1_OAI21X1_849 gnd vdd FILL
XFILL_0_OAI21X1_667 gnd vdd FILL
XFILL_9_18_0 gnd vdd FILL
XFILL_0_OAI21X1_689 gnd vdd FILL
XFILL_0_OAI21X1_678 gnd vdd FILL
XFILL_1_AND2X2_13 gnd vdd FILL
XFILL_1_AND2X2_24 gnd vdd FILL
XFILL_3_DFFPOSX1_19 gnd vdd FILL
XFILL_13_16_1 gnd vdd FILL
XFILL_0_OAI21X1_1400 gnd vdd FILL
XFILL_0_NAND2X1_651 gnd vdd FILL
XFILL_0_OAI21X1_1433 gnd vdd FILL
XFILL_0_OAI21X1_1422 gnd vdd FILL
XFILL_0_OAI21X1_1411 gnd vdd FILL
XFILL_0_NAND2X1_640 gnd vdd FILL
XFILL_0_NAND2X1_662 gnd vdd FILL
XFILL_0_NAND2X1_673 gnd vdd FILL
XFILL_0_NAND2X1_684 gnd vdd FILL
XFILL_0_OAI21X1_1466 gnd vdd FILL
XFILL_24_8_1 gnd vdd FILL
XFILL_23_3_0 gnd vdd FILL
XFILL_0_OAI21X1_1455 gnd vdd FILL
XFILL_0_NAND2X1_695 gnd vdd FILL
XFILL_0_OAI21X1_1444 gnd vdd FILL
XFILL_0_OAI21X1_1477 gnd vdd FILL
XFILL_0_OAI21X1_1488 gnd vdd FILL
XFILL_0_OAI21X1_1499 gnd vdd FILL
XFILL_4_DFFPOSX1_6 gnd vdd FILL
XFILL_0_BUFX2_8 gnd vdd FILL
XFILL_5_DFFPOSX1_660 gnd vdd FILL
XFILL_5_DFFPOSX1_671 gnd vdd FILL
XFILL_5_DFFPOSX1_682 gnd vdd FILL
XFILL_5_DFFPOSX1_693 gnd vdd FILL
XFILL_18_15_1 gnd vdd FILL
XFILL_7_9_1 gnd vdd FILL
XFILL_6_4_0 gnd vdd FILL
XFILL_4_DFFPOSX1_261 gnd vdd FILL
XFILL_0_NAND2X1_19 gnd vdd FILL
XFILL_4_DFFPOSX1_272 gnd vdd FILL
XFILL_31_17_1 gnd vdd FILL
XFILL_4_DFFPOSX1_250 gnd vdd FILL
XFILL_4_DFFPOSX1_283 gnd vdd FILL
XFILL_12_11_0 gnd vdd FILL
XFILL_4_DFFPOSX1_294 gnd vdd FILL
XFILL_2_BUFX4_382 gnd vdd FILL
XFILL_15_8_1 gnd vdd FILL
XFILL_0_INVX2_8 gnd vdd FILL
XFILL_14_3_0 gnd vdd FILL
XFILL_1_BUFX2_151 gnd vdd FILL
XFILL_1_BUFX2_162 gnd vdd FILL
XFILL_1_BUFX2_140 gnd vdd FILL
XFILL_1_BUFX2_195 gnd vdd FILL
XFILL_1_BUFX2_184 gnd vdd FILL
XFILL_0_BUFX2_900 gnd vdd FILL
XFILL_0_BUFX2_911 gnd vdd FILL
XFILL_0_BUFX2_933 gnd vdd FILL
XFILL_0_BUFX2_922 gnd vdd FILL
XFILL_1_OAI21X1_1106 gnd vdd FILL
XFILL_1_OAI21X1_1128 gnd vdd FILL
XFILL_1_OAI21X1_1117 gnd vdd FILL
XINVX1_210 NOR3X1_18/A gnd INVX1_210/Y vdd INVX1
XDFFPOSX1_509 BUFX2_539/A CLKBUF1_60/Y OAI21X1_567/Y gnd vdd DFFPOSX1
XOAI21X1_190 BUFX4_6/A BUFX4_370/Y BUFX2_960/A gnd OAI21X1_191/C vdd OAI21X1
XFILL_0_BUFX2_944 gnd vdd FILL
XFILL_1_DFFPOSX1_718 gnd vdd FILL
XFILL_0_BUFX2_955 gnd vdd FILL
XINVX1_221 INVX1_221/A gnd INVX1_221/Y vdd INVX1
XFILL_1_DFFPOSX1_729 gnd vdd FILL
XFILL_0_BUFX2_966 gnd vdd FILL
XFILL_1_DFFPOSX1_707 gnd vdd FILL
XFILL_1_OAI21X1_1139 gnd vdd FILL
XFILL_0_BUFX2_999 gnd vdd FILL
XFILL_0_BUFX2_988 gnd vdd FILL
XFILL_0_BUFX2_977 gnd vdd FILL
XFILL_36_16_1 gnd vdd FILL
XFILL_17_10_0 gnd vdd FILL
XFILL_6_DFFPOSX1_377 gnd vdd FILL
XNAND2X1_32 BUFX2_858/A BUFX4_207/Y gnd OAI21X1_32/C vdd NAND2X1
XFILL_6_DFFPOSX1_399 gnd vdd FILL
XNAND2X1_43 BUFX2_870/A BUFX4_183/Y gnd OAI21X1_43/C vdd NAND2X1
XFILL_6_DFFPOSX1_388 gnd vdd FILL
XNAND2X1_10 BUFX2_853/A BUFX4_233/Y gnd OAI21X1_10/C vdd NAND2X1
XNAND2X1_21 BUFX2_846/A BUFX4_237/Y gnd OAI21X1_21/C vdd NAND2X1
XNAND2X1_65 BUFX2_894/A BUFX4_223/Y gnd OAI21X1_65/C vdd NAND2X1
XNAND2X1_54 BUFX2_882/A BUFX4_222/Y gnd OAI21X1_54/C vdd NAND2X1
XNAND2X1_76 BUFX2_427/A OAI21X1_6/A gnd NAND2X1_76/Y vdd NAND2X1
XFILL_30_12_0 gnd vdd FILL
XFILL_0_XNOR2X1_72 gnd vdd FILL
XNAND2X1_98 BUFX2_412/A BUFX4_378/Y gnd NAND2X1_98/Y vdd NAND2X1
XFILL_0_XNOR2X1_50 gnd vdd FILL
XNAND2X1_87 BUFX2_400/A BUFX4_388/Y gnd NAND2X1_87/Y vdd NAND2X1
XFILL_0_XNOR2X1_61 gnd vdd FILL
XFILL_0_XNOR2X1_83 gnd vdd FILL
XFILL_1_NAND2X1_118 gnd vdd FILL
XFILL_0_XNOR2X1_94 gnd vdd FILL
XFILL_1_NAND2X1_107 gnd vdd FILL
XFILL_0_DFFPOSX1_319 gnd vdd FILL
XFILL_35_1 gnd vdd FILL
XFILL_0_DFFPOSX1_308 gnd vdd FILL
XFILL_0_NOR3X1_15 gnd vdd FILL
XOAI21X1_1431 INVX2_105/Y INVX1_221/Y OAI21X1_1431/C gnd OAI21X1_1433/A vdd OAI21X1
XOAI21X1_1420 OAI21X1_1420/A AOI21X1_60/Y OAI21X1_1420/C gnd OAI21X1_1420/Y vdd OAI21X1
XFILL_1_OAI21X1_1651 gnd vdd FILL
XFILL_1_OAI21X1_1640 gnd vdd FILL
XOAI21X1_1475 XNOR2X1_99/Y BUFX4_301/Y OAI21X1_1475/C gnd OAI21X1_1475/Y vdd OAI21X1
XFILL_0_BUFX4_292 gnd vdd FILL
XOAI21X1_1464 INVX2_98/A INVX2_109/Y OAI21X1_1464/C gnd OAI21X1_1466/A vdd OAI21X1
XFILL_0_BUFX4_281 gnd vdd FILL
XFILL_0_BUFX4_270 gnd vdd FILL
XOAI21X1_1442 OAI21X1_1442/A INVX8_2/A OAI21X1_1442/C gnd OAI21X1_1442/Y vdd OAI21X1
XOAI21X1_1453 XNOR2X1_95/Y INVX8_2/A OAI21X1_1453/C gnd OAI21X1_1453/Y vdd OAI21X1
XFILL_4_NOR3X1_14 gnd vdd FILL
XFILL_1_OAI21X1_1662 gnd vdd FILL
XFILL_1_OAI21X1_1684 gnd vdd FILL
XFILL_1_OAI21X1_1673 gnd vdd FILL
XOAI21X1_1486 NOR2X1_154/A INVX1_223/A OAI21X1_1486/C gnd OAI21X1_1488/A vdd OAI21X1
XOAI21X1_1497 INVX1_223/A INVX2_100/Y INVX2_78/Y gnd NAND2X1_638/A vdd OAI21X1
XFILL_0_OAI21X1_420 gnd vdd FILL
XFILL_0_OAI21X1_431 gnd vdd FILL
XFILL_1_OAI21X1_602 gnd vdd FILL
XFILL_1_OAI21X1_1695 gnd vdd FILL
XFILL_1_OAI21X1_635 gnd vdd FILL
XFILL_0_OAI21X1_464 gnd vdd FILL
XFILL_1_NOR2X1_207 gnd vdd FILL
XFILL_1_OAI21X1_613 gnd vdd FILL
XFILL_1_OAI21X1_624 gnd vdd FILL
XFILL_0_OAI21X1_453 gnd vdd FILL
XFILL_0_OAI21X1_442 gnd vdd FILL
XFILL_1_OAI21X1_657 gnd vdd FILL
XFILL_1_OAI21X1_646 gnd vdd FILL
XFILL_0_OAI21X1_497 gnd vdd FILL
XFILL_0_OAI21X1_486 gnd vdd FILL
XFILL_0_OAI21X1_475 gnd vdd FILL
XFILL_1_OAI21X1_668 gnd vdd FILL
XFILL_3_NOR3X1_8 gnd vdd FILL
XFILL_1_OAI21X1_679 gnd vdd FILL
XFILL_35_11_0 gnd vdd FILL
XFILL_0_OAI21X1_1230 gnd vdd FILL
XFILL_0_OAI21X1_1241 gnd vdd FILL
XFILL_0_NAND2X1_470 gnd vdd FILL
XFILL_1_NAND2X1_641 gnd vdd FILL
XFILL_1_NAND2X1_630 gnd vdd FILL
XFILL_0_DFFPOSX1_820 gnd vdd FILL
XFILL_1_NAND2X1_652 gnd vdd FILL
XFILL_0_OAI21X1_1252 gnd vdd FILL
XFILL_0_NAND2X1_492 gnd vdd FILL
XFILL_0_NAND2X1_481 gnd vdd FILL
XFILL_0_OAI21X1_1263 gnd vdd FILL
XFILL_0_OAI21X1_1274 gnd vdd FILL
XFILL_0_DFFPOSX1_842 gnd vdd FILL
XFILL_1_NAND2X1_674 gnd vdd FILL
XFILL_1_NAND2X1_685 gnd vdd FILL
XFILL_0_DFFPOSX1_831 gnd vdd FILL
XFILL_0_DFFPOSX1_875 gnd vdd FILL
XFILL_1_NAND2X1_696 gnd vdd FILL
XFILL_0_DFFPOSX1_886 gnd vdd FILL
XFILL_0_OAI21X1_1285 gnd vdd FILL
XFILL_0_DFFPOSX1_853 gnd vdd FILL
XFILL_0_OAI21X1_1296 gnd vdd FILL
XFILL_0_DFFPOSX1_864 gnd vdd FILL
XDFFPOSX1_1027 BUFX2_665/A CLKBUF1_32/Y OAI21X1_1604/Y gnd vdd DFFPOSX1
XDFFPOSX1_1005 BUFX2_650/A CLKBUF1_65/Y OAI21X1_1582/Y gnd vdd DFFPOSX1
XDFFPOSX1_1016 BUFX2_653/A CLKBUF1_73/Y OAI21X1_1593/Y gnd vdd DFFPOSX1
XFILL_0_DFFPOSX1_897 gnd vdd FILL
XFILL_5_DFFPOSX1_490 gnd vdd FILL
XFILL_0_BUFX2_218 gnd vdd FILL
XFILL_0_BUFX2_229 gnd vdd FILL
XFILL_0_BUFX2_207 gnd vdd FILL
XFILL_0_AOI21X1_50 gnd vdd FILL
XFILL_0_AOI21X1_61 gnd vdd FILL
XFILL_2_DFFPOSX1_903 gnd vdd FILL
XFILL_2_DFFPOSX1_914 gnd vdd FILL
XFILL_2_OAI21X1_1324 gnd vdd FILL
XFILL_2_DFFPOSX1_936 gnd vdd FILL
XFILL_2_DFFPOSX1_947 gnd vdd FILL
XFILL_2_DFFPOSX1_925 gnd vdd FILL
XFILL_2_DFFPOSX1_958 gnd vdd FILL
XFILL_2_DFFPOSX1_969 gnd vdd FILL
XFILL_6_DFFPOSX1_1010 gnd vdd FILL
XFILL_6_DFFPOSX1_1032 gnd vdd FILL
XFILL_6_DFFPOSX1_1021 gnd vdd FILL
XFILL_30_6_1 gnd vdd FILL
XFILL_3_XNOR2X1_38 gnd vdd FILL
XFILL_3_XNOR2X1_27 gnd vdd FILL
XDFFPOSX1_306 BUFX2_975/A CLKBUF1_25/Y OAI21X1_229/Y gnd vdd DFFPOSX1
XDFFPOSX1_328 BUFX2_999/A CLKBUF1_7/Y OAI21X1_273/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_730 gnd vdd FILL
XDFFPOSX1_317 BUFX2_987/A CLKBUF1_27/Y OAI21X1_251/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_504 gnd vdd FILL
XFILL_0_BUFX2_741 gnd vdd FILL
XFILL_0_BUFX2_774 gnd vdd FILL
XFILL_0_BUFX2_752 gnd vdd FILL
XFILL_0_BUFX2_763 gnd vdd FILL
XDFFPOSX1_339 BUFX2_1011/A CLKBUF1_7/Y OAI21X1_295/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_785 gnd vdd FILL
XFILL_1_DFFPOSX1_515 gnd vdd FILL
XFILL_1_DFFPOSX1_537 gnd vdd FILL
XFILL_0_NOR2X1_92 gnd vdd FILL
XFILL_1_DFFPOSX1_526 gnd vdd FILL
XFILL_1_DFFPOSX1_548 gnd vdd FILL
XFILL_0_NOR2X1_81 gnd vdd FILL
XFILL_0_NOR2X1_70 gnd vdd FILL
XFILL_0_BUFX2_796 gnd vdd FILL
XNAND2X1_409 BUFX2_62/A BUFX4_353/Y gnd NAND2X1_409/Y vdd NAND2X1
XFILL_1_DFFPOSX1_559 gnd vdd FILL
XFILL_6_DFFPOSX1_130 gnd vdd FILL
XFILL_6_DFFPOSX1_152 gnd vdd FILL
XFILL_3_DFFPOSX1_3 gnd vdd FILL
XFILL_6_DFFPOSX1_141 gnd vdd FILL
XFILL_6_DFFPOSX1_185 gnd vdd FILL
XFILL_6_DFFPOSX1_163 gnd vdd FILL
XFILL_6_DFFPOSX1_174 gnd vdd FILL
XFILL_38_7_1 gnd vdd FILL
XFILL_37_2_0 gnd vdd FILL
XBUFX4_382 BUFX4_386/A gnd BUFX4_382/Y vdd BUFX4
XBUFX4_360 BUFX4_381/A gnd BUFX4_360/Y vdd BUFX4
XBUFX4_371 BUFX4_378/A gnd OAI21X1_5/A vdd BUFX4
XFILL_0_DFFPOSX1_105 gnd vdd FILL
XFILL_0_DFFPOSX1_127 gnd vdd FILL
XFILL_0_DFFPOSX1_138 gnd vdd FILL
XFILL_0_DFFPOSX1_116 gnd vdd FILL
XFILL_0_DFFPOSX1_149 gnd vdd FILL
XOAI21X1_915 BUFX4_143/Y INVX1_112/Y OAI21X1_915/C gnd OAI21X1_915/Y vdd OAI21X1
XFILL_21_6_1 gnd vdd FILL
XFILL_20_1_0 gnd vdd FILL
XOAI21X1_904 INVX1_105/Y BUFX4_189/Y OAI21X1_904/C gnd OAI21X1_904/Y vdd OAI21X1
XFILL_0_NAND2X1_3 gnd vdd FILL
XOAI21X1_948 BUFX4_11/Y BUFX4_341/Y BUFX2_338/A gnd OAI21X1_949/C vdd OAI21X1
XOAI21X1_937 BUFX4_143/Y INVX1_123/Y OAI21X1_937/C gnd OAI21X1_937/Y vdd OAI21X1
XFILL_3_DFFPOSX1_609 gnd vdd FILL
XOAI21X1_926 BUFX4_4/A OAI21X1_4/A BUFX2_356/A gnd OAI21X1_927/C vdd OAI21X1
XOAI21X1_959 BUFX4_154/Y INVX1_134/Y OAI21X1_959/C gnd OAI21X1_959/Y vdd OAI21X1
XFILL_21_17_0 gnd vdd FILL
XOAI21X1_1250 BUFX4_101/Y BUFX4_340/Y BUFX2_136/A gnd OAI21X1_1251/C vdd OAI21X1
XDFFPOSX1_840 BUFX2_91/A CLKBUF1_89/Y OAI21X1_1154/Y gnd vdd DFFPOSX1
XOAI21X1_1261 AOI21X1_46/Y OAI21X1_1261/B OAI21X1_1261/C gnd OAI21X1_1261/Y vdd OAI21X1
XDFFPOSX1_851 BUFX2_103/A CLKBUF1_89/Y OAI21X1_1170/Y gnd vdd DFFPOSX1
XOAI21X1_1283 BUFX4_6/A BUFX4_344/Y BUFX2_149/A gnd OAI21X1_1284/C vdd OAI21X1
XOAI21X1_1272 NOR3X1_18/C OR2X2_17/Y MUX2X1_2/S gnd NOR2X1_188/B vdd OAI21X1
XDFFPOSX1_884 BUFX2_133/A CLKBUF1_11/Y OAI21X1_1241/Y gnd vdd DFFPOSX1
XOAI21X1_1294 XNOR2X1_81/Y BUFX4_128/Y OAI21X1_1294/C gnd OAI21X1_1294/Y vdd OAI21X1
XFILL_1_OAI21X1_1481 gnd vdd FILL
XDFFPOSX1_873 BUFX2_130/A CLKBUF1_78/Y OAI21X1_1211/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1470 gnd vdd FILL
XFILL_1_OAI21X1_1492 gnd vdd FILL
XINVX2_12 bundleStartMajId_i[58] gnd INVX2_12/Y vdd INVX2
XDFFPOSX1_862 BUFX2_115/A CLKBUF1_20/Y OAI21X1_1189/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_410 gnd vdd FILL
XFILL_0_OAI21X1_261 gnd vdd FILL
XFILL_0_OAI21X1_272 gnd vdd FILL
XFILL_0_OAI21X1_250 gnd vdd FILL
XFILL_1_OAI21X1_454 gnd vdd FILL
XINVX2_34 bundleStartMajId_i[12] gnd INVX2_34/Y vdd INVX2
XINVX2_45 INVX2_45/A gnd INVX2_45/Y vdd INVX2
XFILL_2_OAI21X1_614 gnd vdd FILL
XINVX2_23 bundleStartMajId_i[33] gnd NOR3X1_7/A vdd INVX2
XDFFPOSX1_895 MUX2X1_2/B CLKBUF1_34/Y NOR2X1_189/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_421 gnd vdd FILL
XFILL_1_OAI21X1_432 gnd vdd FILL
XFILL_1_OAI21X1_443 gnd vdd FILL
XFILL_0_OAI21X1_294 gnd vdd FILL
XINVX2_67 bundleAddress_i[48] gnd INVX2_67/Y vdd INVX2
XINVX2_56 bundleAddress_i[60] gnd INVX2_56/Y vdd INVX2
XFILL_0_OAI21X1_283 gnd vdd FILL
XFILL_1_OAI21X1_476 gnd vdd FILL
XFILL_1_OAI21X1_487 gnd vdd FILL
XFILL_1_OAI21X1_465 gnd vdd FILL
XINVX2_78 bundleAddress_i[25] gnd INVX2_78/Y vdd INVX2
XFILL_1_OAI21X1_498 gnd vdd FILL
XFILL_2_OAI21X1_669 gnd vdd FILL
XINVX2_89 bundleAddress_i[5] gnd INVX2_89/Y vdd INVX2
XBUFX2_308 BUFX2_308/A gnd instr2_o[9] vdd BUFX2
XFILL_29_7_1 gnd vdd FILL
XFILL_28_2_0 gnd vdd FILL
XFILL_0_AOI21X1_8 gnd vdd FILL
XFILL_4_7_1 gnd vdd FILL
XFILL_3_2_0 gnd vdd FILL
XBUFX2_319 BUFX2_319/A gnd instr2_o[27] vdd BUFX2
XFILL_1_INVX4_23 gnd vdd FILL
XFILL_1_INVX4_45 gnd vdd FILL
XFILL_1_BUFX4_202 gnd vdd FILL
XFILL_1_BUFX4_213 gnd vdd FILL
XFILL_1_NAND2X1_460 gnd vdd FILL
XFILL_1_NAND2X1_471 gnd vdd FILL
XOAI21X1_19 INVX2_157/Y BUFX4_191/Y OAI21X1_19/C gnd OAI21X1_19/Y vdd OAI21X1
XFILL_1_BUFX4_235 gnd vdd FILL
XFILL_1_NAND2X1_493 gnd vdd FILL
XFILL_1_BUFX4_246 gnd vdd FILL
XFILL_1_NAND2X1_482 gnd vdd FILL
XFILL_0_DFFPOSX1_650 gnd vdd FILL
XFILL_0_OAI21X1_1082 gnd vdd FILL
XFILL_1_BUFX4_224 gnd vdd FILL
XFILL_0_DFFPOSX1_661 gnd vdd FILL
XFILL_0_OAI21X1_1071 gnd vdd FILL
XFILL_0_OAI21X1_1093 gnd vdd FILL
XFILL_0_OAI21X1_1060 gnd vdd FILL
XFILL_0_DFFPOSX1_672 gnd vdd FILL
XFILL_0_DFFPOSX1_683 gnd vdd FILL
XFILL_0_DFFPOSX1_694 gnd vdd FILL
XFILL_1_BUFX4_279 gnd vdd FILL
XFILL_1_BUFX4_257 gnd vdd FILL
XFILL_26_16_0 gnd vdd FILL
XFILL_12_6_1 gnd vdd FILL
XFILL_11_1_0 gnd vdd FILL
XFILL_1_BUFX4_268 gnd vdd FILL
XFILL_0_DFFPOSX1_17 gnd vdd FILL
XFILL_0_DFFPOSX1_39 gnd vdd FILL
XFILL_2_BUFX4_40 gnd vdd FILL
XFILL_0_DFFPOSX1_28 gnd vdd FILL
XFILL_2_XNOR2X1_6 gnd vdd FILL
XFILL_19_2_0 gnd vdd FILL
XFILL_2_DFFPOSX1_700 gnd vdd FILL
XBUFX2_820 BUFX2_820/A gnd tid1_o[15] vdd BUFX2
XFILL_2_DFFPOSX1_711 gnd vdd FILL
XFILL_2_DFFPOSX1_722 gnd vdd FILL
XFILL_2_OAI21X1_1132 gnd vdd FILL
XBUFX2_831 NAND2X1_2/A gnd tid1_o[5] vdd BUFX2
XFILL_2_DFFPOSX1_755 gnd vdd FILL
XFILL_2_DFFPOSX1_744 gnd vdd FILL
XFILL_2_DFFPOSX1_733 gnd vdd FILL
XFILL_2_OAI21X1_1187 gnd vdd FILL
XFILL_1_17_0 gnd vdd FILL
XBUFX2_842 NAND2X1_9/A gnd tid2_o[62] vdd BUFX2
XBUFX2_853 BUFX2_853/A gnd tid2_o[61] vdd BUFX2
XFILL_2_DFFPOSX1_766 gnd vdd FILL
XBUFX2_864 BUFX2_864/A gnd tid2_o[60] vdd BUFX2
XBUFX2_875 BUFX2_875/A gnd tid2_o[59] vdd BUFX2
XFILL_2_DFFPOSX1_788 gnd vdd FILL
XBUFX2_897 BUFX2_897/A gnd tid2_o[57] vdd BUFX2
XFILL_2_DFFPOSX1_777 gnd vdd FILL
XFILL_0_NOR2X1_204 gnd vdd FILL
XFILL_2_DFFPOSX1_799 gnd vdd FILL
XBUFX2_886 BUFX2_886/A gnd tid2_o[58] vdd BUFX2
XFILL_0_NOR2X1_215 gnd vdd FILL
XFILL_0_NOR2X1_226 gnd vdd FILL
XFILL_12_3 gnd vdd FILL
XFILL_3_CLKBUF1_6 gnd vdd FILL
XDFFPOSX1_103 BUFX2_800/A CLKBUF1_94/Y OAI21X1_1777/Y gnd vdd DFFPOSX1
XDFFPOSX1_114 BUFX2_783/A CLKBUF1_25/Y OAI21X1_1788/Y gnd vdd DFFPOSX1
XDFFPOSX1_125 BUFX2_795/A CLKBUF1_3/Y OAI21X1_1799/Y gnd vdd DFFPOSX1
XDFFPOSX1_136 BUFX2_807/A CLKBUF1_16/Y OAI21X1_1810/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_323 gnd vdd FILL
XFILL_1_DFFPOSX1_301 gnd vdd FILL
XFILL_1_DFFPOSX1_312 gnd vdd FILL
XFILL_0_BUFX2_560 gnd vdd FILL
XFILL_1_DFFPOSX1_345 gnd vdd FILL
XDFFPOSX1_147 BUFX2_819/A CLKBUF1_16/Y OAI21X1_1821/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_356 gnd vdd FILL
XDFFPOSX1_158 NAND2X1_2/A CLKBUF1_33/Y OAI21X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_169 BUFX2_886/A CLKBUF1_37/Y OAI21X1_13/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_582 gnd vdd FILL
XFILL_0_BUFX2_593 gnd vdd FILL
XFILL_1_DFFPOSX1_334 gnd vdd FILL
XFILL_0_BUFX2_571 gnd vdd FILL
XNAND2X1_217 BUFX2_492/A BUFX4_204/Y gnd OAI21X1_459/C vdd NAND2X1
XFILL_1_DFFPOSX1_378 gnd vdd FILL
XFILL_1_DFFPOSX1_367 gnd vdd FILL
XFILL_1_DFFPOSX1_389 gnd vdd FILL
XNAND2X1_206 bundleStartMajId_i[30] bundleStartMajId_i[29] gnd OR2X2_8/A vdd NAND2X1
XNAND2X1_239 BUFX2_503/A BUFX4_204/Y gnd OAI21X1_477/C vdd NAND2X1
XNAND2X1_228 BUFX2_498/A BUFX4_215/Y gnd OAI21X1_469/C vdd NAND2X1
XFILL_4_DFFPOSX1_816 gnd vdd FILL
XFILL_4_DFFPOSX1_838 gnd vdd FILL
XFILL_4_DFFPOSX1_805 gnd vdd FILL
XFILL_6_16_0 gnd vdd FILL
XFILL_4_DFFPOSX1_827 gnd vdd FILL
XFILL_4_DFFPOSX1_849 gnd vdd FILL
XFILL_4_CLKBUF1_61 gnd vdd FILL
XFILL_4_CLKBUF1_50 gnd vdd FILL
XFILL_10_14_1 gnd vdd FILL
XBUFX4_190 BUFX4_22/Y gnd BUFX4_190/Y vdd BUFX4
XFILL_0_BUFX2_10 gnd vdd FILL
XFILL_0_INVX1_90 gnd vdd FILL
XFILL_0_BUFX2_21 gnd vdd FILL
XFILL_4_CLKBUF1_72 gnd vdd FILL
XFILL_4_CLKBUF1_83 gnd vdd FILL
XFILL_4_CLKBUF1_94 gnd vdd FILL
XFILL_0_BUFX2_43 gnd vdd FILL
XFILL_0_BUFX2_54 gnd vdd FILL
XFILL_0_BUFX2_32 gnd vdd FILL
XFILL_0_BUFX2_65 gnd vdd FILL
XFILL_1_BUFX2_728 gnd vdd FILL
XFILL_0_BUFX2_87 gnd vdd FILL
XFILL_1_NOR2X1_46 gnd vdd FILL
XFILL_1_BUFX2_717 gnd vdd FILL
XFILL_0_BUFX2_76 gnd vdd FILL
XFILL_1_NOR2X1_24 gnd vdd FILL
XFILL_1_NOR2X1_57 gnd vdd FILL
XOAI21X1_712 INVX1_36/A OR2X2_5/A OR2X2_5/B gnd OAI21X1_713/C vdd OAI21X1
XFILL_1_BUFX2_739 gnd vdd FILL
XOAI21X1_723 BUFX4_142/Y BUFX4_37/Y BUFX2_600/A gnd OAI21X1_724/C vdd OAI21X1
XFILL_1_NOR2X1_68 gnd vdd FILL
XOAI21X1_701 NOR2X1_11/B NOR2X1_105/A OAI21X1_701/C gnd OAI21X1_703/A vdd OAI21X1
XFILL_0_BUFX2_98 gnd vdd FILL
XFILL_3_DFFPOSX1_406 gnd vdd FILL
XOAI21X1_745 XNOR2X1_48/Y BUFX4_295/Y OAI21X1_745/C gnd OAI21X1_745/Y vdd OAI21X1
XOAI21X1_756 BUFX4_142/Y BUFX4_54/Y BUFX2_613/A gnd OAI21X1_757/C vdd OAI21X1
XOAI21X1_734 INVX1_38/Y OR2X2_4/A BUFX4_287/Y gnd OAI21X1_736/A vdd OAI21X1
XOAI21X1_767 INVX1_42/Y BUFX4_287/Y OAI21X1_767/C gnd OAI21X1_767/Y vdd OAI21X1
XFILL_3_DFFPOSX1_428 gnd vdd FILL
XFILL_3_DFFPOSX1_417 gnd vdd FILL
XFILL_3_DFFPOSX1_439 gnd vdd FILL
XOAI21X1_778 OAI21X1_778/A BUFX4_299/Y OAI21X1_778/C gnd OAI21X1_778/Y vdd OAI21X1
XOAI21X1_789 OAI21X1_789/A BUFX4_300/Y OAI21X1_789/C gnd OAI21X1_789/Y vdd OAI21X1
XOAI21X1_1080 BUFX4_381/Y INVX1_177/Y NAND2X1_446/Y gnd OAI21X1_1080/Y vdd OAI21X1
XOAI21X1_1091 BUFX4_357/Y INVX4_45/Y NAND2X1_457/Y gnd OAI21X1_1091/Y vdd OAI21X1
XDFFPOSX1_670 BUFX2_308/A CLKBUF1_95/Y OAI21X1_898/Y gnd vdd DFFPOSX1
XDFFPOSX1_692 BUFX2_329/A CLKBUF1_61/Y OAI21X1_933/Y gnd vdd DFFPOSX1
XDFFPOSX1_681 BUFX2_326/A CLKBUF1_42/Y OAI21X1_911/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_890 gnd vdd FILL
XFILL_1_OAI21X1_262 gnd vdd FILL
XFILL_1_OAI21X1_251 gnd vdd FILL
XFILL_1_OAI21X1_240 gnd vdd FILL
XFILL_0_NOR2X1_1 gnd vdd FILL
XNAND2X1_740 BUFX2_795/A BUFX4_363/Y gnd NAND2X1_740/Y vdd NAND2X1
XNAND2X1_762 BUFX2_819/A BUFX4_336/Y gnd NAND2X1_762/Y vdd NAND2X1
XFILL_1_OAI21X1_295 gnd vdd FILL
XFILL_1_OAI21X1_273 gnd vdd FILL
XNAND2X1_751 BUFX2_807/A BUFX4_311/Y gnd NAND2X1_751/Y vdd NAND2X1
XFILL_1_OAI21X1_284 gnd vdd FILL
XFILL_2_OAI21X1_488 gnd vdd FILL
XFILL_15_13_1 gnd vdd FILL
XFILL_2_XNOR2X1_13 gnd vdd FILL
XBUFX2_105 BUFX2_105/A gnd addr2_o[18] vdd BUFX2
XFILL_2_XNOR2X1_46 gnd vdd FILL
XFILL_2_XNOR2X1_35 gnd vdd FILL
XBUFX2_116 BUFX2_116/A gnd addr2_o[8] vdd BUFX2
XFILL_2_XNOR2X1_24 gnd vdd FILL
XBUFX2_138 BUFX2_138/A gnd addr3_o[46] vdd BUFX2
XBUFX2_127 BUFX2_127/A gnd addr2_o[55] vdd BUFX2
XFILL_2_XNOR2X1_57 gnd vdd FILL
XBUFX2_149 BUFX2_149/A gnd addr3_o[36] vdd BUFX2
XFILL_2_XNOR2X1_79 gnd vdd FILL
XFILL_2_XNOR2X1_68 gnd vdd FILL
XFILL_1_NAND2X1_290 gnd vdd FILL
XFILL_0_DFFPOSX1_480 gnd vdd FILL
XFILL_0_DFFPOSX1_491 gnd vdd FILL
XBUFX2_1008 BUFX2_1008/A gnd tid4_o[19] vdd BUFX2
XBUFX2_1019 BUFX2_1019/A gnd tid4_o[9] vdd BUFX2
XFILL_3_DFFPOSX1_940 gnd vdd FILL
XFILL_3_DFFPOSX1_962 gnd vdd FILL
XFILL_3_DFFPOSX1_951 gnd vdd FILL
XFILL_3_DFFPOSX1_984 gnd vdd FILL
XFILL_3_DFFPOSX1_973 gnd vdd FILL
XFILL_3_DFFPOSX1_995 gnd vdd FILL
XFILL_1_DFFPOSX1_18 gnd vdd FILL
XFILL_1_DFFPOSX1_29 gnd vdd FILL
XFILL_33_14_1 gnd vdd FILL
XBUFX4_52 BUFX4_72/A gnd BUFX4_52/Y vdd BUFX4
XBUFX4_41 BUFX4_71/A gnd BUFX4_41/Y vdd BUFX4
XBUFX4_30 BUFX4_82/A gnd BUFX4_30/Y vdd BUFX4
XBUFX4_63 BUFX4_82/A gnd BUFX4_63/Y vdd BUFX4
XBUFX4_85 clock_i gnd BUFX4_85/Y vdd BUFX4
XBUFX4_96 BUFX4_1/A gnd BUFX4_96/Y vdd BUFX4
XBUFX4_74 BUFX4_82/A gnd BUFX4_74/Y vdd BUFX4
XFILL_0_OAI21X1_1807 gnd vdd FILL
XFILL_2_DFFPOSX1_541 gnd vdd FILL
XFILL_2_DFFPOSX1_530 gnd vdd FILL
XBUFX2_650 BUFX2_650/A gnd pid1_o[30] vdd BUFX2
XFILL_35_5_1 gnd vdd FILL
XFILL_34_0_0 gnd vdd FILL
XBUFX2_661 BUFX2_661/A gnd pid1_o[29] vdd BUFX2
XFILL_0_OAI21X1_1818 gnd vdd FILL
XBUFX2_672 BUFX2_672/A gnd pid1_o[28] vdd BUFX2
XFILL_2_DFFPOSX1_563 gnd vdd FILL
XFILL_0_OAI21X1_1829 gnd vdd FILL
XFILL_2_DFFPOSX1_574 gnd vdd FILL
XFILL_2_DFFPOSX1_552 gnd vdd FILL
XFILL_2_DFFPOSX1_585 gnd vdd FILL
XBUFX2_694 BUFX2_694/A gnd pid2_o[11] vdd BUFX2
XFILL_2_DFFPOSX1_596 gnd vdd FILL
XBUFX2_683 BUFX2_683/A gnd pid2_o[21] vdd BUFX2
XOR2X2_11 OR2X2_11/A bundleStartMajId_i[15] gnd OR2X2_11/Y vdd OR2X2
XFILL_1_DFFPOSX1_131 gnd vdd FILL
XOR2X2_4 OR2X2_4/A OR2X2_4/B gnd OR2X2_4/Y vdd OR2X2
XFILL_1_DFFPOSX1_120 gnd vdd FILL
XINVX2_190 bundleTid_i[19] gnd INVX2_190/Y vdd INVX2
XFILL_1_DFFPOSX1_153 gnd vdd FILL
XFILL_1_DFFPOSX1_164 gnd vdd FILL
XFILL_0_BUFX2_390 gnd vdd FILL
XFILL_2_AOI21X1_35 gnd vdd FILL
XFILL_1_DFFPOSX1_142 gnd vdd FILL
XFILL_38_13_1 gnd vdd FILL
XFILL_1_DFFPOSX1_175 gnd vdd FILL
XFILL_1_DFFPOSX1_197 gnd vdd FILL
XFILL_1_DFFPOSX1_186 gnd vdd FILL
XXNOR2X1_6 INVX1_10/A INVX4_7/Y gnd XNOR2X1_6/Y vdd XNOR2X1
XFILL_4_DFFPOSX1_613 gnd vdd FILL
XFILL_4_DFFPOSX1_602 gnd vdd FILL
XFILL_4_DFFPOSX1_624 gnd vdd FILL
XFILL_4_DFFPOSX1_635 gnd vdd FILL
XFILL_4_DFFPOSX1_646 gnd vdd FILL
XFILL_4_DFFPOSX1_679 gnd vdd FILL
XFILL_4_DFFPOSX1_668 gnd vdd FILL
XFILL_4_DFFPOSX1_657 gnd vdd FILL
XFILL_26_5_1 gnd vdd FILL
XFILL_25_0_0 gnd vdd FILL
XFILL_1_5_1 gnd vdd FILL
XFILL_0_0_0 gnd vdd FILL
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XFILL_1_BUFX2_536 gnd vdd FILL
XFILL_1_BUFX2_525 gnd vdd FILL
XFILL_1_BUFX2_569 gnd vdd FILL
XFILL_3_DFFPOSX1_203 gnd vdd FILL
XOAI21X1_520 BUFX4_7/A BUFX4_358/Y BUFX2_582/A gnd OAI21X1_521/C vdd OAI21X1
XOAI21X1_531 INVX4_30/Y OR2X2_1/A INVX4_4/Y gnd OAI21X1_532/C vdd OAI21X1
XFILL_3_DFFPOSX1_214 gnd vdd FILL
XFILL_3_DFFPOSX1_225 gnd vdd FILL
XOAI21X1_553 OR2X2_10/B OR2X2_5/A OR2X2_5/B gnd OAI21X1_554/C vdd OAI21X1
XOAI21X1_575 NOR2X1_70/B OAI21X1_575/B INVX4_13/Y gnd NAND3X1_16/C vdd OAI21X1
XOAI21X1_542 BUFX4_93/Y BUFX4_372/Y BUFX2_528/A gnd OAI21X1_543/C vdd OAI21X1
XFILL_3_DFFPOSX1_236 gnd vdd FILL
XOAI21X1_564 BUFX4_10/A BUFX4_383/Y BUFX2_538/A gnd OAI21X1_565/C vdd OAI21X1
XFILL_3_DFFPOSX1_258 gnd vdd FILL
XFILL_3_DFFPOSX1_247 gnd vdd FILL
XOAI21X1_597 OR2X2_9/A INVX2_48/Y INVX2_26/Y gnd OAI21X1_598/C vdd OAI21X1
XFILL_3_DFFPOSX1_269 gnd vdd FILL
XOAI21X1_586 XNOR2X1_34/Y BUFX4_131/Y OAI21X1_586/C gnd OAI21X1_586/Y vdd OAI21X1
XFILL_6_DFFPOSX1_718 gnd vdd FILL
XFILL_6_DFFPOSX1_707 gnd vdd FILL
XFILL_9_6_1 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XNAND2X1_581 BUFX4_242/Y NAND2X1_581/B gnd NAND2X1_581/Y vdd NAND2X1
XNAND2X1_570 BUFX2_113/A BUFX4_201/Y gnd NAND2X1_570/Y vdd NAND2X1
XNAND2X1_592 bundleAddress_i[54] bundleAddress_i[53] gnd NOR2X1_180/B vdd NAND2X1
XFILL_2_OAI21X1_285 gnd vdd FILL
XFILL_17_5_1 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XFILL_1_DFFPOSX1_1027 gnd vdd FILL
XFILL_1_DFFPOSX1_1005 gnd vdd FILL
XFILL_5_DFFPOSX1_308 gnd vdd FILL
XFILL_1_DFFPOSX1_1016 gnd vdd FILL
XFILL_5_DFFPOSX1_319 gnd vdd FILL
XOAI21X1_1805 BUFX4_366/Y INVX2_177/Y NAND2X1_746/Y gnd OAI21X1_1805/Y vdd OAI21X1
XOAI21X1_1827 BUFX4_380/Y INVX2_199/Y NAND2X1_768/Y gnd OAI21X1_1827/Y vdd OAI21X1
XOAI21X1_1816 BUFX4_384/Y INVX2_188/Y NAND2X1_757/Y gnd OAI21X1_1816/Y vdd OAI21X1
XFILL_3_DFFPOSX1_792 gnd vdd FILL
XFILL_0_OAI21X1_805 gnd vdd FILL
XFILL_3_DFFPOSX1_770 gnd vdd FILL
XFILL_3_DFFPOSX1_781 gnd vdd FILL
XFILL_0_OAI21X1_838 gnd vdd FILL
XFILL_0_OAI21X1_827 gnd vdd FILL
XFILL_3_CLKBUF1_91 gnd vdd FILL
XFILL_3_CLKBUF1_80 gnd vdd FILL
XFILL_0_OAI21X1_816 gnd vdd FILL
XFILL_0_OAI21X1_849 gnd vdd FILL
XFILL_2_DFFPOSX1_19 gnd vdd FILL
XFILL_0_OAI21X1_1604 gnd vdd FILL
XFILL_0_OAI21X1_1615 gnd vdd FILL
XFILL_0_OAI21X1_1637 gnd vdd FILL
XFILL_0_OAI21X1_1648 gnd vdd FILL
XFILL_2_DFFPOSX1_382 gnd vdd FILL
XFILL_0_OAI21X1_1626 gnd vdd FILL
XBUFX2_480 BUFX2_480/A gnd majID2_o[60] vdd BUFX2
XFILL_2_DFFPOSX1_360 gnd vdd FILL
XFILL_2_DFFPOSX1_371 gnd vdd FILL
XFILL_0_OAI21X1_1659 gnd vdd FILL
XFILL_2_DFFPOSX1_393 gnd vdd FILL
XBUFX2_491 BUFX2_491/A gnd majID2_o[59] vdd BUFX2
XFILL_5_DFFPOSX1_820 gnd vdd FILL
XFILL_5_DFFPOSX1_831 gnd vdd FILL
XFILL_5_DFFPOSX1_853 gnd vdd FILL
XFILL_5_DFFPOSX1_842 gnd vdd FILL
XFILL_5_DFFPOSX1_864 gnd vdd FILL
XFILL_5_DFFPOSX1_875 gnd vdd FILL
XFILL_5_DFFPOSX1_886 gnd vdd FILL
XFILL_1_XNOR2X1_21 gnd vdd FILL
XFILL_5_DFFPOSX1_897 gnd vdd FILL
XFILL_1_XNOR2X1_10 gnd vdd FILL
XFILL_1_XNOR2X1_32 gnd vdd FILL
XFILL_1_XNOR2X1_43 gnd vdd FILL
XFILL_1_XNOR2X1_54 gnd vdd FILL
XFILL_1_XNOR2X1_76 gnd vdd FILL
XFILL_1_XNOR2X1_98 gnd vdd FILL
XFILL_1_XNOR2X1_65 gnd vdd FILL
XFILL_1_XNOR2X1_87 gnd vdd FILL
XFILL_4_DFFPOSX1_1009 gnd vdd FILL
XFILL_4_DFFPOSX1_421 gnd vdd FILL
XFILL_4_DFFPOSX1_410 gnd vdd FILL
XFILL_4_DFFPOSX1_443 gnd vdd FILL
XFILL_4_DFFPOSX1_432 gnd vdd FILL
XFILL_4_DFFPOSX1_454 gnd vdd FILL
XFILL_4_DFFPOSX1_476 gnd vdd FILL
XFILL_4_DFFPOSX1_487 gnd vdd FILL
XFILL_4_DFFPOSX1_465 gnd vdd FILL
XFILL_4_DFFPOSX1_498 gnd vdd FILL
XFILL_29_18_1 gnd vdd FILL
XFILL_1_BUFX2_322 gnd vdd FILL
XFILL_1_BUFX2_333 gnd vdd FILL
XFILL_1_BUFX2_344 gnd vdd FILL
XFILL_1_BUFX2_388 gnd vdd FILL
XFILL_1_BUFX2_366 gnd vdd FILL
XFILL_23_14_0 gnd vdd FILL
XFILL_1_BUFX2_377 gnd vdd FILL
XOAI21X1_350 BUFX4_337/Y INVX2_21/Y NAND2X1_94/Y gnd OAI21X1_350/Y vdd OAI21X1
XAND2X2_6 bundleStartMajId_i[34] bundleStartMajId_i[33] gnd AND2X2_6/Y vdd AND2X2
XOAI21X1_372 BUFX4_372/Y NOR3X1_2/A OAI21X1_372/C gnd OAI21X1_372/Y vdd OAI21X1
XOAI21X1_383 BUFX4_335/Y INVX2_36/Y OAI21X1_383/C gnd OAI21X1_383/Y vdd OAI21X1
XOAI21X1_361 BUFX4_373/Y INVX4_15/Y OAI21X1_361/C gnd OAI21X1_361/Y vdd OAI21X1
XOAI21X1_394 INVX4_1/Y INVX2_8/Y INVX2_9/Y gnd OAI21X1_395/C vdd OAI21X1
XFILL_6_DFFPOSX1_559 gnd vdd FILL
XFILL_0_NAND2X1_107 gnd vdd FILL
XFILL_0_INVX1_110 gnd vdd FILL
XFILL_0_INVX1_121 gnd vdd FILL
XFILL_0_NAND2X1_129 gnd vdd FILL
XFILL_0_NAND2X1_118 gnd vdd FILL
XFILL_0_INVX1_154 gnd vdd FILL
XFILL_0_INVX1_143 gnd vdd FILL
XFILL_1_AOI21X1_21 gnd vdd FILL
XFILL_1_AOI21X1_10 gnd vdd FILL
XFILL_1_AOI21X1_32 gnd vdd FILL
XFILL_0_INVX1_132 gnd vdd FILL
XFILL_0_INVX1_165 gnd vdd FILL
XFILL_0_INVX1_176 gnd vdd FILL
XFILL_1_AOI21X1_54 gnd vdd FILL
XFILL_1_AOI21X1_65 gnd vdd FILL
XFILL_0_INVX1_198 gnd vdd FILL
XFILL_1_AOI21X1_43 gnd vdd FILL
XFILL_0_INVX1_187 gnd vdd FILL
XFILL_32_3_1 gnd vdd FILL
XFILL_28_13_0 gnd vdd FILL
XFILL_5_DFFPOSX1_116 gnd vdd FILL
XFILL_5_DFFPOSX1_105 gnd vdd FILL
XFILL_5_DFFPOSX1_127 gnd vdd FILL
XFILL_5_DFFPOSX1_138 gnd vdd FILL
XFILL_5_DFFPOSX1_149 gnd vdd FILL
XFILL_1_OAI21X1_1800 gnd vdd FILL
XOAI21X1_1613 bundleLen_i[1] bundleLen_i[0] INVX8_4/A gnd BUFX4_26/A vdd OAI21X1
XOAI21X1_1602 BUFX4_352/Y INVX2_138/Y NAND2X1_671/Y gnd OAI21X1_1602/Y vdd OAI21X1
XOAI21X1_1624 INVX2_127/Y BUFX4_195/Y NAND2X1_692/Y gnd DFFPOSX1_14/D vdd OAI21X1
XFILL_1_OAI21X1_1811 gnd vdd FILL
XFILL_1_OAI21X1_1822 gnd vdd FILL
XOAI21X1_1646 BUFX4_5/Y BUFX4_341/Y BUFX2_713/A gnd OAI21X1_1647/C vdd OAI21X1
XOAI21X1_1635 INVX2_138/Y BUFX4_211/Y NAND2X1_703/Y gnd DFFPOSX1_25/D vdd OAI21X1
XOAI21X1_1657 BUFX4_154/Y INVX2_122/Y OAI21X1_1657/C gnd DFFPOSX1_41/D vdd OAI21X1
XOAI21X1_1679 BUFX4_126/Y INVX2_133/Y OAI21X1_1679/C gnd DFFPOSX1_52/D vdd OAI21X1
XOAI21X1_1668 BUFX4_101/Y BUFX4_347/Y BUFX2_716/A gnd OAI21X1_1669/C vdd OAI21X1
XFILL_0_OAI21X1_613 gnd vdd FILL
XFILL_0_OAI21X1_602 gnd vdd FILL
XFILL_0_OAI21X1_646 gnd vdd FILL
XFILL_0_OAI21X1_635 gnd vdd FILL
XFILL_1_OAI21X1_828 gnd vdd FILL
XFILL_1_OAI21X1_806 gnd vdd FILL
XFILL_0_OAI21X1_624 gnd vdd FILL
XFILL_1_OAI21X1_817 gnd vdd FILL
XFILL_0_OAI21X1_657 gnd vdd FILL
XFILL_1_OAI21X1_839 gnd vdd FILL
XFILL_0_OAI21X1_668 gnd vdd FILL
XFILL_9_18_1 gnd vdd FILL
XFILL_0_OAI21X1_679 gnd vdd FILL
XFILL_1_AND2X2_14 gnd vdd FILL
XFILL_1_AND2X2_25 gnd vdd FILL
XFILL_3_14_0 gnd vdd FILL
XFILL_0_NAND2X1_663 gnd vdd FILL
XFILL_0_NAND2X1_652 gnd vdd FILL
XFILL_0_OAI21X1_1401 gnd vdd FILL
XFILL_0_OAI21X1_1423 gnd vdd FILL
XFILL_0_OAI21X1_1412 gnd vdd FILL
XFILL_0_NAND2X1_641 gnd vdd FILL
XFILL_0_NAND2X1_630 gnd vdd FILL
XFILL_2_DFFPOSX1_190 gnd vdd FILL
XFILL_0_NAND2X1_696 gnd vdd FILL
XFILL_0_OAI21X1_1434 gnd vdd FILL
XFILL_0_OAI21X1_1456 gnd vdd FILL
XFILL_0_OAI21X1_1467 gnd vdd FILL
XFILL_0_OAI21X1_1445 gnd vdd FILL
XFILL_0_NAND2X1_674 gnd vdd FILL
XFILL_0_NAND2X1_685 gnd vdd FILL
XFILL_0_OAI21X1_1478 gnd vdd FILL
XFILL_23_3_1 gnd vdd FILL
XFILL_0_OAI21X1_1489 gnd vdd FILL
XFILL_4_DFFPOSX1_7 gnd vdd FILL
XFILL_5_DFFPOSX1_672 gnd vdd FILL
XFILL_0_BUFX2_9 gnd vdd FILL
XFILL_5_DFFPOSX1_650 gnd vdd FILL
XFILL_5_DFFPOSX1_661 gnd vdd FILL
XFILL_5_DFFPOSX1_683 gnd vdd FILL
XFILL_5_DFFPOSX1_694 gnd vdd FILL
XFILL_8_13_0 gnd vdd FILL
XFILL_6_4_1 gnd vdd FILL
XFILL_4_DFFPOSX1_262 gnd vdd FILL
XFILL_4_DFFPOSX1_240 gnd vdd FILL
XFILL_4_DFFPOSX1_251 gnd vdd FILL
XFILL_2_OAI21X1_1528 gnd vdd FILL
XFILL_4_DFFPOSX1_273 gnd vdd FILL
XFILL_4_DFFPOSX1_284 gnd vdd FILL
XFILL_4_DFFPOSX1_295 gnd vdd FILL
XFILL_12_11_1 gnd vdd FILL
XFILL_2_BUFX4_350 gnd vdd FILL
XFILL_0_INVX2_9 gnd vdd FILL
XFILL_14_3_1 gnd vdd FILL
XFILL_1_BUFX2_141 gnd vdd FILL
XFILL_1_BUFX2_130 gnd vdd FILL
XFILL_1_BUFX2_185 gnd vdd FILL
XFILL_1_BUFX2_174 gnd vdd FILL
XFILL_0_BUFX2_912 gnd vdd FILL
XOAI21X1_180 BUFX4_247/Y BUFX4_352/Y BUFX2_955/A gnd OAI21X1_181/C vdd OAI21X1
XINVX1_200 INVX1_200/A gnd INVX1_200/Y vdd INVX1
XFILL_1_OAI21X1_1107 gnd vdd FILL
XFILL_0_BUFX2_923 gnd vdd FILL
XFILL_1_OAI21X1_1118 gnd vdd FILL
XFILL_1_OAI21X1_1129 gnd vdd FILL
XFILL_0_BUFX2_934 gnd vdd FILL
XFILL_0_BUFX2_901 gnd vdd FILL
XOAI21X1_191 BUFX4_169/Y INVX2_3/Y OAI21X1_191/C gnd OAI21X1_191/Y vdd OAI21X1
XFILL_0_BUFX2_945 gnd vdd FILL
XINVX1_211 INVX1_211/A gnd INVX1_211/Y vdd INVX1
XFILL_0_BUFX2_956 gnd vdd FILL
XINVX1_222 INVX1_222/A gnd INVX1_222/Y vdd INVX1
XFILL_1_DFFPOSX1_719 gnd vdd FILL
XFILL_1_DFFPOSX1_708 gnd vdd FILL
XFILL_0_BUFX2_967 gnd vdd FILL
XFILL_0_BUFX2_989 gnd vdd FILL
XFILL_0_BUFX2_978 gnd vdd FILL
XFILL_6_DFFPOSX1_323 gnd vdd FILL
XFILL_6_DFFPOSX1_312 gnd vdd FILL
XFILL_6_DFFPOSX1_334 gnd vdd FILL
XFILL_6_DFFPOSX1_345 gnd vdd FILL
XFILL_6_DFFPOSX1_356 gnd vdd FILL
XFILL_6_DFFPOSX1_367 gnd vdd FILL
XNAND2X1_22 BUFX2_847/A BUFX4_218/Y gnd OAI21X1_22/C vdd NAND2X1
XNAND2X1_33 BUFX2_859/A BUFX4_191/Y gnd OAI21X1_33/C vdd NAND2X1
XFILL_17_10_1 gnd vdd FILL
XNAND2X1_11 BUFX2_864/A BUFX4_222/Y gnd OAI21X1_11/C vdd NAND2X1
XNAND2X1_55 BUFX2_883/A BUFX4_207/Y gnd OAI21X1_55/C vdd NAND2X1
XNAND2X1_44 BUFX2_871/A BUFX4_223/Y gnd OAI21X1_44/C vdd NAND2X1
XNAND2X1_66 BUFX2_895/A BUFX4_190/Y gnd OAI21X1_66/C vdd NAND2X1
XNAND2X1_77 BUFX2_438/A BUFX4_355/Y gnd NAND2X1_77/Y vdd NAND2X1
XFILL_30_12_1 gnd vdd FILL
XFILL_0_XNOR2X1_62 gnd vdd FILL
XFILL_0_XNOR2X1_51 gnd vdd FILL
XFILL_0_XNOR2X1_40 gnd vdd FILL
XNAND2X1_88 BUFX2_401/A BUFX4_355/Y gnd NAND2X1_88/Y vdd NAND2X1
XNAND2X1_99 BUFX2_413/A BUFX4_383/Y gnd NAND2X1_99/Y vdd NAND2X1
XFILL_0_XNOR2X1_73 gnd vdd FILL
XFILL_1_NAND2X1_119 gnd vdd FILL
XFILL_0_XNOR2X1_95 gnd vdd FILL
XFILL_0_XNOR2X1_84 gnd vdd FILL
XFILL_0_DFFPOSX1_309 gnd vdd FILL
XFILL_35_2 gnd vdd FILL
XFILL_28_1 gnd vdd FILL
XFILL_0_NOR3X1_16 gnd vdd FILL
XOAI21X1_1432 BUFX4_127/Y BUFX4_44/Y BUFX2_201/A gnd OAI21X1_1433/C vdd OAI21X1
XOAI21X1_1421 INVX2_108/Y INVX2_96/A INVX2_65/Y gnd OAI21X1_1422/C vdd OAI21X1
XOAI21X1_1410 INVX2_94/Y INVX4_50/Y OAI21X1_1410/C gnd OAI21X1_1412/A vdd OAI21X1
XFILL_0_BUFX4_260 gnd vdd FILL
XFILL_1_OAI21X1_1630 gnd vdd FILL
XFILL_0_BUFX4_293 gnd vdd FILL
XOAI21X1_1465 BUFX4_138/Y BUFX4_55/Y BUFX2_214/A gnd OAI21X1_1466/C vdd OAI21X1
XFILL_0_BUFX4_282 gnd vdd FILL
XOAI21X1_1454 BUFX4_174/Y BUFX4_71/Y BUFX2_210/A gnd OAI21X1_1455/C vdd OAI21X1
XFILL_0_BUFX4_271 gnd vdd FILL
XOAI21X1_1443 NOR2X1_221/Y bundleAddress_i[43] BUFX4_286/Y gnd OAI21X1_1445/B vdd
+ OAI21X1
XFILL_1_OAI21X1_1641 gnd vdd FILL
XFILL_1_OAI21X1_1674 gnd vdd FILL
XFILL_1_OAI21X1_1663 gnd vdd FILL
XFILL_1_OAI21X1_1652 gnd vdd FILL
XOAI21X1_1476 XNOR2X1_99/A INVX4_39/Y INVX2_74/Y gnd OAI21X1_1477/C vdd OAI21X1
XFILL_1_OAI21X1_1685 gnd vdd FILL
XFILL_1_OAI21X1_603 gnd vdd FILL
XFILL_0_OAI21X1_421 gnd vdd FILL
XOAI21X1_1487 BUFX4_152/Y BUFX4_28/Y BUFX2_222/A gnd OAI21X1_1488/C vdd OAI21X1
XFILL_0_OAI21X1_410 gnd vdd FILL
XOAI21X1_1498 BUFX4_152/Y BUFX4_78/Y BUFX2_225/A gnd OAI21X1_1499/C vdd OAI21X1
XFILL_1_OAI21X1_1696 gnd vdd FILL
XFILL_0_OAI21X1_454 gnd vdd FILL
XFILL_1_OAI21X1_614 gnd vdd FILL
XFILL_1_OAI21X1_636 gnd vdd FILL
XFILL_0_OAI21X1_465 gnd vdd FILL
XFILL_1_OAI21X1_625 gnd vdd FILL
XFILL_0_OAI21X1_432 gnd vdd FILL
XFILL_0_OAI21X1_443 gnd vdd FILL
XFILL_1_OAI21X1_647 gnd vdd FILL
XFILL_2_OAI21X1_829 gnd vdd FILL
XFILL_0_OAI21X1_498 gnd vdd FILL
XFILL_0_OAI21X1_476 gnd vdd FILL
XFILL_0_OAI21X1_487 gnd vdd FILL
XFILL_1_OAI21X1_658 gnd vdd FILL
XFILL_19_18_0 gnd vdd FILL
XFILL_1_OAI21X1_669 gnd vdd FILL
XFILL_3_NOR3X1_9 gnd vdd FILL
XFILL_35_11_1 gnd vdd FILL
XFILL_0_DFFPOSX1_810 gnd vdd FILL
XFILL_0_NAND2X1_471 gnd vdd FILL
XFILL_0_OAI21X1_1231 gnd vdd FILL
XFILL_0_OAI21X1_1242 gnd vdd FILL
XFILL_0_OAI21X1_1220 gnd vdd FILL
XFILL_1_NAND2X1_642 gnd vdd FILL
XFILL_1_NAND2X1_631 gnd vdd FILL
XFILL_0_NAND2X1_460 gnd vdd FILL
XFILL_1_NAND2X1_620 gnd vdd FILL
XFILL_0_DFFPOSX1_821 gnd vdd FILL
XFILL_0_DFFPOSX1_832 gnd vdd FILL
XFILL_0_NAND2X1_493 gnd vdd FILL
XFILL_0_OAI21X1_1253 gnd vdd FILL
XFILL_0_NAND2X1_482 gnd vdd FILL
XFILL_1_NAND2X1_653 gnd vdd FILL
XFILL_0_OAI21X1_1264 gnd vdd FILL
XFILL_0_OAI21X1_1275 gnd vdd FILL
XFILL_0_DFFPOSX1_843 gnd vdd FILL
XFILL_1_NAND2X1_675 gnd vdd FILL
XFILL_1_NAND2X1_697 gnd vdd FILL
XFILL_0_DFFPOSX1_876 gnd vdd FILL
XFILL_0_OAI21X1_1297 gnd vdd FILL
XFILL_0_OAI21X1_1286 gnd vdd FILL
XFILL_0_DFFPOSX1_854 gnd vdd FILL
XFILL_1_NAND2X1_686 gnd vdd FILL
XFILL_0_DFFPOSX1_865 gnd vdd FILL
XFILL_0_DFFPOSX1_887 gnd vdd FILL
XDFFPOSX1_1017 BUFX2_654/A CLKBUF1_3/Y OAI21X1_1594/Y gnd vdd DFFPOSX1
XDFFPOSX1_1006 BUFX2_661/A CLKBUF1_99/Y OAI21X1_1583/Y gnd vdd DFFPOSX1
XFILL_0_DFFPOSX1_898 gnd vdd FILL
XFILL_5_DFFPOSX1_480 gnd vdd FILL
XDFFPOSX1_1028 BUFX2_666/A CLKBUF1_51/Y OAI21X1_1605/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_219 gnd vdd FILL
XFILL_5_DFFPOSX1_491 gnd vdd FILL
XFILL_0_BUFX2_208 gnd vdd FILL
XFILL_0_AOI21X1_40 gnd vdd FILL
XFILL_0_AOI21X1_62 gnd vdd FILL
XFILL_0_AOI21X1_51 gnd vdd FILL
XFILL_2_DFFPOSX1_904 gnd vdd FILL
XFILL_2_DFFPOSX1_915 gnd vdd FILL
XFILL_2_DFFPOSX1_948 gnd vdd FILL
XFILL_2_DFFPOSX1_937 gnd vdd FILL
XFILL_2_OAI21X1_1369 gnd vdd FILL
XFILL_2_OAI21X1_1358 gnd vdd FILL
XFILL_2_DFFPOSX1_926 gnd vdd FILL
XFILL_2_DFFPOSX1_959 gnd vdd FILL
XFILL_3_XNOR2X1_17 gnd vdd FILL
XFILL_3_XNOR2X1_39 gnd vdd FILL
XFILL_0_BUFX2_742 gnd vdd FILL
XFILL_0_BUFX2_720 gnd vdd FILL
XDFFPOSX1_318 BUFX2_988/A CLKBUF1_7/Y OAI21X1_253/Y gnd vdd DFFPOSX1
XDFFPOSX1_307 BUFX2_976/A CLKBUF1_74/Y OAI21X1_231/Y gnd vdd DFFPOSX1
XDFFPOSX1_329 BUFX2_1000/A CLKBUF1_70/Y OAI21X1_275/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_731 gnd vdd FILL
XFILL_1_DFFPOSX1_505 gnd vdd FILL
XFILL_0_NOR2X1_60 gnd vdd FILL
XFILL_0_BUFX2_775 gnd vdd FILL
XFILL_0_BUFX2_753 gnd vdd FILL
XFILL_0_BUFX2_764 gnd vdd FILL
XFILL_0_NOR2X1_93 gnd vdd FILL
XFILL_1_DFFPOSX1_516 gnd vdd FILL
XFILL_1_DFFPOSX1_527 gnd vdd FILL
XFILL_0_NOR2X1_82 gnd vdd FILL
XFILL_1_DFFPOSX1_538 gnd vdd FILL
XFILL_0_NOR2X1_71 gnd vdd FILL
XFILL_0_BUFX2_797 gnd vdd FILL
XFILL_0_BUFX2_786 gnd vdd FILL
XFILL_1_DFFPOSX1_549 gnd vdd FILL
XFILL_6_DFFPOSX1_120 gnd vdd FILL
XFILL_3_DFFPOSX1_4 gnd vdd FILL
XFILL_37_2_1 gnd vdd FILL
XBUFX4_361 BUFX4_380/A gnd BUFX4_361/Y vdd BUFX4
XBUFX4_372 BUFX4_388/A gnd BUFX4_372/Y vdd BUFX4
XBUFX4_350 BUFX4_384/A gnd BUFX4_350/Y vdd BUFX4
XBUFX4_383 BUFX4_385/A gnd BUFX4_383/Y vdd BUFX4
XFILL_0_DFFPOSX1_117 gnd vdd FILL
XFILL_0_DFFPOSX1_106 gnd vdd FILL
XFILL_0_DFFPOSX1_128 gnd vdd FILL
XFILL_0_DFFPOSX1_139 gnd vdd FILL
XOAI21X1_905 INVX1_106/Y BUFX4_189/Y OAI21X1_905/C gnd OAI21X1_905/Y vdd OAI21X1
XOAI21X1_916 BUFX4_96/Y OAI21X1_7/A BUFX2_351/A gnd OAI21X1_917/C vdd OAI21X1
XOAI21X1_949 BUFX4_165/Y INVX1_129/Y OAI21X1_949/C gnd OAI21X1_949/Y vdd OAI21X1
XFILL_20_1_1 gnd vdd FILL
XOAI21X1_938 BUFX4_111/Y BUFX4_330/Y BUFX2_332/A gnd OAI21X1_939/C vdd OAI21X1
XOAI21X1_927 BUFX4_124/Y INVX1_118/Y OAI21X1_927/C gnd OAI21X1_927/Y vdd OAI21X1
XFILL_0_NAND2X1_4 gnd vdd FILL
XOAI21X1_1240 BUFX4_10/A BUFX4_386/Y BUFX2_133/A gnd OAI21X1_1241/C vdd OAI21X1
XFILL_21_17_1 gnd vdd FILL
XOAI21X1_1251 XNOR2X1_77/Y BUFX4_150/Y OAI21X1_1251/C gnd OAI21X1_1251/Y vdd OAI21X1
XDFFPOSX1_841 BUFX2_92/A CLKBUF1_95/Y OAI21X1_1156/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1460 gnd vdd FILL
XOAI21X1_1262 BUFX4_5/Y BUFX4_324/Y BUFX2_140/A gnd OAI21X1_1263/C vdd OAI21X1
XOAI21X1_1273 BUFX4_4/A OAI21X1_5/A BUFX2_144/A gnd OAI21X1_1274/C vdd OAI21X1
XDFFPOSX1_830 BUFX2_80/A CLKBUF1_52/Y OAI21X1_1141/Y gnd vdd DFFPOSX1
XDFFPOSX1_874 BUFX2_141/A CLKBUF1_74/Y OAI21X1_1213/Y gnd vdd DFFPOSX1
XOAI21X1_1295 BUFX4_99/Y BUFX4_381/Y BUFX2_155/A gnd OAI21X1_1296/C vdd OAI21X1
XFILL_0_OAI21X1_240 gnd vdd FILL
XFILL_1_OAI21X1_1471 gnd vdd FILL
XFILL_1_OAI21X1_1482 gnd vdd FILL
XDFFPOSX1_852 BUFX2_104/A CLKBUF1_68/Y OAI21X1_1172/Y gnd vdd DFFPOSX1
XOAI21X1_1284 XNOR2X1_80/Y OR2X2_20/B OAI21X1_1284/C gnd OAI21X1_1284/Y vdd OAI21X1
XFILL_1_OAI21X1_1493 gnd vdd FILL
XFILL_1_OAI21X1_411 gnd vdd FILL
XFILL_1_OAI21X1_400 gnd vdd FILL
XDFFPOSX1_863 BUFX2_116/A CLKBUF1_20/Y OAI21X1_1191/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_273 gnd vdd FILL
XFILL_0_OAI21X1_262 gnd vdd FILL
XFILL_0_OAI21X1_251 gnd vdd FILL
XDFFPOSX1_885 BUFX2_134/A CLKBUF1_50/Y OAI21X1_1245/Y gnd vdd DFFPOSX1
XDFFPOSX1_896 BUFX2_146/A CLKBUF1_60/Y OAI21X1_1277/Y gnd vdd DFFPOSX1
XINVX2_35 bundleStartMajId_i[11] gnd NOR3X1_8/A vdd INVX2
XFILL_2_OAI21X1_604 gnd vdd FILL
XINVX2_24 bundleStartMajId_i[32] gnd INVX2_24/Y vdd INVX2
XFILL_1_OAI21X1_422 gnd vdd FILL
XFILL_1_OAI21X1_444 gnd vdd FILL
XINVX2_13 bundleStartMajId_i[56] gnd INVX2_13/Y vdd INVX2
XFILL_1_OAI21X1_433 gnd vdd FILL
XFILL_0_OAI21X1_295 gnd vdd FILL
XINVX2_68 bundleAddress_i[46] gnd INVX2_68/Y vdd INVX2
XINVX2_57 bundleAddress_i[59] gnd INVX2_57/Y vdd INVX2
XFILL_1_OAI21X1_477 gnd vdd FILL
XFILL_1_OAI21X1_455 gnd vdd FILL
XINVX2_46 INVX2_46/A gnd INVX2_46/Y vdd INVX2
XINVX2_79 bundleAddress_i[23] gnd INVX2_79/Y vdd INVX2
XFILL_1_OAI21X1_466 gnd vdd FILL
XFILL_0_OAI21X1_284 gnd vdd FILL
XFILL_1_OAI21X1_499 gnd vdd FILL
XFILL_1_OAI21X1_488 gnd vdd FILL
XFILL_0_AOI21X1_9 gnd vdd FILL
XBUFX2_309 BUFX2_309/A gnd instr2_o[8] vdd BUFX2
XFILL_28_2_1 gnd vdd FILL
XFILL_3_2_1 gnd vdd FILL
XFILL_1_INVX4_24 gnd vdd FILL
XFILL_1_INVX4_13 gnd vdd FILL
XFILL_0_OAI21X1_1050 gnd vdd FILL
XFILL_1_BUFX4_203 gnd vdd FILL
XFILL_1_NAND2X1_450 gnd vdd FILL
XFILL_0_DFFPOSX1_640 gnd vdd FILL
XFILL_1_NAND2X1_472 gnd vdd FILL
XFILL_0_OAI21X1_1083 gnd vdd FILL
XFILL_1_NAND2X1_483 gnd vdd FILL
XFILL_1_NAND2X1_461 gnd vdd FILL
XFILL_0_DFFPOSX1_651 gnd vdd FILL
XFILL_0_OAI21X1_1061 gnd vdd FILL
XFILL_0_NAND2X1_290 gnd vdd FILL
XFILL_1_BUFX4_225 gnd vdd FILL
XFILL_1_BUFX4_236 gnd vdd FILL
XFILL_1_BUFX4_214 gnd vdd FILL
XFILL_0_OAI21X1_1072 gnd vdd FILL
XFILL_0_DFFPOSX1_662 gnd vdd FILL
XFILL_1_BUFX4_247 gnd vdd FILL
XFILL_1_BUFX4_269 gnd vdd FILL
XFILL_26_16_1 gnd vdd FILL
XFILL_0_OAI21X1_1094 gnd vdd FILL
XFILL_1_BUFX4_258 gnd vdd FILL
XFILL_0_DFFPOSX1_673 gnd vdd FILL
XFILL_0_DFFPOSX1_684 gnd vdd FILL
XFILL_0_DFFPOSX1_695 gnd vdd FILL
XFILL_11_1_1 gnd vdd FILL
XFILL_20_12_0 gnd vdd FILL
XFILL_0_DFFPOSX1_18 gnd vdd FILL
XFILL_0_DFFPOSX1_29 gnd vdd FILL
XFILL_2_XNOR2X1_7 gnd vdd FILL
XFILL_2_BUFX4_85 gnd vdd FILL
XFILL_2_DFFPOSX1_701 gnd vdd FILL
XBUFX2_821 BUFX2_821/A gnd tid1_o[14] vdd BUFX2
XBUFX2_810 BUFX2_810/A gnd tid1_o[24] vdd BUFX2
XFILL_19_2_1 gnd vdd FILL
XFILL_2_DFFPOSX1_712 gnd vdd FILL
XFILL_2_DFFPOSX1_723 gnd vdd FILL
XFILL_2_DFFPOSX1_756 gnd vdd FILL
XFILL_2_DFFPOSX1_745 gnd vdd FILL
XFILL_2_DFFPOSX1_734 gnd vdd FILL
XFILL_1_17_1 gnd vdd FILL
XBUFX2_832 NAND2X1_3/A gnd tid1_o[4] vdd BUFX2
XBUFX2_843 BUFX2_843/A gnd tid2_o[53] vdd BUFX2
XBUFX2_854 BUFX2_854/A gnd tid2_o[43] vdd BUFX2
XBUFX2_887 BUFX2_887/A gnd tid2_o[13] vdd BUFX2
XBUFX2_865 BUFX2_865/A gnd tid2_o[33] vdd BUFX2
XFILL_2_DFFPOSX1_789 gnd vdd FILL
XFILL_2_DFFPOSX1_778 gnd vdd FILL
XBUFX2_898 BUFX2_898/A gnd tid2_o[3] vdd BUFX2
XBUFX2_876 BUFX2_876/A gnd tid2_o[23] vdd BUFX2
XFILL_2_DFFPOSX1_767 gnd vdd FILL
XFILL_0_NOR2X1_216 gnd vdd FILL
XFILL_0_NOR2X1_205 gnd vdd FILL
XFILL_0_NOR2X1_227 gnd vdd FILL
XFILL_31_9_0 gnd vdd FILL
XFILL_12_4 gnd vdd FILL
XFILL_25_11_0 gnd vdd FILL
XFILL_3_CLKBUF1_7 gnd vdd FILL
XDFFPOSX1_104 BUFX2_811/A CLKBUF1_59/Y OAI21X1_1778/Y gnd vdd DFFPOSX1
XDFFPOSX1_126 BUFX2_796/A CLKBUF1_3/Y OAI21X1_1800/Y gnd vdd DFFPOSX1
XDFFPOSX1_115 BUFX2_784/A CLKBUF1_39/Y OAI21X1_1789/Y gnd vdd DFFPOSX1
XDFFPOSX1_137 BUFX2_808/A CLKBUF1_39/Y OAI21X1_1811/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_313 gnd vdd FILL
XFILL_1_DFFPOSX1_302 gnd vdd FILL
XFILL_0_BUFX2_550 gnd vdd FILL
XDFFPOSX1_148 BUFX2_820/A CLKBUF1_7/Y OAI21X1_1822/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_346 gnd vdd FILL
XFILL_1_DFFPOSX1_335 gnd vdd FILL
XFILL_0_BUFX2_572 gnd vdd FILL
XFILL_0_BUFX2_561 gnd vdd FILL
XDFFPOSX1_159 NAND2X1_3/A CLKBUF1_51/Y OAI21X1_3/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_583 gnd vdd FILL
XFILL_1_DFFPOSX1_324 gnd vdd FILL
XFILL_1_DFFPOSX1_357 gnd vdd FILL
XFILL_1_DFFPOSX1_368 gnd vdd FILL
XFILL_1_DFFPOSX1_379 gnd vdd FILL
XFILL_0_BUFX2_594 gnd vdd FILL
XNAND2X1_207 BUFX2_485/A BUFX4_194/Y gnd OAI21X1_452/C vdd NAND2X1
XNAND2X1_218 bundleStartMajId_i[22] NOR2X1_35/Y gnd OAI21X1_462/A vdd NAND2X1
XNAND2X1_229 BUFX2_499/A BUFX4_182/Y gnd OAI21X1_471/C vdd NAND2X1
XFILL_4_DFFPOSX1_806 gnd vdd FILL
XFILL_4_DFFPOSX1_817 gnd vdd FILL
XFILL_4_DFFPOSX1_828 gnd vdd FILL
XFILL_4_DFFPOSX1_839 gnd vdd FILL
XFILL_6_16_1 gnd vdd FILL
XBUFX4_191 BUFX4_26/Y gnd BUFX4_191/Y vdd BUFX4
XBUFX4_180 BUFX4_24/Y gnd BUFX4_180/Y vdd BUFX4
XFILL_4_CLKBUF1_40 gnd vdd FILL
XFILL_4_CLKBUF1_51 gnd vdd FILL
XFILL_0_INVX1_91 gnd vdd FILL
XFILL_0_BUFX2_11 gnd vdd FILL
XFILL_4_CLKBUF1_73 gnd vdd FILL
XFILL_0_INVX1_80 gnd vdd FILL
XFILL_4_CLKBUF1_84 gnd vdd FILL
XFILL_0_12_0 gnd vdd FILL
XFILL_0_BUFX2_22 gnd vdd FILL
XFILL_0_BUFX2_44 gnd vdd FILL
XFILL_0_BUFX2_33 gnd vdd FILL
XFILL_0_BUFX2_77 gnd vdd FILL
XFILL_0_BUFX2_88 gnd vdd FILL
XFILL_0_BUFX2_66 gnd vdd FILL
XFILL_22_9_0 gnd vdd FILL
XFILL_0_BUFX2_55 gnd vdd FILL
XFILL_1_NOR2X1_36 gnd vdd FILL
XFILL_1_BUFX2_707 gnd vdd FILL
XFILL_1_BUFX2_718 gnd vdd FILL
XFILL_1_NOR2X1_14 gnd vdd FILL
XFILL_0_BUFX2_99 gnd vdd FILL
XOAI21X1_702 BUFX4_145/Y BUFX4_63/Y BUFX2_592/A gnd OAI21X1_703/C vdd OAI21X1
XFILL_1_NOR2X1_47 gnd vdd FILL
XOAI21X1_713 OR2X2_5/Y INVX1_36/A OAI21X1_713/C gnd OAI21X1_715/A vdd OAI21X1
XOAI21X1_724 OAI21X1_724/A BUFX4_300/Y OAI21X1_724/C gnd OAI21X1_724/Y vdd OAI21X1
XFILL_1_NOR2X1_69 gnd vdd FILL
XFILL_1_NOR2X1_58 gnd vdd FILL
XFILL_3_DFFPOSX1_418 gnd vdd FILL
XFILL_3_DFFPOSX1_407 gnd vdd FILL
XOAI21X1_757 INVX1_41/Y OAI21X1_757/B OAI21X1_757/C gnd OAI21X1_757/Y vdd OAI21X1
XOAI21X1_746 AOI21X1_33/Y NOR3X1_7/Y BUFX4_287/Y gnd OAI21X1_747/C vdd OAI21X1
XOAI21X1_735 BUFX4_174/Y BUFX4_79/Y BUFX2_604/A gnd OAI21X1_736/C vdd OAI21X1
XOAI21X1_768 BUFX4_142/Y BUFX4_37/Y BUFX2_618/A gnd OAI21X1_769/C vdd OAI21X1
XOAI21X1_779 NOR2X1_114/B NOR3X1_3/A INVX4_21/Y gnd OAI21X1_780/C vdd OAI21X1
XFILL_3_DFFPOSX1_429 gnd vdd FILL
XOAI21X1_1081 BUFX4_342/Y INVX2_81/Y NAND2X1_447/Y gnd OAI21X1_1081/Y vdd OAI21X1
XOAI21X1_1070 BUFX4_324/Y INVX4_40/Y NAND2X1_436/Y gnd OAI21X1_1070/Y vdd OAI21X1
XDFFPOSX1_660 BUFX2_297/A CLKBUF1_42/Y OAI21X1_888/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1290 gnd vdd FILL
XDFFPOSX1_693 BUFX2_330/A CLKBUF1_54/Y OAI21X1_935/Y gnd vdd DFFPOSX1
XDFFPOSX1_671 BUFX2_309/A CLKBUF1_10/Y OAI21X1_899/Y gnd vdd DFFPOSX1
XOAI21X1_1092 BUFX4_343/Y INVX2_88/Y NAND2X1_458/Y gnd OAI21X1_1092/Y vdd OAI21X1
XDFFPOSX1_682 BUFX2_337/A CLKBUF1_56/Y OAI21X1_913/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_880 gnd vdd FILL
XNAND2X1_730 BUFX2_784/A BUFX4_368/Y gnd NAND2X1_730/Y vdd NAND2X1
XFILL_1_OAI21X1_252 gnd vdd FILL
XFILL_1_OAI21X1_230 gnd vdd FILL
XFILL_1_OAI21X1_241 gnd vdd FILL
XFILL_1_DFFPOSX1_891 gnd vdd FILL
XFILL_0_NOR2X1_2 gnd vdd FILL
XFILL_2_OAI21X1_412 gnd vdd FILL
XFILL_2_OAI21X1_401 gnd vdd FILL
XNAND2X1_741 BUFX2_796/A BUFX4_363/Y gnd NAND2X1_741/Y vdd NAND2X1
XNAND2X1_752 BUFX2_808/A BUFX4_329/Y gnd NAND2X1_752/Y vdd NAND2X1
XNAND2X1_763 BUFX2_820/A BUFX4_377/Y gnd NAND2X1_763/Y vdd NAND2X1
XFILL_1_OAI21X1_296 gnd vdd FILL
XFILL_1_OAI21X1_274 gnd vdd FILL
XFILL_1_OAI21X1_263 gnd vdd FILL
XFILL_2_OAI21X1_434 gnd vdd FILL
XFILL_2_OAI21X1_467 gnd vdd FILL
XFILL_1_OAI21X1_285 gnd vdd FILL
XFILL_5_11_0 gnd vdd FILL
XFILL_2_XNOR2X1_14 gnd vdd FILL
XBUFX2_106 BUFX2_106/A gnd addr2_o[17] vdd BUFX2
XFILL_2_XNOR2X1_36 gnd vdd FILL
XFILL_2_XNOR2X1_25 gnd vdd FILL
XFILL_2_XNOR2X1_47 gnd vdd FILL
XBUFX2_117 BUFX2_117/A gnd addr2_o[7] vdd BUFX2
XBUFX2_139 BUFX2_139/A gnd addr3_o[45] vdd BUFX2
XFILL_2_XNOR2X1_58 gnd vdd FILL
XFILL_2_XNOR2X1_69 gnd vdd FILL
XBUFX2_128 BUFX2_128/A gnd addr2_o[54] vdd BUFX2
XFILL_13_9_0 gnd vdd FILL
XFILL_1_NAND2X1_291 gnd vdd FILL
XFILL_2_DFFPOSX1_1 gnd vdd FILL
XFILL_0_DFFPOSX1_470 gnd vdd FILL
XFILL_0_DFFPOSX1_481 gnd vdd FILL
XFILL_0_DFFPOSX1_492 gnd vdd FILL
XBUFX2_1009 BUFX2_1009/A gnd tid4_o[18] vdd BUFX2
XFILL_3_DFFPOSX1_941 gnd vdd FILL
XFILL_3_DFFPOSX1_930 gnd vdd FILL
XFILL_3_DFFPOSX1_952 gnd vdd FILL
XFILL_3_DFFPOSX1_963 gnd vdd FILL
XFILL_3_DFFPOSX1_974 gnd vdd FILL
XFILL_3_DFFPOSX1_985 gnd vdd FILL
XFILL_3_DFFPOSX1_996 gnd vdd FILL
XFILL_1_DFFPOSX1_19 gnd vdd FILL
XBUFX4_20 BUFX4_26/A gnd BUFX4_20/Y vdd BUFX4
XBUFX4_42 BUFX4_75/A gnd BUFX4_42/Y vdd BUFX4
XBUFX4_53 BUFX4_59/A gnd BUFX4_53/Y vdd BUFX4
XBUFX4_31 BUFX4_79/A gnd BUFX4_31/Y vdd BUFX4
XFILL_2_OAI21X1_990 gnd vdd FILL
XBUFX4_75 BUFX4_75/A gnd BUFX4_75/Y vdd BUFX4
XBUFX4_64 BUFX4_64/A gnd BUFX4_64/Y vdd BUFX4
XBUFX4_86 clock_i gnd BUFX4_86/Y vdd BUFX4
XFILL_0_OAI21X1_1808 gnd vdd FILL
XBUFX4_97 BUFX4_4/A gnd BUFX4_97/Y vdd BUFX4
XFILL_2_DFFPOSX1_520 gnd vdd FILL
XFILL_2_DFFPOSX1_531 gnd vdd FILL
XFILL_11_17_0 gnd vdd FILL
XFILL_0_OAI21X1_1819 gnd vdd FILL
XBUFX2_651 BUFX2_651/A gnd pid1_o[21] vdd BUFX2
XFILL_34_0_1 gnd vdd FILL
XFILL_2_DFFPOSX1_542 gnd vdd FILL
XBUFX2_662 BUFX2_662/A gnd pid1_o[11] vdd BUFX2
XBUFX2_640 BUFX2_640/A gnd majID4_o[4] vdd BUFX2
XFILL_2_DFFPOSX1_564 gnd vdd FILL
XBUFX2_673 BUFX2_673/A gnd pid1_o[1] vdd BUFX2
XFILL_2_DFFPOSX1_553 gnd vdd FILL
XBUFX2_695 BUFX2_695/A gnd pid2_o[10] vdd BUFX2
XBUFX2_684 BUFX2_684/A gnd pid2_o[20] vdd BUFX2
XFILL_2_DFFPOSX1_575 gnd vdd FILL
XFILL_2_DFFPOSX1_586 gnd vdd FILL
XFILL_2_DFFPOSX1_597 gnd vdd FILL
XFILL_10_1 gnd vdd FILL
XOR2X2_12 OR2X2_12/A bundleStartMajId_i[7] gnd OR2X2_12/Y vdd OR2X2
XFILL_1_DFFPOSX1_121 gnd vdd FILL
XFILL_2_AOI21X1_14 gnd vdd FILL
XOR2X2_5 OR2X2_5/A OR2X2_5/B gnd OR2X2_5/Y vdd OR2X2
XFILL_1_DFFPOSX1_110 gnd vdd FILL
XINVX2_180 bundleTid_i[29] gnd INVX2_180/Y vdd INVX2
XFILL_0_BUFX2_380 gnd vdd FILL
XINVX2_191 bundleTid_i[18] gnd INVX2_191/Y vdd INVX2
XFILL_1_DFFPOSX1_154 gnd vdd FILL
XFILL_1_DFFPOSX1_143 gnd vdd FILL
XFILL_0_BUFX2_391 gnd vdd FILL
XFILL_1_DFFPOSX1_165 gnd vdd FILL
XFILL_1_DFFPOSX1_132 gnd vdd FILL
XFILL_1_DFFPOSX1_198 gnd vdd FILL
XFILL_1_DFFPOSX1_176 gnd vdd FILL
XFILL_1_DFFPOSX1_187 gnd vdd FILL
XXNOR2X1_7 XNOR2X1_7/A bundleStartMajId_i[42] gnd XNOR2X1_7/Y vdd XNOR2X1
XFILL_4_DFFPOSX1_603 gnd vdd FILL
XFILL_4_DFFPOSX1_636 gnd vdd FILL
XFILL_16_16_0 gnd vdd FILL
XFILL_4_DFFPOSX1_625 gnd vdd FILL
XFILL_4_DFFPOSX1_614 gnd vdd FILL
XFILL_4_DFFPOSX1_647 gnd vdd FILL
XFILL_4_DFFPOSX1_658 gnd vdd FILL
XFILL_4_DFFPOSX1_669 gnd vdd FILL
XFILL_25_0_1 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XFILL_1_BUFX2_504 gnd vdd FILL
XFILL_1_BUFX2_515 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XFILL_1_BUFX2_526 gnd vdd FILL
XFILL_1_BUFX2_559 gnd vdd FILL
XOAI21X1_510 INVX1_24/A NOR2X1_59/B OAI21X1_510/C gnd OAI21X1_512/A vdd OAI21X1
XFILL_1_BUFX2_548 gnd vdd FILL
XOAI21X1_532 NOR2X1_104/A INVX4_30/Y OAI21X1_532/C gnd OAI21X1_534/A vdd OAI21X1
XOAI21X1_521 OAI21X1_521/A BUFX4_163/Y OAI21X1_521/C gnd OAI21X1_521/Y vdd OAI21X1
XFILL_3_DFFPOSX1_237 gnd vdd FILL
XFILL_3_DFFPOSX1_215 gnd vdd FILL
XOAI21X1_554 OR2X2_5/Y OR2X2_10/B OAI21X1_554/C gnd OAI21X1_556/A vdd OAI21X1
XOAI21X1_543 XNOR2X1_27/Y BUFX4_167/Y OAI21X1_543/C gnd OAI21X1_543/Y vdd OAI21X1
XFILL_3_DFFPOSX1_226 gnd vdd FILL
XFILL_3_DFFPOSX1_204 gnd vdd FILL
XOAI21X1_565 XNOR2X1_31/Y BUFX4_130/Y OAI21X1_565/C gnd OAI21X1_565/Y vdd OAI21X1
XFILL_3_DFFPOSX1_248 gnd vdd FILL
XFILL_3_DFFPOSX1_259 gnd vdd FILL
XOAI21X1_576 INVX1_28/Y INVX8_6/A NAND3X1_16/Y gnd OAI21X1_576/Y vdd OAI21X1
XOAI21X1_598 OR2X2_9/Y NOR3X1_6/B OAI21X1_598/C gnd OAI21X1_600/A vdd OAI21X1
XOAI21X1_587 OR2X2_9/A INVX4_15/Y INVX1_2/Y gnd OAI21X1_588/C vdd OAI21X1
XDFFPOSX1_490 BUFX2_577/A CLKBUF1_46/Y OAI21X1_517/Y gnd vdd DFFPOSX1
XFILL_2_OAI21X1_220 gnd vdd FILL
XFILL_8_1_1 gnd vdd FILL
XFILL_34_17_0 gnd vdd FILL
XFILL_2_OAI21X1_253 gnd vdd FILL
XNAND2X1_560 BUFX2_108/A BUFX4_203/Y gnd NAND2X1_560/Y vdd NAND2X1
XNAND2X1_571 bundleAddress_i[13] bundleAddress_i[12] gnd NAND2X1_571/Y vdd NAND2X1
XNAND2X1_593 INVX4_47/A NOR2X1_180/Y gnd INVX1_201/A vdd NAND2X1
XNAND2X1_582 BUFX2_119/A BUFX4_187/Y gnd NAND2X1_582/Y vdd NAND2X1
XFILL_16_0_1 gnd vdd FILL
XFILL_5_DFFPOSX1_309 gnd vdd FILL
XFILL_1_DFFPOSX1_1017 gnd vdd FILL
XFILL_1_DFFPOSX1_1006 gnd vdd FILL
XFILL_1_DFFPOSX1_1028 gnd vdd FILL
XOAI21X1_1806 BUFX4_320/Y INVX2_178/Y NAND2X1_747/Y gnd OAI21X1_1806/Y vdd OAI21X1
XOAI21X1_1828 BUFX4_352/Y INVX2_200/Y NAND2X1_769/Y gnd OAI21X1_1828/Y vdd OAI21X1
XOAI21X1_1817 BUFX4_313/Y INVX2_189/Y NAND2X1_758/Y gnd OAI21X1_1817/Y vdd OAI21X1
XFILL_3_DFFPOSX1_771 gnd vdd FILL
XFILL_3_DFFPOSX1_760 gnd vdd FILL
XFILL_3_DFFPOSX1_782 gnd vdd FILL
XFILL_3_CLKBUF1_70 gnd vdd FILL
XFILL_0_OAI21X1_839 gnd vdd FILL
XFILL_0_OAI21X1_828 gnd vdd FILL
XFILL_0_OAI21X1_806 gnd vdd FILL
XFILL_3_DFFPOSX1_793 gnd vdd FILL
XFILL_0_OAI21X1_817 gnd vdd FILL
XFILL_3_CLKBUF1_81 gnd vdd FILL
XFILL_3_CLKBUF1_92 gnd vdd FILL
XFILL_36_8_0 gnd vdd FILL
XFILL_0_OAI21X1_1616 gnd vdd FILL
XFILL_0_OAI21X1_1605 gnd vdd FILL
XFILL_0_OAI21X1_1649 gnd vdd FILL
XBUFX2_481 BUFX2_481/A gnd majID2_o[33] vdd BUFX2
XFILL_0_OAI21X1_1627 gnd vdd FILL
XBUFX2_470 BUFX2_470/A gnd majID2_o[43] vdd BUFX2
XFILL_2_DFFPOSX1_350 gnd vdd FILL
XFILL_0_OAI21X1_1638 gnd vdd FILL
XFILL_2_DFFPOSX1_361 gnd vdd FILL
XFILL_2_DFFPOSX1_372 gnd vdd FILL
XFILL_2_DFFPOSX1_383 gnd vdd FILL
XFILL_2_DFFPOSX1_394 gnd vdd FILL
XBUFX2_492 BUFX2_492/A gnd majID2_o[23] vdd BUFX2
XFILL_5_DFFPOSX1_821 gnd vdd FILL
XFILL_5_DFFPOSX1_810 gnd vdd FILL
XFILL_5_DFFPOSX1_832 gnd vdd FILL
XFILL_5_DFFPOSX1_854 gnd vdd FILL
XFILL_5_DFFPOSX1_843 gnd vdd FILL
XFILL_5_DFFPOSX1_887 gnd vdd FILL
XFILL_5_DFFPOSX1_876 gnd vdd FILL
XFILL_5_DFFPOSX1_898 gnd vdd FILL
XFILL_1_XNOR2X1_22 gnd vdd FILL
XFILL_5_DFFPOSX1_865 gnd vdd FILL
XFILL_1_XNOR2X1_11 gnd vdd FILL
XFILL_1_XNOR2X1_55 gnd vdd FILL
XFILL_1_XNOR2X1_33 gnd vdd FILL
XFILL_1_XNOR2X1_44 gnd vdd FILL
XFILL_1_XNOR2X1_77 gnd vdd FILL
XFILL_1_XNOR2X1_66 gnd vdd FILL
XFILL_1_XNOR2X1_88 gnd vdd FILL
XFILL_1_XNOR2X1_99 gnd vdd FILL
XFILL_4_DFFPOSX1_400 gnd vdd FILL
XFILL_4_DFFPOSX1_411 gnd vdd FILL
XFILL_4_DFFPOSX1_422 gnd vdd FILL
XFILL_4_DFFPOSX1_433 gnd vdd FILL
XFILL_4_DFFPOSX1_455 gnd vdd FILL
XFILL_4_DFFPOSX1_444 gnd vdd FILL
XFILL_4_DFFPOSX1_477 gnd vdd FILL
XFILL_4_DFFPOSX1_466 gnd vdd FILL
XFILL_4_DFFPOSX1_488 gnd vdd FILL
XFILL_27_8_0 gnd vdd FILL
XFILL_4_DFFPOSX1_499 gnd vdd FILL
XFILL_2_8_0 gnd vdd FILL
XFILL_1_BUFX2_301 gnd vdd FILL
XFILL_1_BUFX2_323 gnd vdd FILL
XFILL_1_BUFX2_312 gnd vdd FILL
XOAI21X1_340 BUFX4_358/Y INVX4_5/Y NAND2X1_84/Y gnd OAI21X1_340/Y vdd OAI21X1
XFILL_10_7_0 gnd vdd FILL
XFILL_1_BUFX2_356 gnd vdd FILL
XFILL_1_BUFX2_367 gnd vdd FILL
XFILL_23_14_1 gnd vdd FILL
XAND2X2_7 AND2X2_7/A AND2X2_7/B gnd AND2X2_7/Y vdd AND2X2
XOAI21X1_373 BUFX4_345/Y INVX2_30/Y OAI21X1_373/C gnd OAI21X1_373/Y vdd OAI21X1
XOAI21X1_351 BUFX4_337/Y INVX4_9/Y NAND2X1_95/Y gnd OAI21X1_351/Y vdd OAI21X1
XOAI21X1_362 BUFX4_373/Y INVX1_2/Y OAI21X1_362/C gnd OAI21X1_362/Y vdd OAI21X1
XOAI21X1_384 BUFX4_319/Y INVX2_37/Y OAI21X1_384/C gnd OAI21X1_384/Y vdd OAI21X1
XOAI21X1_395 INVX4_1/Y INVX1_24/A OAI21X1_395/C gnd OAI21X1_396/A vdd OAI21X1
XFILL_6_DFFPOSX1_516 gnd vdd FILL
XFILL_6_DFFPOSX1_527 gnd vdd FILL
XFILL_6_DFFPOSX1_505 gnd vdd FILL
XFILL_6_DFFPOSX1_538 gnd vdd FILL
XFILL_6_DFFPOSX1_549 gnd vdd FILL
XNAND2X1_390 BUFX2_306/A BUFX4_184/Y gnd OAI21X1_896/C vdd NAND2X1
XFILL_0_NAND2X1_108 gnd vdd FILL
XFILL_0_NAND2X1_119 gnd vdd FILL
XFILL_18_8_0 gnd vdd FILL
XFILL_0_INVX1_122 gnd vdd FILL
XFILL_0_INVX1_100 gnd vdd FILL
XFILL_0_INVX1_111 gnd vdd FILL
XFILL_0_INVX1_144 gnd vdd FILL
XFILL_0_INVX1_133 gnd vdd FILL
XFILL_1_AOI21X1_22 gnd vdd FILL
XFILL_1_AOI21X1_11 gnd vdd FILL
XFILL_1_AOI21X1_33 gnd vdd FILL
XFILL_0_INVX1_155 gnd vdd FILL
XFILL_0_INVX1_166 gnd vdd FILL
XFILL_0_INVX1_177 gnd vdd FILL
XFILL_1_AOI21X1_66 gnd vdd FILL
XFILL_1_AOI21X1_44 gnd vdd FILL
XFILL_0_INVX1_188 gnd vdd FILL
XFILL_1_AOI21X1_55 gnd vdd FILL
XFILL_5_DFFPOSX1_117 gnd vdd FILL
XFILL_28_13_1 gnd vdd FILL
XFILL_5_DFFPOSX1_106 gnd vdd FILL
XFILL_0_INVX1_199 gnd vdd FILL
XFILL_5_DFFPOSX1_139 gnd vdd FILL
XFILL_5_DFFPOSX1_128 gnd vdd FILL
XFILL_1_BUFX2_890 gnd vdd FILL
XOAI21X1_1614 INVX2_117/Y BUFX4_203/Y NAND2X1_682/Y gnd DFFPOSX1_4/D vdd OAI21X1
XOAI21X1_1603 BUFX4_359/Y INVX2_139/Y NAND2X1_672/Y gnd OAI21X1_1603/Y vdd OAI21X1
XFILL_1_OAI21X1_1801 gnd vdd FILL
XFILL_1_OAI21X1_1812 gnd vdd FILL
XOAI21X1_1647 BUFX4_172/Y INVX2_117/Y OAI21X1_1647/C gnd DFFPOSX1_36/D vdd OAI21X1
XOAI21X1_1636 INVX2_139/Y BUFX4_223/Y NAND2X1_704/Y gnd DFFPOSX1_26/D vdd OAI21X1
XFILL_1_OAI21X1_1823 gnd vdd FILL
XOAI21X1_1625 INVX2_128/Y BUFX4_211/Y NAND2X1_693/Y gnd DFFPOSX1_15/D vdd OAI21X1
XOAI21X1_1669 BUFX4_151/Y INVX2_128/Y OAI21X1_1669/C gnd DFFPOSX1_47/D vdd OAI21X1
XFILL_0_OAI21X1_614 gnd vdd FILL
XFILL_3_DFFPOSX1_590 gnd vdd FILL
XFILL_0_OAI21X1_603 gnd vdd FILL
XOAI21X1_1658 BUFX4_7/A OAI21X1_6/A BUFX2_741/A gnd OAI21X1_1659/C vdd OAI21X1
XFILL_0_OAI21X1_647 gnd vdd FILL
XFILL_1_OAI21X1_807 gnd vdd FILL
XFILL_0_OAI21X1_636 gnd vdd FILL
XFILL_0_OAI21X1_625 gnd vdd FILL
XFILL_1_OAI21X1_818 gnd vdd FILL
XFILL_1_OAI21X1_829 gnd vdd FILL
XFILL_0_OAI21X1_658 gnd vdd FILL
XFILL_0_OAI21X1_669 gnd vdd FILL
XFILL_1_AND2X2_26 gnd vdd FILL
XFILL_1_AND2X2_15 gnd vdd FILL
XFILL_0_NAND2X1_620 gnd vdd FILL
XFILL_3_14_1 gnd vdd FILL
XFILL_0_OAI21X1_1413 gnd vdd FILL
XFILL_0_OAI21X1_1402 gnd vdd FILL
XFILL_0_NAND2X1_653 gnd vdd FILL
XFILL_0_OAI21X1_1424 gnd vdd FILL
XFILL_0_NAND2X1_642 gnd vdd FILL
XFILL_0_NAND2X1_631 gnd vdd FILL
XFILL_2_DFFPOSX1_191 gnd vdd FILL
XFILL_2_DFFPOSX1_180 gnd vdd FILL
XFILL_0_NAND2X1_664 gnd vdd FILL
XFILL_0_OAI21X1_1435 gnd vdd FILL
XFILL_0_OAI21X1_1457 gnd vdd FILL
XFILL_0_NAND2X1_686 gnd vdd FILL
XFILL_0_OAI21X1_1446 gnd vdd FILL
XFILL_0_NAND2X1_675 gnd vdd FILL
XFILL_0_NAND2X1_697 gnd vdd FILL
XFILL_0_OAI21X1_1479 gnd vdd FILL
XFILL_0_OAI21X1_1468 gnd vdd FILL
XFILL_4_DFFPOSX1_8 gnd vdd FILL
XFILL_5_DFFPOSX1_662 gnd vdd FILL
XFILL_5_DFFPOSX1_640 gnd vdd FILL
XFILL_5_DFFPOSX1_651 gnd vdd FILL
XFILL_5_DFFPOSX1_673 gnd vdd FILL
XFILL_5_DFFPOSX1_695 gnd vdd FILL
XFILL_5_DFFPOSX1_684 gnd vdd FILL
XFILL_8_13_1 gnd vdd FILL
XFILL_4_DFFPOSX1_230 gnd vdd FILL
XFILL_4_DFFPOSX1_252 gnd vdd FILL
XFILL_4_DFFPOSX1_263 gnd vdd FILL
XFILL_4_DFFPOSX1_241 gnd vdd FILL
XFILL_4_DFFPOSX1_296 gnd vdd FILL
XFILL_4_DFFPOSX1_285 gnd vdd FILL
XFILL_4_DFFPOSX1_274 gnd vdd FILL
XFILL_1_BUFX2_120 gnd vdd FILL
XFILL_1_BUFX2_153 gnd vdd FILL
XFILL_1_BUFX2_175 gnd vdd FILL
XFILL_1_BUFX2_164 gnd vdd FILL
XFILL_0_BUFX2_924 gnd vdd FILL
XFILL_1_BUFX2_197 gnd vdd FILL
XOAI21X1_181 BUFX4_143/Y INVX2_200/Y OAI21X1_181/C gnd OAI21X1_181/Y vdd OAI21X1
XFILL_1_OAI21X1_1108 gnd vdd FILL
XINVX1_201 INVX1_201/A gnd INVX1_201/Y vdd INVX1
XFILL_0_BUFX2_913 gnd vdd FILL
XFILL_0_BUFX2_902 gnd vdd FILL
XFILL_1_OAI21X1_1119 gnd vdd FILL
XOAI21X1_170 BUFX4_96/Y BUFX4_330/Y BUFX2_949/A gnd OAI21X1_171/C vdd OAI21X1
XOAI21X1_192 BUFX4_109/Y BUFX4_354/Y BUFX2_962/A gnd OAI21X1_193/C vdd OAI21X1
XFILL_0_BUFX2_957 gnd vdd FILL
XINVX1_212 INVX1_212/A gnd INVX1_212/Y vdd INVX1
XFILL_0_BUFX2_935 gnd vdd FILL
XINVX1_223 INVX1_223/A gnd INVX1_223/Y vdd INVX1
XFILL_0_BUFX2_946 gnd vdd FILL
XFILL_1_DFFPOSX1_709 gnd vdd FILL
XFILL_0_BUFX2_968 gnd vdd FILL
XFILL_0_BUFX2_979 gnd vdd FILL
XFILL_6_DFFPOSX1_302 gnd vdd FILL
XNAND2X1_23 BUFX2_848/A BUFX4_216/Y gnd OAI21X1_23/C vdd NAND2X1
XNAND2X1_34 BUFX2_860/A BUFX4_191/Y gnd OAI21X1_34/C vdd NAND2X1
XNAND2X1_12 BUFX2_875/A BUFX4_197/Y gnd OAI21X1_12/C vdd NAND2X1
XNAND2X1_56 BUFX2_884/A BUFX4_191/Y gnd OAI21X1_56/C vdd NAND2X1
XNAND2X1_45 BUFX2_872/A BUFX4_200/Y gnd OAI21X1_45/C vdd NAND2X1
XFILL_2_INVX8_2 gnd vdd FILL
XNAND2X1_67 BUFX2_896/A OAI21X1_9/B gnd OAI21X1_67/C vdd NAND2X1
XFILL_0_XNOR2X1_30 gnd vdd FILL
XFILL_0_XNOR2X1_63 gnd vdd FILL
XFILL_0_XNOR2X1_52 gnd vdd FILL
XNAND2X1_89 BUFX2_402/A BUFX4_387/Y gnd NAND2X1_89/Y vdd NAND2X1
XFILL_0_XNOR2X1_41 gnd vdd FILL
XNAND2X1_78 BUFX2_449/A BUFX4_355/Y gnd NAND2X1_78/Y vdd NAND2X1
XFILL_0_XNOR2X1_74 gnd vdd FILL
XFILL_0_XNOR2X1_85 gnd vdd FILL
XFILL_0_XNOR2X1_96 gnd vdd FILL
XFILL_33_6_0 gnd vdd FILL
XFILL_0_NOR3X1_17 gnd vdd FILL
XFILL_0_BUFX4_250 gnd vdd FILL
XOAI21X1_1422 NOR2X1_183/A INVX2_108/Y OAI21X1_1422/C gnd OAI21X1_1424/A vdd OAI21X1
XOAI21X1_1400 BUFX4_151/Y BUFX4_75/A BUFX2_249/A gnd OAI21X1_1401/C vdd OAI21X1
XOAI21X1_1411 BUFX4_145/Y BUFX4_72/Y BUFX2_256/A gnd OAI21X1_1412/C vdd OAI21X1
XFILL_1_OAI21X1_1642 gnd vdd FILL
XFILL_1_OAI21X1_1631 gnd vdd FILL
XOAI21X1_1433 OAI21X1_1433/A BUFX4_291/Y OAI21X1_1433/C gnd OAI21X1_1433/Y vdd OAI21X1
XFILL_0_BUFX4_272 gnd vdd FILL
XOAI21X1_1466 OAI21X1_1466/A BUFX4_292/Y OAI21X1_1466/C gnd OAI21X1_1466/Y vdd OAI21X1
XFILL_0_BUFX4_283 gnd vdd FILL
XFILL_0_BUFX4_294 gnd vdd FILL
XOAI21X1_1455 XNOR2X1_96/Y INVX8_2/A OAI21X1_1455/C gnd OAI21X1_1455/Y vdd OAI21X1
XOAI21X1_1444 BUFX4_124/Y BUFX4_27/Y BUFX2_206/A gnd OAI21X1_1445/C vdd OAI21X1
XFILL_0_BUFX4_261 gnd vdd FILL
XFILL_1_OAI21X1_1620 gnd vdd FILL
XFILL_1_OAI21X1_1675 gnd vdd FILL
XFILL_1_OAI21X1_1653 gnd vdd FILL
XFILL_1_OAI21X1_1664 gnd vdd FILL
XOAI21X1_1477 INVX2_99/Y XNOR2X1_99/A OAI21X1_1477/C gnd OAI21X1_1479/A vdd OAI21X1
XFILL_4_NOR3X1_16 gnd vdd FILL
XFILL_0_OAI21X1_411 gnd vdd FILL
XFILL_0_OAI21X1_422 gnd vdd FILL
XFILL_0_OAI21X1_400 gnd vdd FILL
XOAI21X1_1488 OAI21X1_1488/A BUFX4_294/Y OAI21X1_1488/C gnd OAI21X1_1488/Y vdd OAI21X1
XOAI21X1_1499 NAND2X1_638/Y BUFX4_294/Y OAI21X1_1499/C gnd OAI21X1_1499/Y vdd OAI21X1
XFILL_1_OAI21X1_626 gnd vdd FILL
XFILL_1_OAI21X1_1686 gnd vdd FILL
XFILL_1_OAI21X1_1697 gnd vdd FILL
XFILL_0_OAI21X1_455 gnd vdd FILL
XFILL_1_NOR2X1_209 gnd vdd FILL
XFILL_1_OAI21X1_615 gnd vdd FILL
XFILL_1_OAI21X1_604 gnd vdd FILL
XFILL_0_OAI21X1_444 gnd vdd FILL
XFILL_0_OAI21X1_433 gnd vdd FILL
XFILL_1_OAI21X1_648 gnd vdd FILL
XFILL_0_OAI21X1_477 gnd vdd FILL
XFILL_1_OAI21X1_659 gnd vdd FILL
XFILL_0_OAI21X1_488 gnd vdd FILL
XFILL_19_18_1 gnd vdd FILL
XFILL_2_OAI21X1_819 gnd vdd FILL
XFILL_1_OAI21X1_637 gnd vdd FILL
XFILL_0_OAI21X1_466 gnd vdd FILL
XFILL_6_DFFPOSX1_880 gnd vdd FILL
XFILL_3_DFFPOSX1_1030 gnd vdd FILL
XFILL_0_OAI21X1_499 gnd vdd FILL
XFILL_6_DFFPOSX1_891 gnd vdd FILL
XFILL_13_14_0 gnd vdd FILL
XFILL_0_OAI21X1_1232 gnd vdd FILL
XFILL_0_OAI21X1_1221 gnd vdd FILL
XFILL_0_NAND2X1_450 gnd vdd FILL
XFILL_0_OAI21X1_1210 gnd vdd FILL
XFILL_0_NAND2X1_461 gnd vdd FILL
XFILL_1_NAND2X1_621 gnd vdd FILL
XFILL_0_DFFPOSX1_800 gnd vdd FILL
XFILL_1_NAND2X1_665 gnd vdd FILL
XFILL_0_DFFPOSX1_822 gnd vdd FILL
XFILL_0_OAI21X1_1254 gnd vdd FILL
XFILL_0_OAI21X1_1243 gnd vdd FILL
XFILL_0_NAND2X1_472 gnd vdd FILL
XFILL_0_DFFPOSX1_811 gnd vdd FILL
XFILL_0_NAND2X1_494 gnd vdd FILL
XFILL_0_DFFPOSX1_833 gnd vdd FILL
XFILL_24_6_0 gnd vdd FILL
XFILL_0_NAND2X1_483 gnd vdd FILL
XFILL_0_OAI21X1_1265 gnd vdd FILL
XFILL_1_NAND2X1_643 gnd vdd FILL
XFILL_1_NAND2X1_698 gnd vdd FILL
XFILL_0_DFFPOSX1_877 gnd vdd FILL
XFILL_0_DFFPOSX1_855 gnd vdd FILL
XFILL_0_OAI21X1_1287 gnd vdd FILL
XFILL_0_OAI21X1_1298 gnd vdd FILL
XFILL_0_DFFPOSX1_866 gnd vdd FILL
XFILL_0_OAI21X1_1276 gnd vdd FILL
XFILL_0_DFFPOSX1_844 gnd vdd FILL
XDFFPOSX1_1018 BUFX2_655/A CLKBUF1_8/Y OAI21X1_1595/Y gnd vdd DFFPOSX1
XFILL_0_DFFPOSX1_888 gnd vdd FILL
XDFFPOSX1_1007 BUFX2_672/A CLKBUF1_3/Y OAI21X1_1584/Y gnd vdd DFFPOSX1
XFILL_0_DFFPOSX1_899 gnd vdd FILL
XFILL_5_DFFPOSX1_470 gnd vdd FILL
XFILL_5_DFFPOSX1_481 gnd vdd FILL
XDFFPOSX1_1029 BUFX2_667/A CLKBUF1_52/Y OAI21X1_1606/Y gnd vdd DFFPOSX1
XFILL_5_DFFPOSX1_492 gnd vdd FILL
XFILL_0_BUFX2_209 gnd vdd FILL
XFILL_0_AOI21X1_41 gnd vdd FILL
XFILL_0_AOI21X1_30 gnd vdd FILL
XFILL_0_AOI21X1_52 gnd vdd FILL
XFILL_0_AOI21X1_63 gnd vdd FILL
XFILL_18_13_0 gnd vdd FILL
XFILL_7_7_0 gnd vdd FILL
XFILL_31_15_0 gnd vdd FILL
XFILL_2_DFFPOSX1_905 gnd vdd FILL
XFILL_2_DFFPOSX1_949 gnd vdd FILL
XFILL_2_DFFPOSX1_938 gnd vdd FILL
XFILL_2_DFFPOSX1_916 gnd vdd FILL
XFILL_2_DFFPOSX1_927 gnd vdd FILL
XFILL_2_BUFX4_170 gnd vdd FILL
XFILL_6_DFFPOSX1_1001 gnd vdd FILL
XFILL_6_DFFPOSX1_1012 gnd vdd FILL
XFILL_6_DFFPOSX1_1023 gnd vdd FILL
XFILL_15_6_0 gnd vdd FILL
XFILL_3_XNOR2X1_18 gnd vdd FILL
XFILL_3_XNOR2X1_29 gnd vdd FILL
XFILL_0_BUFX2_710 gnd vdd FILL
XFILL_0_BUFX2_721 gnd vdd FILL
XDFFPOSX1_319 BUFX2_989/A CLKBUF1_17/Y OAI21X1_255/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_732 gnd vdd FILL
XDFFPOSX1_308 BUFX2_977/A CLKBUF1_50/Y OAI21X1_233/Y gnd vdd DFFPOSX1
XFILL_0_NOR2X1_50 gnd vdd FILL
XFILL_0_BUFX2_776 gnd vdd FILL
XFILL_0_BUFX2_754 gnd vdd FILL
XFILL_0_BUFX2_765 gnd vdd FILL
XFILL_0_NOR2X1_94 gnd vdd FILL
XFILL_1_DFFPOSX1_539 gnd vdd FILL
XFILL_1_DFFPOSX1_528 gnd vdd FILL
XFILL_0_NOR2X1_72 gnd vdd FILL
XFILL_0_NOR2X1_83 gnd vdd FILL
XFILL_0_NOR2X1_61 gnd vdd FILL
XFILL_1_DFFPOSX1_506 gnd vdd FILL
XFILL_1_DFFPOSX1_517 gnd vdd FILL
XFILL_0_BUFX2_743 gnd vdd FILL
XFILL_0_BUFX2_787 gnd vdd FILL
XFILL_0_BUFX2_798 gnd vdd FILL
XFILL_6_DFFPOSX1_143 gnd vdd FILL
XFILL_3_DFFPOSX1_5 gnd vdd FILL
XFILL_36_14_0 gnd vdd FILL
XFILL_6_DFFPOSX1_154 gnd vdd FILL
XFILL_6_DFFPOSX1_176 gnd vdd FILL
XFILL_6_DFFPOSX1_165 gnd vdd FILL
XFILL_6_DFFPOSX1_198 gnd vdd FILL
XFILL_6_DFFPOSX1_187 gnd vdd FILL
XBUFX4_340 BUFX4_385/A gnd BUFX4_340/Y vdd BUFX4
XBUFX4_351 BUFX4_385/A gnd BUFX4_351/Y vdd BUFX4
XBUFX4_362 BUFX4_376/A gnd BUFX4_362/Y vdd BUFX4
XBUFX4_373 BUFX4_386/A gnd BUFX4_373/Y vdd BUFX4
XBUFX4_384 BUFX4_384/A gnd BUFX4_384/Y vdd BUFX4
XFILL_0_DFFPOSX1_118 gnd vdd FILL
XFILL_0_DFFPOSX1_107 gnd vdd FILL
XFILL_0_DFFPOSX1_129 gnd vdd FILL
XOAI21X1_906 INVX1_107/Y BUFX4_228/Y OAI21X1_906/C gnd OAI21X1_906/Y vdd OAI21X1
XOAI21X1_928 BUFX4_247/Y BUFX4_329/Y BUFX2_327/A gnd OAI21X1_929/C vdd OAI21X1
XOAI21X1_939 BUFX4_141/Y INVX1_124/Y OAI21X1_939/C gnd OAI21X1_939/Y vdd OAI21X1
XFILL_0_NAND2X1_5 gnd vdd FILL
XOAI21X1_917 BUFX4_154/Y INVX1_113/Y OAI21X1_917/C gnd OAI21X1_917/Y vdd OAI21X1
XOAI21X1_1230 BUFX4_8/A BUFX4_382/Y BUFX2_191/A gnd OAI21X1_1231/C vdd OAI21X1
XOAI21X1_1241 OAI21X1_1241/A BUFX4_146/Y OAI21X1_1241/C gnd OAI21X1_1241/Y vdd OAI21X1
XDFFPOSX1_820 BUFX2_69/A CLKBUF1_11/Y OAI21X1_1124/Y gnd vdd DFFPOSX1
XOAI21X1_1252 INVX1_200/Y INVX2_67/Y INVX4_34/Y gnd OAI21X1_1253/C vdd OAI21X1
XOAI21X1_1263 XNOR2X1_78/Y BUFX4_129/Y OAI21X1_1263/C gnd OAI21X1_1263/Y vdd OAI21X1
XFILL_1_OAI21X1_1450 gnd vdd FILL
XOAI21X1_1274 NOR2X1_187/Y NOR2X1_188/B OAI21X1_1274/C gnd OAI21X1_1274/Y vdd OAI21X1
XDFFPOSX1_842 BUFX2_93/A CLKBUF1_28/Y OAI21X1_1158/Y gnd vdd DFFPOSX1
XDFFPOSX1_831 BUFX2_81/A CLKBUF1_34/Y OAI21X1_1142/Y gnd vdd DFFPOSX1
XDFFPOSX1_875 BUFX2_152/A CLKBUF1_12/Y OAI21X1_1215/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_230 gnd vdd FILL
XFILL_1_OAI21X1_1472 gnd vdd FILL
XOAI21X1_1285 BUFX4_4/A BUFX4_317/Y BUFX2_150/A gnd OAI21X1_1287/C vdd OAI21X1
XDFFPOSX1_853 BUFX2_105/A CLKBUF1_68/Y OAI21X1_1173/Y gnd vdd DFFPOSX1
XOAI21X1_1296 AOI21X1_49/Y NAND2X1_607/Y OAI21X1_1296/C gnd OAI21X1_1296/Y vdd OAI21X1
XFILL_1_OAI21X1_1461 gnd vdd FILL
XFILL_1_OAI21X1_1483 gnd vdd FILL
XDFFPOSX1_864 BUFX2_117/A CLKBUF1_20/Y OAI21X1_1193/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_401 gnd vdd FILL
XFILL_0_OAI21X1_252 gnd vdd FILL
XFILL_0_OAI21X1_263 gnd vdd FILL
XDFFPOSX1_886 BUFX2_135/A CLKBUF1_5/Y OAI21X1_1249/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_241 gnd vdd FILL
XFILL_1_OAI21X1_445 gnd vdd FILL
XDFFPOSX1_897 BUFX2_147/A CLKBUF1_35/Y OAI21X1_1280/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1494 gnd vdd FILL
XFILL_1_OAI21X1_423 gnd vdd FILL
XINVX2_25 bundleStartMajId_i[31] gnd OR2X2_15/B vdd INVX2
XINVX2_36 bundleStartMajId_i[8] gnd INVX2_36/Y vdd INVX2
XFILL_1_OAI21X1_412 gnd vdd FILL
XFILL_1_OAI21X1_434 gnd vdd FILL
XINVX2_14 bundleStartMajId_i[55] gnd NOR2X1_5/A vdd INVX2
XINVX2_58 bundleAddress_i[58] gnd INVX2_58/Y vdd INVX2
XFILL_0_OAI21X1_296 gnd vdd FILL
XFILL_0_OAI21X1_274 gnd vdd FILL
XFILL_1_OAI21X1_478 gnd vdd FILL
XFILL_2_OAI21X1_627 gnd vdd FILL
XFILL_1_OAI21X1_456 gnd vdd FILL
XINVX2_47 NOR3X1_4/A gnd INVX2_47/Y vdd INVX2
XINVX2_69 bundleAddress_i[45] gnd INVX2_69/Y vdd INVX2
XFILL_1_OAI21X1_467 gnd vdd FILL
XFILL_0_OAI21X1_285 gnd vdd FILL
XFILL_1_OAI21X1_489 gnd vdd FILL
XFILL_1_INVX4_25 gnd vdd FILL
XFILL_1_INVX4_36 gnd vdd FILL
XFILL_0_OAI21X1_1040 gnd vdd FILL
XFILL_1_BUFX4_204 gnd vdd FILL
XFILL_0_OAI21X1_1051 gnd vdd FILL
XFILL_0_DFFPOSX1_630 gnd vdd FILL
XFILL_0_OAI21X1_1084 gnd vdd FILL
XFILL_0_OAI21X1_1062 gnd vdd FILL
XFILL_1_NAND2X1_462 gnd vdd FILL
XFILL_0_NAND2X1_291 gnd vdd FILL
XFILL_0_DFFPOSX1_652 gnd vdd FILL
XFILL_0_OAI21X1_1073 gnd vdd FILL
XFILL_1_BUFX4_215 gnd vdd FILL
XFILL_1_BUFX4_237 gnd vdd FILL
XFILL_0_DFFPOSX1_641 gnd vdd FILL
XFILL_0_NAND2X1_280 gnd vdd FILL
XFILL_1_BUFX4_226 gnd vdd FILL
XFILL_1_BUFX4_248 gnd vdd FILL
XFILL_1_NAND2X1_495 gnd vdd FILL
XFILL_0_OAI21X1_1095 gnd vdd FILL
XFILL_1_BUFX4_259 gnd vdd FILL
XFILL_0_DFFPOSX1_663 gnd vdd FILL
XFILL_0_DFFPOSX1_674 gnd vdd FILL
XFILL_0_DFFPOSX1_685 gnd vdd FILL
XFILL_0_DFFPOSX1_696 gnd vdd FILL
XFILL_20_12_1 gnd vdd FILL
XFILL_2_BUFX4_20 gnd vdd FILL
XFILL_0_DFFPOSX1_19 gnd vdd FILL
XFILL_2_BUFX4_53 gnd vdd FILL
XFILL_2_XNOR2X1_8 gnd vdd FILL
XFILL_1_OAI21X1_990 gnd vdd FILL
XFILL_2_OAI21X1_1101 gnd vdd FILL
XFILL_2_DFFPOSX1_713 gnd vdd FILL
XBUFX2_811 BUFX2_811/A gnd tid1_o[59] vdd BUFX2
XFILL_2_DFFPOSX1_702 gnd vdd FILL
XBUFX2_800 BUFX2_800/A gnd tid1_o[60] vdd BUFX2
XBUFX2_822 BUFX2_822/A gnd tid1_o[58] vdd BUFX2
XBUFX2_844 BUFX2_844/A gnd tid2_o[52] vdd BUFX2
XFILL_2_DFFPOSX1_746 gnd vdd FILL
XFILL_2_DFFPOSX1_757 gnd vdd FILL
XBUFX2_855 BUFX2_855/A gnd tid2_o[42] vdd BUFX2
XFILL_2_DFFPOSX1_735 gnd vdd FILL
XBUFX2_833 BUFX2_833/A gnd tid1_o[57] vdd BUFX2
XFILL_2_DFFPOSX1_724 gnd vdd FILL
XBUFX2_877 BUFX2_877/A gnd tid2_o[22] vdd BUFX2
XBUFX2_888 BUFX2_888/A gnd tid2_o[12] vdd BUFX2
XBUFX2_866 BUFX2_866/A gnd tid2_o[32] vdd BUFX2
XFILL_2_DFFPOSX1_779 gnd vdd FILL
XFILL_2_DFFPOSX1_768 gnd vdd FILL
XFILL_0_NOR2X1_217 gnd vdd FILL
XBUFX2_899 BUFX2_899/A gnd tid2_o[2] vdd BUFX2
XFILL_0_NOR2X1_206 gnd vdd FILL
XFILL_0_NOR2X1_228 gnd vdd FILL
XFILL_31_9_1 gnd vdd FILL
XFILL_30_4_0 gnd vdd FILL
XFILL_25_11_1 gnd vdd FILL
XFILL_3_CLKBUF1_8 gnd vdd FILL
XDFFPOSX1_127 BUFX2_797/A CLKBUF1_32/Y OAI21X1_1801/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_303 gnd vdd FILL
XFILL_0_BUFX2_540 gnd vdd FILL
XDFFPOSX1_116 BUFX2_785/A CLKBUF1_47/Y OAI21X1_1790/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_314 gnd vdd FILL
XFILL_0_BUFX2_551 gnd vdd FILL
XDFFPOSX1_105 BUFX2_822/A CLKBUF1_71/Y OAI21X1_1779/Y gnd vdd DFFPOSX1
XDFFPOSX1_138 BUFX2_809/A CLKBUF1_86/Y OAI21X1_1812/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_336 gnd vdd FILL
XFILL_1_DFFPOSX1_325 gnd vdd FILL
XFILL_0_BUFX2_584 gnd vdd FILL
XDFFPOSX1_149 BUFX2_821/A CLKBUF1_21/Y OAI21X1_1823/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_347 gnd vdd FILL
XFILL_0_BUFX2_573 gnd vdd FILL
XFILL_0_BUFX2_562 gnd vdd FILL
XFILL_0_BUFX2_595 gnd vdd FILL
XFILL_1_DFFPOSX1_358 gnd vdd FILL
XNAND2X1_208 BUFX2_486/A BUFX4_236/Y gnd OAI21X1_453/C vdd NAND2X1
XFILL_1_DFFPOSX1_369 gnd vdd FILL
XNAND2X1_219 OAI21X1_460/Y OAI21X1_462/A gnd OAI21X1_461/A vdd NAND2X1
XFILL_4_DFFPOSX1_818 gnd vdd FILL
XFILL_4_DFFPOSX1_807 gnd vdd FILL
XFILL_4_DFFPOSX1_829 gnd vdd FILL
XFILL_38_5_0 gnd vdd FILL
XBUFX4_170 BUFX4_14/Y gnd BUFX4_170/Y vdd BUFX4
XFILL_4_CLKBUF1_41 gnd vdd FILL
XFILL_0_INVX1_70 gnd vdd FILL
XBUFX4_181 BUFX4_20/Y gnd BUFX4_181/Y vdd BUFX4
XFILL_4_CLKBUF1_52 gnd vdd FILL
XFILL_4_CLKBUF1_74 gnd vdd FILL
XFILL_4_CLKBUF1_63 gnd vdd FILL
XFILL_4_CLKBUF1_85 gnd vdd FILL
XFILL_0_BUFX2_12 gnd vdd FILL
XFILL_0_INVX1_92 gnd vdd FILL
XFILL_0_12_1 gnd vdd FILL
XBUFX4_192 BUFX4_26/Y gnd BUFX4_192/Y vdd BUFX4
XNOR2X1_230 bundleAddress_i[8] INVX1_226/Y gnd NOR2X1_230/Y vdd NOR2X1
XFILL_0_INVX1_81 gnd vdd FILL
XFILL_0_BUFX2_23 gnd vdd FILL
XFILL_4_CLKBUF1_96 gnd vdd FILL
XFILL_0_BUFX2_45 gnd vdd FILL
XFILL_0_BUFX2_34 gnd vdd FILL
XFILL_0_BUFX2_67 gnd vdd FILL
XFILL_22_9_1 gnd vdd FILL
XFILL_0_BUFX2_56 gnd vdd FILL
XFILL_1_BUFX2_708 gnd vdd FILL
XFILL_0_BUFX2_78 gnd vdd FILL
XFILL_1_NOR2X1_26 gnd vdd FILL
XFILL_1_NOR2X1_15 gnd vdd FILL
XFILL_0_BUFX2_89 gnd vdd FILL
XOAI21X1_714 BUFX4_171/Y BUFX4_48/Y BUFX2_596/A gnd OAI21X1_715/C vdd OAI21X1
XOAI21X1_703 OAI21X1_703/A BUFX4_290/Y OAI21X1_703/C gnd OAI21X1_703/Y vdd OAI21X1
XFILL_21_4_0 gnd vdd FILL
XFILL_1_NOR2X1_48 gnd vdd FILL
XFILL_1_NOR2X1_59 gnd vdd FILL
XOAI21X1_758 BUFX4_171/Y BUFX4_48/Y BUFX2_614/A gnd OAI21X1_759/C vdd OAI21X1
XOAI21X1_747 INVX1_39/Y BUFX4_286/Y OAI21X1_747/C gnd OAI21X1_747/Y vdd OAI21X1
XOAI21X1_736 OAI21X1_736/A AOI21X1_32/Y OAI21X1_736/C gnd OAI21X1_736/Y vdd OAI21X1
XFILL_3_DFFPOSX1_408 gnd vdd FILL
XFILL_3_DFFPOSX1_419 gnd vdd FILL
XOAI21X1_725 BUFX4_177/Y BUFX4_33/Y BUFX2_601/A gnd OAI21X1_726/C vdd OAI21X1
XOAI21X1_769 XNOR2X1_51/Y BUFX4_300/Y OAI21X1_769/C gnd OAI21X1_769/Y vdd OAI21X1
XDFFPOSX1_650 BUFX2_305/A CLKBUF1_78/Y OAI21X1_878/Y gnd vdd DFFPOSX1
XOAI21X1_1082 BUFX4_360/Y INVX1_178/Y NAND2X1_448/Y gnd OAI21X1_1082/Y vdd OAI21X1
XOAI21X1_1071 BUFX4_384/Y INVX2_76/Y NAND2X1_437/Y gnd OAI21X1_1071/Y vdd OAI21X1
XOAI21X1_1060 BUFX4_354/Y INVX1_175/Y NAND2X1_426/Y gnd OAI21X1_1060/Y vdd OAI21X1
XDFFPOSX1_672 BUFX2_310/A CLKBUF1_101/Y OAI21X1_900/Y gnd vdd DFFPOSX1
XDFFPOSX1_683 BUFX2_348/A CLKBUF1_39/Y OAI21X1_915/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1291 gnd vdd FILL
XDFFPOSX1_661 BUFX2_298/A CLKBUF1_32/Y OAI21X1_889/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_870 gnd vdd FILL
XFILL_1_OAI21X1_1280 gnd vdd FILL
XOAI21X1_1093 BUFX4_343/Y INVX1_180/Y NAND2X1_459/Y gnd OAI21X1_1093/Y vdd OAI21X1
XDFFPOSX1_694 BUFX2_331/A CLKBUF1_96/Y OAI21X1_937/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_881 gnd vdd FILL
XFILL_1_OAI21X1_253 gnd vdd FILL
XFILL_1_OAI21X1_231 gnd vdd FILL
XFILL_1_OAI21X1_242 gnd vdd FILL
XFILL_0_NOR2X1_3 gnd vdd FILL
XFILL_1_DFFPOSX1_892 gnd vdd FILL
XFILL_1_OAI21X1_220 gnd vdd FILL
XNAND2X1_720 BUFX2_822/A BUFX4_374/Y gnd NAND2X1_720/Y vdd NAND2X1
XNAND2X1_742 BUFX2_797/A BUFX4_332/Y gnd NAND2X1_742/Y vdd NAND2X1
XNAND2X1_753 BUFX2_809/A BUFX4_313/Y gnd NAND2X1_753/Y vdd NAND2X1
XFILL_1_OAI21X1_275 gnd vdd FILL
XNAND2X1_764 BUFX2_821/A BUFX4_313/Y gnd NAND2X1_764/Y vdd NAND2X1
XFILL_1_OAI21X1_286 gnd vdd FILL
XNAND2X1_731 BUFX2_785/A BUFX4_334/Y gnd NAND2X1_731/Y vdd NAND2X1
XFILL_1_OAI21X1_264 gnd vdd FILL
XFILL_2_OAI21X1_435 gnd vdd FILL
XFILL_1_OAI21X1_297 gnd vdd FILL
XFILL_5_11_1 gnd vdd FILL
XFILL_29_5_0 gnd vdd FILL
XBUFX2_107 BUFX2_107/A gnd addr2_o[16] vdd BUFX2
XFILL_2_XNOR2X1_15 gnd vdd FILL
XFILL_2_XNOR2X1_37 gnd vdd FILL
XFILL_2_XNOR2X1_26 gnd vdd FILL
XFILL_4_5_0 gnd vdd FILL
XBUFX2_129 BUFX2_129/A gnd addr3_o[63] vdd BUFX2
XFILL_2_XNOR2X1_59 gnd vdd FILL
XFILL_2_XNOR2X1_48 gnd vdd FILL
XBUFX2_118 BUFX2_118/A gnd addr2_o[6] vdd BUFX2
XFILL_0_DFFPOSX1_460 gnd vdd FILL
XFILL_1_NAND2X1_292 gnd vdd FILL
XFILL_13_9_1 gnd vdd FILL
XFILL_1_NAND2X1_281 gnd vdd FILL
XFILL_2_DFFPOSX1_2 gnd vdd FILL
XFILL_1_NAND2X1_270 gnd vdd FILL
XFILL_0_DFFPOSX1_493 gnd vdd FILL
XFILL_0_DFFPOSX1_471 gnd vdd FILL
XFILL_0_DFFPOSX1_482 gnd vdd FILL
XINVX8_1 INVX8_1/A gnd INVX8_1/Y vdd INVX8
XFILL_12_4_0 gnd vdd FILL
XFILL_3_DFFPOSX1_920 gnd vdd FILL
XFILL_3_DFFPOSX1_931 gnd vdd FILL
XFILL_3_DFFPOSX1_942 gnd vdd FILL
XFILL_3_DFFPOSX1_953 gnd vdd FILL
XFILL_3_DFFPOSX1_964 gnd vdd FILL
XFILL_3_DFFPOSX1_975 gnd vdd FILL
XFILL_3_DFFPOSX1_997 gnd vdd FILL
XFILL_3_DFFPOSX1_986 gnd vdd FILL
XBUFX4_10 BUFX4_10/A gnd BUFX4_10/Y vdd BUFX4
XFILL_2_OAI21X1_980 gnd vdd FILL
XBUFX4_43 BUFX4_64/A gnd BUFX4_43/Y vdd BUFX4
XBUFX4_32 BUFX4_59/A gnd BUFX4_32/Y vdd BUFX4
XBUFX4_21 BUFX4_26/A gnd BUFX4_21/Y vdd BUFX4
XBUFX4_65 BUFX4_82/A gnd BUFX4_65/Y vdd BUFX4
XBUFX4_87 clock_i gnd BUFX4_87/Y vdd BUFX4
XBUFX4_54 BUFX4_71/A gnd BUFX4_54/Y vdd BUFX4
XBUFX4_76 BUFX4_82/A gnd BUFX4_76/Y vdd BUFX4
XFILL_2_DFFPOSX1_510 gnd vdd FILL
XBUFX4_98 BUFX4_2/A gnd BUFX4_98/Y vdd BUFX4
XFILL_2_DFFPOSX1_521 gnd vdd FILL
XFILL_2_DFFPOSX1_532 gnd vdd FILL
XFILL_11_17_1 gnd vdd FILL
XBUFX2_630 BUFX2_630/A gnd majID4_o[58] vdd BUFX2
XFILL_2_DFFPOSX1_543 gnd vdd FILL
XBUFX2_663 BUFX2_663/A gnd pid1_o[10] vdd BUFX2
XBUFX2_652 BUFX2_652/A gnd pid1_o[20] vdd BUFX2
XFILL_0_OAI21X1_1809 gnd vdd FILL
XFILL_2_DFFPOSX1_565 gnd vdd FILL
XBUFX2_641 BUFX2_641/A gnd majID4_o[57] vdd BUFX2
XFILL_2_DFFPOSX1_554 gnd vdd FILL
XBUFX2_696 BUFX2_696/A gnd pid2_o[9] vdd BUFX2
XFILL_2_DFFPOSX1_598 gnd vdd FILL
XFILL_2_DFFPOSX1_587 gnd vdd FILL
XBUFX2_685 BUFX2_685/A gnd pid2_o[19] vdd BUFX2
XFILL_2_DFFPOSX1_576 gnd vdd FILL
XBUFX2_674 BUFX2_674/A gnd pid1_o[0] vdd BUFX2
XOR2X2_13 OR2X2_13/A OR2X2_13/B gnd OR2X2_13/Y vdd OR2X2
XFILL_1_DFFPOSX1_111 gnd vdd FILL
XFILL_1_DFFPOSX1_100 gnd vdd FILL
XFILL_1_DFFPOSX1_122 gnd vdd FILL
XOR2X2_6 OR2X2_6/A OR2X2_6/B gnd OR2X2_6/Y vdd OR2X2
XFILL_2_AOI21X1_15 gnd vdd FILL
XINVX2_170 bundleTid_i[39] gnd INVX2_170/Y vdd INVX2
XFILL_1_DFFPOSX1_133 gnd vdd FILL
XFILL_0_BUFX2_381 gnd vdd FILL
XFILL_1_DFFPOSX1_144 gnd vdd FILL
XINVX2_181 bundleTid_i[28] gnd INVX2_181/Y vdd INVX2
XFILL_1_DFFPOSX1_155 gnd vdd FILL
XINVX2_192 bundleTid_i[17] gnd INVX2_192/Y vdd INVX2
XFILL_0_BUFX2_370 gnd vdd FILL
XFILL_0_BUFX2_392 gnd vdd FILL
XFILL_1_DFFPOSX1_188 gnd vdd FILL
XFILL_1_DFFPOSX1_166 gnd vdd FILL
XFILL_1_DFFPOSX1_177 gnd vdd FILL
XXNOR2X1_8 AND2X2_3/Y bundleStartMajId_i[41] gnd XNOR2X1_8/Y vdd XNOR2X1
XFILL_4_DFFPOSX1_604 gnd vdd FILL
XFILL_1_DFFPOSX1_199 gnd vdd FILL
XFILL_4_DFFPOSX1_615 gnd vdd FILL
XFILL_16_16_1 gnd vdd FILL
XFILL_4_DFFPOSX1_626 gnd vdd FILL
XFILL_4_DFFPOSX1_637 gnd vdd FILL
XFILL_4_DFFPOSX1_648 gnd vdd FILL
XFILL_4_DFFPOSX1_659 gnd vdd FILL
XFILL_10_12_0 gnd vdd FILL
XFILL_1_BUFX2_505 gnd vdd FILL
XFILL_2_AND2X2_7 gnd vdd FILL
XOAI21X1_500 BUFX4_93/Y BUFX4_362/Y BUFX2_521/A gnd OAI21X1_501/C vdd OAI21X1
XFILL_1_BUFX2_538 gnd vdd FILL
XFILL_1_BUFX2_549 gnd vdd FILL
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XOAI21X1_511 BUFX4_7/A BUFX4_355/Y BUFX2_555/A gnd OAI21X1_512/C vdd OAI21X1
XOAI21X1_522 INVX4_29/Y NOR2X1_4/B NOR2X1_5/A gnd OAI21X1_522/Y vdd OAI21X1
XOAI21X1_566 BUFX4_10/A BUFX4_378/Y BUFX2_539/A gnd OAI21X1_567/C vdd OAI21X1
XOAI21X1_555 BUFX4_10/A BUFX4_319/Y BUFX2_532/A gnd OAI21X1_556/C vdd OAI21X1
XOAI21X1_533 BUFX4_112/Y BUFX4_372/Y BUFX2_524/A gnd OAI21X1_534/C vdd OAI21X1
XFILL_3_DFFPOSX1_205 gnd vdd FILL
XOAI21X1_544 BUFX4_9/Y BUFX4_345/Y BUFX2_529/A gnd OAI21X1_546/C vdd OAI21X1
XFILL_3_DFFPOSX1_216 gnd vdd FILL
XFILL_3_DFFPOSX1_227 gnd vdd FILL
XFILL_3_DFFPOSX1_249 gnd vdd FILL
XFILL_3_DFFPOSX1_238 gnd vdd FILL
XOAI21X1_577 BUFX4_108/Y BUFX4_378/Y BUFX2_543/A gnd OAI21X1_578/C vdd OAI21X1
XOAI21X1_599 BUFX4_10/A BUFX4_346/Y BUFX2_552/A gnd OAI21X1_600/C vdd OAI21X1
XOAI21X1_588 OR2X2_8/A OR2X2_9/A OAI21X1_588/C gnd OAI21X1_590/A vdd OAI21X1
XFILL_6_DFFPOSX1_709 gnd vdd FILL
XDFFPOSX1_480 BUFX2_514/A CLKBUF1_9/Y OAI21X1_494/Y gnd vdd DFFPOSX1
XDFFPOSX1_491 BUFX2_582/A CLKBUF1_94/Y OAI21X1_521/Y gnd vdd DFFPOSX1
XFILL_34_17_1 gnd vdd FILL
XNAND2X1_561 bundleAddress_i[16] bundleAddress_i[15] gnd INVX1_195/A vdd NAND2X1
XNAND2X1_550 BUFX2_102/A INVX8_1/A gnd NAND2X1_550/Y vdd NAND2X1
XNAND2X1_572 BUFX4_239/Y NAND2X1_572/B gnd NAND2X1_572/Y vdd NAND2X1
XFILL_2_OAI21X1_298 gnd vdd FILL
XNAND2X1_594 bundleAddress_i[50] INVX2_96/Y gnd NOR2X1_183/A vdd NAND2X1
XNAND2X1_583 BUFX2_120/A BUFX4_188/Y gnd NAND2X1_583/Y vdd NAND2X1
XFILL_15_11_0 gnd vdd FILL
XFILL_1_DFFPOSX1_1018 gnd vdd FILL
XFILL_1_DFFPOSX1_1007 gnd vdd FILL
XFILL_1_DFFPOSX1_1029 gnd vdd FILL
XFILL_0_DFFPOSX1_290 gnd vdd FILL
XOAI21X1_1807 BUFX4_329/Y INVX2_179/Y NAND2X1_748/Y gnd OAI21X1_1807/Y vdd OAI21X1
XOAI21X1_1818 BUFX4_336/Y INVX2_190/Y NAND2X1_759/Y gnd OAI21X1_1818/Y vdd OAI21X1
XFILL_3_DFFPOSX1_750 gnd vdd FILL
XOAI21X1_1829 BUFX4_367/Y INVX2_201/Y NAND2X1_770/Y gnd OAI21X1_1829/Y vdd OAI21X1
XFILL_3_DFFPOSX1_761 gnd vdd FILL
XFILL_3_DFFPOSX1_772 gnd vdd FILL
XFILL_3_CLKBUF1_60 gnd vdd FILL
XFILL_3_DFFPOSX1_783 gnd vdd FILL
XFILL_3_CLKBUF1_93 gnd vdd FILL
XFILL_0_OAI21X1_829 gnd vdd FILL
XFILL_0_OAI21X1_807 gnd vdd FILL
XFILL_0_OAI21X1_818 gnd vdd FILL
XFILL_3_CLKBUF1_82 gnd vdd FILL
XFILL_3_CLKBUF1_71 gnd vdd FILL
XFILL_3_DFFPOSX1_794 gnd vdd FILL
XFILL_33_12_0 gnd vdd FILL
XFILL_36_8_1 gnd vdd FILL
XFILL_35_3_0 gnd vdd FILL
XFILL_2_DFFPOSX1_340 gnd vdd FILL
XFILL_0_OAI21X1_1606 gnd vdd FILL
XFILL_0_OAI21X1_1628 gnd vdd FILL
XFILL_0_OAI21X1_1639 gnd vdd FILL
XBUFX2_460 BUFX2_460/A gnd majID2_o[52] vdd BUFX2
XBUFX2_471 BUFX2_471/A gnd majID2_o[42] vdd BUFX2
XFILL_2_DFFPOSX1_373 gnd vdd FILL
XFILL_0_OAI21X1_1617 gnd vdd FILL
XFILL_2_DFFPOSX1_362 gnd vdd FILL
XFILL_2_DFFPOSX1_351 gnd vdd FILL
XFILL_2_DFFPOSX1_395 gnd vdd FILL
XBUFX2_493 BUFX2_493/A gnd majID2_o[22] vdd BUFX2
XBUFX2_482 INVX1_14/A gnd majID2_o[32] vdd BUFX2
XFILL_2_DFFPOSX1_384 gnd vdd FILL
XFILL_5_DFFPOSX1_822 gnd vdd FILL
XFILL_5_DFFPOSX1_811 gnd vdd FILL
XFILL_5_DFFPOSX1_800 gnd vdd FILL
XFILL_5_DFFPOSX1_855 gnd vdd FILL
XFILL_5_DFFPOSX1_833 gnd vdd FILL
XFILL_5_DFFPOSX1_844 gnd vdd FILL
XFILL_5_DFFPOSX1_888 gnd vdd FILL
XFILL_5_DFFPOSX1_877 gnd vdd FILL
XFILL_5_DFFPOSX1_866 gnd vdd FILL
XFILL_1_XNOR2X1_12 gnd vdd FILL
XFILL_1_XNOR2X1_23 gnd vdd FILL
XFILL_5_DFFPOSX1_899 gnd vdd FILL
XFILL_1_XNOR2X1_45 gnd vdd FILL
XFILL_1_XNOR2X1_34 gnd vdd FILL
XFILL_1_XNOR2X1_56 gnd vdd FILL
XFILL_1_XNOR2X1_89 gnd vdd FILL
XFILL_1_XNOR2X1_78 gnd vdd FILL
XFILL_1_XNOR2X1_67 gnd vdd FILL
XFILL_38_11_0 gnd vdd FILL
XFILL_4_DFFPOSX1_412 gnd vdd FILL
XFILL_4_DFFPOSX1_401 gnd vdd FILL
XFILL_4_DFFPOSX1_445 gnd vdd FILL
XFILL_4_DFFPOSX1_423 gnd vdd FILL
XFILL_4_DFFPOSX1_434 gnd vdd FILL
XFILL_4_DFFPOSX1_478 gnd vdd FILL
XFILL_4_DFFPOSX1_456 gnd vdd FILL
XFILL_4_DFFPOSX1_467 gnd vdd FILL
XFILL_27_8_1 gnd vdd FILL
XFILL_4_DFFPOSX1_489 gnd vdd FILL
XFILL_2_8_1 gnd vdd FILL
XFILL_26_3_0 gnd vdd FILL
XFILL_1_3_0 gnd vdd FILL
XFILL_1_BUFX2_302 gnd vdd FILL
XFILL_1_BUFX2_335 gnd vdd FILL
XFILL_1_BUFX2_379 gnd vdd FILL
XOAI21X1_330 BUFX4_365/Y INVX2_9/Y NAND2X1_74/Y gnd OAI21X1_330/Y vdd OAI21X1
XFILL_10_7_1 gnd vdd FILL
XOAI21X1_341 BUFX4_345/Y INVX1_1/Y NAND2X1_85/Y gnd OAI21X1_341/Y vdd OAI21X1
XFILL_1_BUFX2_357 gnd vdd FILL
XFILL_1_BUFX2_346 gnd vdd FILL
XOAI21X1_374 BUFX4_358/Y INVX2_31/Y OAI21X1_374/C gnd OAI21X1_374/Y vdd OAI21X1
XOAI21X1_352 OAI21X1_2/A INVX4_10/Y NAND2X1_96/Y gnd OAI21X1_352/Y vdd OAI21X1
XOAI21X1_363 BUFX4_337/Y OR2X2_8/B OAI21X1_363/C gnd OAI21X1_363/Y vdd OAI21X1
XOAI21X1_385 BUFX4_356/Y INVX4_25/Y OAI21X1_385/C gnd OAI21X1_385/Y vdd OAI21X1
XOAI21X1_396 OAI21X1_396/A BUFX4_180/Y OAI21X1_396/C gnd OAI21X1_396/Y vdd OAI21X1
XAND2X2_8 NOR3X1_2/Y INVX1_33/A gnd AND2X2_8/Y vdd AND2X2
XFILL_9_4_0 gnd vdd FILL
XNAND2X1_380 BUFX2_295/A BUFX4_186/Y gnd OAI21X1_886/C vdd NAND2X1
XNAND2X1_391 BUFX2_307/A BUFX4_189/Y gnd OAI21X1_897/C vdd NAND2X1
XFILL_0_INVX1_101 gnd vdd FILL
XFILL_0_INVX1_112 gnd vdd FILL
XFILL_18_8_1 gnd vdd FILL
XFILL_0_NAND2X1_109 gnd vdd FILL
XFILL_4_DFFPOSX1_990 gnd vdd FILL
XFILL_0_INVX1_123 gnd vdd FILL
XFILL_0_INVX1_145 gnd vdd FILL
XFILL_1_AOI21X1_23 gnd vdd FILL
XFILL_17_3_0 gnd vdd FILL
XFILL_1_AOI21X1_12 gnd vdd FILL
XFILL_0_INVX1_134 gnd vdd FILL
XFILL_0_INVX1_189 gnd vdd FILL
XFILL_0_INVX1_178 gnd vdd FILL
XFILL_0_INVX1_156 gnd vdd FILL
XFILL_1_AOI21X1_45 gnd vdd FILL
XFILL_1_AOI21X1_34 gnd vdd FILL
XFILL_1_AOI21X1_56 gnd vdd FILL
XFILL_0_INVX1_167 gnd vdd FILL
XFILL_5_DFFPOSX1_107 gnd vdd FILL
XFILL_5_DFFPOSX1_118 gnd vdd FILL
XFILL_5_DFFPOSX1_129 gnd vdd FILL
XOAI21X1_1604 BUFX4_332/Y INVX2_140/Y NAND2X1_673/Y gnd OAI21X1_1604/Y vdd OAI21X1
XOAI21X1_1615 INVX2_118/Y BUFX4_235/Y NAND2X1_683/Y gnd DFFPOSX1_5/D vdd OAI21X1
XOAI21X1_1637 INVX2_140/Y BUFX4_205/Y NAND2X1_705/Y gnd DFFPOSX1_27/D vdd OAI21X1
XOAI21X1_1648 BUFX4_3/Y BUFX4_316/Y BUFX2_714/A gnd OAI21X1_1649/C vdd OAI21X1
XFILL_1_OAI21X1_1824 gnd vdd FILL
XFILL_1_OAI21X1_1813 gnd vdd FILL
XOAI21X1_1626 INVX2_129/Y BUFX4_183/Y NAND2X1_694/Y gnd DFFPOSX1_16/D vdd OAI21X1
XFILL_1_OAI21X1_1802 gnd vdd FILL
XFILL_3_DFFPOSX1_591 gnd vdd FILL
XFILL_3_DFFPOSX1_580 gnd vdd FILL
XFILL_0_OAI21X1_604 gnd vdd FILL
XOAI21X1_1659 BUFX4_173/Y INVX2_123/Y OAI21X1_1659/C gnd DFFPOSX1_42/D vdd OAI21X1
XFILL_0_OAI21X1_626 gnd vdd FILL
XFILL_1_OAI21X1_808 gnd vdd FILL
XFILL_1_OAI21X1_819 gnd vdd FILL
XFILL_0_OAI21X1_637 gnd vdd FILL
XFILL_0_OAI21X1_615 gnd vdd FILL
XFILL_0_OAI21X1_648 gnd vdd FILL
XFILL_0_OAI21X1_659 gnd vdd FILL
XFILL_1_AND2X2_16 gnd vdd FILL
XFILL_1_AND2X2_27 gnd vdd FILL
XFILL_0_NAND2X1_610 gnd vdd FILL
XFILL_0_OAI21X1_1414 gnd vdd FILL
XFILL_0_OAI21X1_1403 gnd vdd FILL
XFILL_0_NAND2X1_632 gnd vdd FILL
XFILL_0_NAND2X1_654 gnd vdd FILL
XFILL_0_NAND2X1_621 gnd vdd FILL
XFILL_0_NAND2X1_643 gnd vdd FILL
XFILL_2_DFFPOSX1_181 gnd vdd FILL
XFILL_0_NAND2X1_665 gnd vdd FILL
XFILL_0_NAND2X1_676 gnd vdd FILL
XFILL_0_OAI21X1_1425 gnd vdd FILL
XFILL_0_OAI21X1_1436 gnd vdd FILL
XFILL_2_DFFPOSX1_170 gnd vdd FILL
XFILL_0_OAI21X1_1458 gnd vdd FILL
XFILL_0_OAI21X1_1447 gnd vdd FILL
XBUFX2_290 INVX1_52/A gnd instr1_o[24] vdd BUFX2
XFILL_0_NAND2X1_687 gnd vdd FILL
XFILL_0_NAND2X1_698 gnd vdd FILL
XFILL_0_OAI21X1_1469 gnd vdd FILL
XFILL_2_DFFPOSX1_192 gnd vdd FILL
XFILL_5_DFFPOSX1_630 gnd vdd FILL
XFILL_4_DFFPOSX1_9 gnd vdd FILL
XFILL_5_DFFPOSX1_652 gnd vdd FILL
XFILL_5_DFFPOSX1_663 gnd vdd FILL
XFILL_5_DFFPOSX1_641 gnd vdd FILL
XFILL_24_17_0 gnd vdd FILL
XFILL_5_DFFPOSX1_696 gnd vdd FILL
XFILL_5_DFFPOSX1_674 gnd vdd FILL
XFILL_5_DFFPOSX1_685 gnd vdd FILL
XFILL_4_DFFPOSX1_220 gnd vdd FILL
XFILL_4_DFFPOSX1_242 gnd vdd FILL
XFILL_2_OAI21X1_1519 gnd vdd FILL
XFILL_4_DFFPOSX1_253 gnd vdd FILL
XFILL_4_DFFPOSX1_231 gnd vdd FILL
XFILL_4_DFFPOSX1_275 gnd vdd FILL
XFILL_4_DFFPOSX1_264 gnd vdd FILL
XFILL_4_DFFPOSX1_297 gnd vdd FILL
XFILL_4_DFFPOSX1_286 gnd vdd FILL
XFILL_2_BUFX4_330 gnd vdd FILL
XFILL_2_BUFX4_363 gnd vdd FILL
XFILL_2_CLKBUF1_90 gnd vdd FILL
XFILL_29_16_0 gnd vdd FILL
XFILL_1_BUFX2_110 gnd vdd FILL
XFILL_1_BUFX2_132 gnd vdd FILL
XFILL_1_BUFX2_143 gnd vdd FILL
XFILL_1_BUFX2_154 gnd vdd FILL
XFILL_1_BUFX2_187 gnd vdd FILL
XFILL_1_BUFX2_198 gnd vdd FILL
XFILL_0_BUFX2_914 gnd vdd FILL
XFILL_0_BUFX2_925 gnd vdd FILL
XOAI21X1_160 BUFX4_4/A BUFX4_336/Y BUFX2_944/A gnd OAI21X1_161/C vdd OAI21X1
XFILL_1_OAI21X1_1109 gnd vdd FILL
XOAI21X1_171 BUFX4_141/Y INVX2_195/Y OAI21X1_171/C gnd OAI21X1_171/Y vdd OAI21X1
XOAI21X1_182 BUFX4_7/A BUFX4_367/Y BUFX2_956/A gnd OAI21X1_183/C vdd OAI21X1
XFILL_0_BUFX2_903 gnd vdd FILL
XFILL_0_BUFX2_958 gnd vdd FILL
XFILL_0_BUFX2_947 gnd vdd FILL
XFILL_0_BUFX2_936 gnd vdd FILL
XINVX1_224 INVX1_224/A gnd INVX1_224/Y vdd INVX1
XINVX1_213 INVX1_213/A gnd INVX1_213/Y vdd INVX1
XINVX1_202 INVX1_202/A gnd INVX1_202/Y vdd INVX1
XOAI21X1_193 BUFX4_124/Y INVX2_4/Y OAI21X1_193/C gnd OAI21X1_193/Y vdd OAI21X1
XFILL_0_BUFX2_969 gnd vdd FILL
XFILL_6_DFFPOSX1_325 gnd vdd FILL
XFILL_6_DFFPOSX1_336 gnd vdd FILL
XFILL_6_DFFPOSX1_358 gnd vdd FILL
XFILL_6_DFFPOSX1_347 gnd vdd FILL
XFILL_6_DFFPOSX1_369 gnd vdd FILL
XNAND2X1_24 BUFX2_849/A BUFX4_223/Y gnd OAI21X1_24/C vdd NAND2X1
XNAND2X1_13 BUFX2_886/A BUFX4_196/Y gnd OAI21X1_13/C vdd NAND2X1
XNAND2X1_35 BUFX2_861/A BUFX4_234/Y gnd OAI21X1_35/C vdd NAND2X1
XNAND2X1_46 BUFX2_873/A BUFX4_193/Y gnd OAI21X1_46/C vdd NAND2X1
XNAND2X1_57 BUFX2_885/A BUFX4_195/Y gnd OAI21X1_57/C vdd NAND2X1
XNAND2X1_68 BUFX2_898/A BUFX4_186/Y gnd OAI21X1_68/C vdd NAND2X1
XFILL_0_XNOR2X1_20 gnd vdd FILL
XFILL_0_XNOR2X1_53 gnd vdd FILL
XFILL_0_XNOR2X1_42 gnd vdd FILL
XFILL_4_17_0 gnd vdd FILL
XNAND2X1_79 BUFX2_454/A BUFX4_355/Y gnd NAND2X1_79/Y vdd NAND2X1
XFILL_0_XNOR2X1_31 gnd vdd FILL
XFILL_0_XNOR2X1_64 gnd vdd FILL
XFILL_0_XNOR2X1_75 gnd vdd FILL
XFILL_0_XNOR2X1_97 gnd vdd FILL
XFILL_0_XNOR2X1_86 gnd vdd FILL
XFILL_33_6_1 gnd vdd FILL
XFILL_32_1_0 gnd vdd FILL
XFILL_0_NOR3X1_18 gnd vdd FILL
XFILL_0_BUFX4_251 gnd vdd FILL
XOAI21X1_1401 XNOR2X1_90/Y BUFX4_290/Y OAI21X1_1401/C gnd OAI21X1_1401/Y vdd OAI21X1
XOAI21X1_1423 BUFX4_146/Y BUFX4_57/Y BUFX2_198/A gnd OAI21X1_1424/C vdd OAI21X1
XOAI21X1_1412 OAI21X1_1412/A BUFX4_290/Y OAI21X1_1412/C gnd OAI21X1_1412/Y vdd OAI21X1
XFILL_0_BUFX4_240 gnd vdd FILL
XFILL_1_OAI21X1_1621 gnd vdd FILL
XFILL_0_BUFX4_273 gnd vdd FILL
XOAI21X1_1434 BUFX4_127/Y BUFX4_41/Y BUFX2_202/A gnd OAI21X1_1435/C vdd OAI21X1
XOAI21X1_1456 BUFX4_159/Y BUFX4_67/Y BUFX2_211/A gnd OAI21X1_1457/C vdd OAI21X1
XFILL_1_OAI21X1_1632 gnd vdd FILL
XFILL_0_BUFX4_284 gnd vdd FILL
XNOR3X1_1 OR2X2_4/Y NOR3X1_1/B NOR3X1_1/C gnd NOR3X1_1/Y vdd NOR3X1
XOAI21X1_1445 INVX1_222/Y OAI21X1_1445/B OAI21X1_1445/C gnd OAI21X1_1445/Y vdd OAI21X1
XFILL_1_OAI21X1_1610 gnd vdd FILL
XFILL_0_BUFX4_262 gnd vdd FILL
XFILL_1_OAI21X1_1676 gnd vdd FILL
XFILL_1_OAI21X1_1665 gnd vdd FILL
XOAI21X1_1478 BUFX4_170/Y BUFX4_39/Y BUFX2_219/A gnd OAI21X1_1479/C vdd OAI21X1
XOAI21X1_1467 INVX2_109/Y INVX2_98/A INVX4_38/Y gnd OAI21X1_1468/C vdd OAI21X1
XFILL_0_BUFX4_295 gnd vdd FILL
XFILL_1_OAI21X1_1654 gnd vdd FILL
XFILL_4_NOR3X1_17 gnd vdd FILL
XFILL_1_OAI21X1_1643 gnd vdd FILL
XOAI21X1_1489 INVX1_223/A NOR2X1_154/A INVX2_77/Y gnd OAI21X1_1490/C vdd OAI21X1
XFILL_0_OAI21X1_412 gnd vdd FILL
XFILL_0_OAI21X1_401 gnd vdd FILL
XFILL_1_OAI21X1_1698 gnd vdd FILL
XFILL_1_OAI21X1_1687 gnd vdd FILL
XFILL_1_OAI21X1_627 gnd vdd FILL
XFILL_0_OAI21X1_456 gnd vdd FILL
XFILL_1_OAI21X1_605 gnd vdd FILL
XFILL_0_OAI21X1_445 gnd vdd FILL
XFILL_1_OAI21X1_616 gnd vdd FILL
XFILL_0_OAI21X1_423 gnd vdd FILL
XFILL_0_OAI21X1_434 gnd vdd FILL
XFILL_1_OAI21X1_649 gnd vdd FILL
XFILL_0_OAI21X1_478 gnd vdd FILL
XFILL_0_OAI21X1_489 gnd vdd FILL
XFILL_1_OAI21X1_638 gnd vdd FILL
XFILL_9_16_0 gnd vdd FILL
XFILL_0_OAI21X1_467 gnd vdd FILL
XFILL_3_DFFPOSX1_1020 gnd vdd FILL
XFILL_3_DFFPOSX1_1031 gnd vdd FILL
XFILL_13_14_1 gnd vdd FILL
XFILL_0_OAI21X1_1233 gnd vdd FILL
XFILL_0_OAI21X1_1222 gnd vdd FILL
XFILL_1_NAND2X1_633 gnd vdd FILL
XFILL_0_OAI21X1_1211 gnd vdd FILL
XFILL_0_NAND2X1_451 gnd vdd FILL
XFILL_0_NAND2X1_462 gnd vdd FILL
XFILL_0_OAI21X1_1200 gnd vdd FILL
XFILL_1_NAND2X1_611 gnd vdd FILL
XFILL_0_NAND2X1_440 gnd vdd FILL
XFILL_0_DFFPOSX1_801 gnd vdd FILL
XFILL_1_NAND2X1_666 gnd vdd FILL
XFILL_0_DFFPOSX1_812 gnd vdd FILL
XFILL_0_NAND2X1_473 gnd vdd FILL
XFILL_0_OAI21X1_1255 gnd vdd FILL
XFILL_0_NAND2X1_484 gnd vdd FILL
XFILL_0_NAND2X1_495 gnd vdd FILL
XFILL_0_DFFPOSX1_823 gnd vdd FILL
XFILL_0_DFFPOSX1_834 gnd vdd FILL
XFILL_0_OAI21X1_1244 gnd vdd FILL
XFILL_24_6_1 gnd vdd FILL
XFILL_2_OR2X2_8 gnd vdd FILL
XFILL_0_OAI21X1_1266 gnd vdd FILL
XFILL_1_NAND2X1_644 gnd vdd FILL
XFILL_1_NAND2X1_699 gnd vdd FILL
XFILL_0_DFFPOSX1_856 gnd vdd FILL
XFILL_0_OAI21X1_1299 gnd vdd FILL
XFILL_23_1_0 gnd vdd FILL
XFILL_0_OAI21X1_1288 gnd vdd FILL
XFILL_0_DFFPOSX1_867 gnd vdd FILL
XFILL_0_OAI21X1_1277 gnd vdd FILL
XFILL_0_DFFPOSX1_845 gnd vdd FILL
XFILL_0_DFFPOSX1_889 gnd vdd FILL
XFILL_0_DFFPOSX1_878 gnd vdd FILL
XDFFPOSX1_1008 BUFX2_675/A CLKBUF1_4/Y OAI21X1_1585/Y gnd vdd DFFPOSX1
XDFFPOSX1_1019 BUFX2_656/A CLKBUF1_57/Y OAI21X1_1596/Y gnd vdd DFFPOSX1
XFILL_5_DFFPOSX1_471 gnd vdd FILL
XFILL_5_DFFPOSX1_460 gnd vdd FILL
XFILL_5_DFFPOSX1_493 gnd vdd FILL
XFILL_5_DFFPOSX1_482 gnd vdd FILL
XFILL_0_AOI21X1_20 gnd vdd FILL
XFILL_0_AOI21X1_31 gnd vdd FILL
XFILL_0_AOI21X1_53 gnd vdd FILL
XFILL_0_AOI21X1_64 gnd vdd FILL
XFILL_0_AOI21X1_42 gnd vdd FILL
XFILL_0_OAI21X1_990 gnd vdd FILL
XFILL_18_13_1 gnd vdd FILL
XFILL_7_7_1 gnd vdd FILL
XFILL_6_2_0 gnd vdd FILL
XFILL_2_OAI21X1_1305 gnd vdd FILL
XFILL_31_15_1 gnd vdd FILL
XFILL_2_OAI21X1_1338 gnd vdd FILL
XFILL_2_DFFPOSX1_906 gnd vdd FILL
XFILL_2_DFFPOSX1_939 gnd vdd FILL
XFILL_2_DFFPOSX1_917 gnd vdd FILL
XFILL_2_OAI21X1_1349 gnd vdd FILL
XFILL_2_DFFPOSX1_928 gnd vdd FILL
XFILL_15_6_1 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XFILL_0_BUFX2_700 gnd vdd FILL
XFILL_3_XNOR2X1_19 gnd vdd FILL
XDFFPOSX1_309 BUFX2_978/A CLKBUF1_65/Y OAI21X1_235/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_722 gnd vdd FILL
XFILL_0_BUFX2_733 gnd vdd FILL
XFILL_0_NOR2X1_51 gnd vdd FILL
XFILL_0_BUFX2_711 gnd vdd FILL
XFILL_0_NOR2X1_40 gnd vdd FILL
XFILL_0_BUFX2_766 gnd vdd FILL
XFILL_0_BUFX2_744 gnd vdd FILL
XFILL_0_BUFX2_755 gnd vdd FILL
XFILL_0_NOR2X1_73 gnd vdd FILL
XFILL_0_NOR2X1_84 gnd vdd FILL
XFILL_1_DFFPOSX1_529 gnd vdd FILL
XFILL_1_DFFPOSX1_507 gnd vdd FILL
XFILL_1_DFFPOSX1_518 gnd vdd FILL
XFILL_0_NOR2X1_62 gnd vdd FILL
XFILL_0_BUFX2_788 gnd vdd FILL
XFILL_0_BUFX2_777 gnd vdd FILL
XFILL_6_DFFPOSX1_100 gnd vdd FILL
XFILL_0_NOR2X1_95 gnd vdd FILL
XFILL_0_BUFX2_799 gnd vdd FILL
XFILL_6_DFFPOSX1_133 gnd vdd FILL
XFILL_6_DFFPOSX1_111 gnd vdd FILL
XFILL_6_DFFPOSX1_122 gnd vdd FILL
XFILL_36_14_1 gnd vdd FILL
XFILL_3_DFFPOSX1_6 gnd vdd FILL
XBUFX4_330 BUFX4_381/A gnd BUFX4_330/Y vdd BUFX4
XBUFX4_363 BUFX4_380/A gnd BUFX4_363/Y vdd BUFX4
XFILL_30_10_0 gnd vdd FILL
XBUFX4_352 BUFX4_376/A gnd BUFX4_352/Y vdd BUFX4
XBUFX4_341 BUFX4_380/A gnd BUFX4_341/Y vdd BUFX4
XBUFX4_385 BUFX4_385/A gnd BUFX4_385/Y vdd BUFX4
XBUFX4_374 BUFX4_384/A gnd BUFX4_374/Y vdd BUFX4
XFILL_0_DFFPOSX1_119 gnd vdd FILL
XFILL_33_1 gnd vdd FILL
XFILL_0_DFFPOSX1_108 gnd vdd FILL
XOAI21X1_907 INVX1_108/Y BUFX4_184/Y OAI21X1_907/C gnd OAI21X1_907/Y vdd OAI21X1
XOAI21X1_929 BUFX4_143/Y INVX1_119/Y OAI21X1_929/C gnd OAI21X1_929/Y vdd OAI21X1
XFILL_0_NAND2X1_6 gnd vdd FILL
XOAI21X1_918 BUFX4_12/Y BUFX4_374/Y BUFX2_352/A gnd OAI21X1_919/C vdd OAI21X1
XOAI21X1_1231 OAI21X1_1231/A BUFX4_126/Y OAI21X1_1231/C gnd OAI21X1_1231/Y vdd OAI21X1
XOAI21X1_1220 OAI21X1_1220/A NOR2X1_177/Y OAI21X1_1220/C gnd OAI21X1_1220/Y vdd OAI21X1
XDFFPOSX1_821 BUFX2_70/A CLKBUF1_65/Y OAI21X1_1126/Y gnd vdd DFFPOSX1
XDFFPOSX1_810 BUFX2_77/A CLKBUF1_101/Y OAI21X1_1102/Y gnd vdd DFFPOSX1
XDFFPOSX1_832 BUFX2_82/A CLKBUF1_14/Y OAI21X1_1143/Y gnd vdd DFFPOSX1
XOAI21X1_1253 INVX2_105/Y NOR2X1_184/B OAI21X1_1253/C gnd OAI21X1_1255/A vdd OAI21X1
XOAI21X1_1242 INVX1_201/A INVX2_96/A INVX2_65/Y gnd OAI21X1_1243/C vdd OAI21X1
XFILL_1_OAI21X1_1440 gnd vdd FILL
XFILL_1_OAI21X1_1451 gnd vdd FILL
XOAI21X1_1264 NOR3X1_18/C INVX4_35/Y INVX1_173/Y gnd OAI21X1_1265/C vdd OAI21X1
XFILL_0_OAI21X1_231 gnd vdd FILL
XFILL_1_OAI21X1_1473 gnd vdd FILL
XFILL_1_OAI21X1_1462 gnd vdd FILL
XOAI21X1_1297 BUFX4_95/Y BUFX4_344/Y BUFX2_156/A gnd OAI21X1_1299/C vdd OAI21X1
XOAI21X1_1286 NOR2X1_194/B INVX1_207/A MUX2X1_2/S gnd OAI21X1_1287/B vdd OAI21X1
XDFFPOSX1_854 BUFX2_106/A CLKBUF1_36/Y OAI21X1_1174/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1484 gnd vdd FILL
XOAI21X1_1275 NOR2X1_193/B INVX1_174/Y INVX1_175/Y gnd NAND2X1_601/B vdd OAI21X1
XFILL_0_OAI21X1_220 gnd vdd FILL
XDFFPOSX1_843 BUFX2_94/A CLKBUF1_62/Y OAI21X1_1159/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_402 gnd vdd FILL
XDFFPOSX1_865 BUFX2_118/A CLKBUF1_20/Y OAI21X1_1195/Y gnd vdd DFFPOSX1
XDFFPOSX1_887 BUFX2_136/A CLKBUF1_65/Y OAI21X1_1251/Y gnd vdd DFFPOSX1
XDFFPOSX1_876 BUFX2_163/A CLKBUF1_101/Y OAI21X1_1217/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_253 gnd vdd FILL
XDFFPOSX1_898 BUFX2_148/A CLKBUF1_55/Y OAI21X1_1282/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_242 gnd vdd FILL
XFILL_1_OAI21X1_1495 gnd vdd FILL
XINVX2_26 bundleStartMajId_i[26] gnd INVX2_26/Y vdd INVX2
XFILL_1_OAI21X1_424 gnd vdd FILL
XINVX2_15 bundleStartMajId_i[53] gnd INVX2_15/Y vdd INVX2
XFILL_1_OAI21X1_413 gnd vdd FILL
XFILL_0_OAI21X1_264 gnd vdd FILL
XFILL_1_OAI21X1_435 gnd vdd FILL
XFILL_0_OAI21X1_297 gnd vdd FILL
XFILL_0_OAI21X1_275 gnd vdd FILL
XINVX2_59 bundleAddress_i[57] gnd INVX2_59/Y vdd INVX2
XFILL_0_OAI21X1_286 gnd vdd FILL
XINVX2_37 bundleStartMajId_i[7] gnd INVX2_37/Y vdd INVX2
XFILL_1_OAI21X1_457 gnd vdd FILL
XFILL_1_OAI21X1_446 gnd vdd FILL
XINVX2_48 INVX2_48/A gnd INVX2_48/Y vdd INVX2
XFILL_1_OAI21X1_468 gnd vdd FILL
XFILL_1_OAI21X1_479 gnd vdd FILL
XFILL_1_INVX4_37 gnd vdd FILL
XFILL_1_INVX4_15 gnd vdd FILL
XFILL_0_OAI21X1_1030 gnd vdd FILL
XFILL_0_OAI21X1_1041 gnd vdd FILL
XFILL_1_NAND2X1_430 gnd vdd FILL
XFILL_1_NAND2X1_441 gnd vdd FILL
XFILL_0_NAND2X1_270 gnd vdd FILL
XFILL_1_BUFX4_216 gnd vdd FILL
XFILL_1_BUFX4_205 gnd vdd FILL
XFILL_1_BUFX4_227 gnd vdd FILL
XFILL_0_OAI21X1_1052 gnd vdd FILL
XFILL_0_OAI21X1_1063 gnd vdd FILL
XFILL_0_DFFPOSX1_642 gnd vdd FILL
XFILL_0_NAND2X1_292 gnd vdd FILL
XFILL_1_NAND2X1_463 gnd vdd FILL
XFILL_0_NAND2X1_281 gnd vdd FILL
XFILL_0_DFFPOSX1_620 gnd vdd FILL
XFILL_0_DFFPOSX1_631 gnd vdd FILL
XFILL_0_OAI21X1_1074 gnd vdd FILL
XFILL_1_NAND2X1_452 gnd vdd FILL
XFILL_0_DFFPOSX1_664 gnd vdd FILL
XFILL_1_BUFX4_249 gnd vdd FILL
XFILL_1_NAND2X1_485 gnd vdd FILL
XFILL_1_NAND2X1_496 gnd vdd FILL
XFILL_0_OAI21X1_1085 gnd vdd FILL
XFILL_1_BUFX4_238 gnd vdd FILL
XFILL_0_OAI21X1_1096 gnd vdd FILL
XFILL_0_DFFPOSX1_675 gnd vdd FILL
XFILL_0_DFFPOSX1_653 gnd vdd FILL
XFILL_0_DFFPOSX1_697 gnd vdd FILL
XFILL_0_DFFPOSX1_686 gnd vdd FILL
XFILL_5_DFFPOSX1_290 gnd vdd FILL
XFILL_2_XNOR2X1_9 gnd vdd FILL
XFILL_1_OAI21X1_991 gnd vdd FILL
XFILL_1_OAI21X1_980 gnd vdd FILL
XFILL_2_BUFX4_98 gnd vdd FILL
XBUFX2_801 BUFX2_801/A gnd tid1_o[33] vdd BUFX2
XFILL_2_DFFPOSX1_714 gnd vdd FILL
XFILL_2_DFFPOSX1_703 gnd vdd FILL
XBUFX2_812 BUFX2_812/A gnd tid1_o[23] vdd BUFX2
XFILL_2_OAI21X1_1135 gnd vdd FILL
XBUFX2_845 BUFX2_845/A gnd tid2_o[51] vdd BUFX2
XBUFX2_823 BUFX2_823/A gnd tid1_o[13] vdd BUFX2
XFILL_2_DFFPOSX1_747 gnd vdd FILL
XFILL_2_DFFPOSX1_725 gnd vdd FILL
XFILL_2_DFFPOSX1_736 gnd vdd FILL
XFILL_2_OAI21X1_1168 gnd vdd FILL
XBUFX2_834 NAND2X1_4/A gnd tid1_o[3] vdd BUFX2
XFILL_2_DFFPOSX1_758 gnd vdd FILL
XBUFX2_856 BUFX2_856/A gnd tid2_o[41] vdd BUFX2
XFILL_2_DFFPOSX1_769 gnd vdd FILL
XBUFX2_867 BUFX2_867/A gnd tid2_o[31] vdd BUFX2
XBUFX2_889 BUFX2_889/A gnd tid2_o[11] vdd BUFX2
XBUFX2_878 BUFX2_878/A gnd tid2_o[21] vdd BUFX2
XFILL_0_NOR2X1_218 gnd vdd FILL
XFILL_0_NOR2X1_207 gnd vdd FILL
XFILL_0_NOR2X1_229 gnd vdd FILL
XFILL_30_4_1 gnd vdd FILL
XFILL_3_CLKBUF1_9 gnd vdd FILL
XDFFPOSX1_117 BUFX2_786/A CLKBUF1_59/Y OAI21X1_1791/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_304 gnd vdd FILL
XDFFPOSX1_106 BUFX2_833/A CLKBUF1_49/Y OAI21X1_1780/Y gnd vdd DFFPOSX1
XDFFPOSX1_128 BUFX2_798/A CLKBUF1_81/Y OAI21X1_1802/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_530 gnd vdd FILL
XFILL_0_BUFX2_541 gnd vdd FILL
XFILL_1_DFFPOSX1_337 gnd vdd FILL
XFILL_1_DFFPOSX1_326 gnd vdd FILL
XFILL_1_DFFPOSX1_315 gnd vdd FILL
XFILL_0_BUFX2_574 gnd vdd FILL
XDFFPOSX1_139 BUFX2_810/A CLKBUF1_67/Y OAI21X1_1813/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_563 gnd vdd FILL
XFILL_0_BUFX2_552 gnd vdd FILL
XFILL_1_DFFPOSX1_348 gnd vdd FILL
XFILL_0_BUFX2_596 gnd vdd FILL
XFILL_0_BUFX2_585 gnd vdd FILL
XFILL_1_DFFPOSX1_359 gnd vdd FILL
XNAND2X1_209 bundleStartMajId_i[31] bundleStartMajId_i[28] gnd NOR2X1_31/B vdd NAND2X1
XFILL_4_DFFPOSX1_808 gnd vdd FILL
XFILL_4_DFFPOSX1_819 gnd vdd FILL
XFILL_38_5_1 gnd vdd FILL
XFILL_37_0_0 gnd vdd FILL
XFILL_4_CLKBUF1_42 gnd vdd FILL
XFILL_4_CLKBUF1_31 gnd vdd FILL
XBUFX4_171 BUFX4_17/Y gnd BUFX4_171/Y vdd BUFX4
XBUFX4_160 BUFX4_15/Y gnd BUFX4_160/Y vdd BUFX4
XFILL_4_CLKBUF1_20 gnd vdd FILL
XFILL_0_INVX1_60 gnd vdd FILL
XBUFX4_182 BUFX4_20/Y gnd BUFX4_182/Y vdd BUFX4
XFILL_0_INVX1_93 gnd vdd FILL
XBUFX4_193 BUFX4_23/Y gnd BUFX4_193/Y vdd BUFX4
XFILL_4_CLKBUF1_86 gnd vdd FILL
XFILL_4_CLKBUF1_64 gnd vdd FILL
XNOR2X1_220 NOR2X1_220/A NOR2X1_220/B gnd INVX4_51/A vdd NOR2X1
XFILL_0_INVX1_82 gnd vdd FILL
XFILL_0_INVX1_71 gnd vdd FILL
XNOR2X1_231 OR2X2_21/B OR2X2_21/A gnd NOR2X1_231/Y vdd NOR2X1
XFILL_4_CLKBUF1_53 gnd vdd FILL
XFILL_0_BUFX2_24 gnd vdd FILL
XFILL_0_BUFX2_13 gnd vdd FILL
XFILL_0_BUFX2_35 gnd vdd FILL
XFILL_4_CLKBUF1_97 gnd vdd FILL
XFILL_0_BUFX2_68 gnd vdd FILL
XFILL_0_BUFX2_57 gnd vdd FILL
XFILL_0_BUFX2_46 gnd vdd FILL
XFILL_1_NOR2X1_27 gnd vdd FILL
XFILL_1_NOR2X1_16 gnd vdd FILL
XFILL_0_BUFX2_79 gnd vdd FILL
XOAI21X1_715 OAI21X1_715/A BUFX4_289/Y OAI21X1_715/C gnd OAI21X1_715/Y vdd OAI21X1
XFILL_21_4_1 gnd vdd FILL
XFILL_1_NOR2X1_49 gnd vdd FILL
XOAI21X1_704 NOR2X1_11/B NOR2X1_105/A INVX2_17/Y gnd OAI21X1_704/Y vdd OAI21X1
XOAI21X1_737 BUFX4_147/Y BUFX4_77/Y BUFX2_605/A gnd OAI21X1_738/C vdd OAI21X1
XFILL_3_DFFPOSX1_409 gnd vdd FILL
XOAI21X1_748 NOR3X1_9/C NOR3X1_9/A OR2X2_15/B gnd OAI21X1_748/Y vdd OAI21X1
XOAI21X1_726 XNOR2X1_45/Y BUFX4_300/Y OAI21X1_726/C gnd OAI21X1_726/Y vdd OAI21X1
XOAI21X1_759 XNOR2X1_49/Y BUFX4_300/Y OAI21X1_759/C gnd OAI21X1_759/Y vdd OAI21X1
XFILL_21_15_0 gnd vdd FILL
XDFFPOSX1_640 INVX1_69/A CLKBUF1_99/Y OAI21X1_868/Y gnd vdd DFFPOSX1
XOAI21X1_1050 BUFX4_340/Y INVX2_66/Y NAND2X1_416/Y gnd OAI21X1_1050/Y vdd OAI21X1
XOAI21X1_1061 OAI21X1_5/A INVX4_37/Y NAND2X1_427/Y gnd OAI21X1_1061/Y vdd OAI21X1
XOAI21X1_1072 BUFX4_370/Y INVX2_77/Y NAND2X1_438/Y gnd OAI21X1_1072/Y vdd OAI21X1
XDFFPOSX1_662 BUFX2_299/A CLKBUF1_39/Y OAI21X1_890/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1292 gnd vdd FILL
XOAI21X1_1083 BUFX4_339/Y INVX2_82/Y NAND2X1_449/Y gnd OAI21X1_1083/Y vdd OAI21X1
XFILL_1_OAI21X1_1281 gnd vdd FILL
XOAI21X1_1094 BUFX4_330/Y INVX2_89/Y NAND2X1_460/Y gnd OAI21X1_1094/Y vdd OAI21X1
XDFFPOSX1_651 BUFX2_316/A CLKBUF1_32/Y OAI21X1_879/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1270 gnd vdd FILL
XDFFPOSX1_673 BUFX2_311/A CLKBUF1_82/Y OAI21X1_901/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_210 gnd vdd FILL
XDFFPOSX1_684 BUFX2_351/A CLKBUF1_37/Y OAI21X1_917/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_860 gnd vdd FILL
XNAND2X1_710 BUFX2_702/A BUFX4_197/Y gnd NAND2X1_710/Y vdd NAND2X1
XFILL_1_DFFPOSX1_882 gnd vdd FILL
XFILL_1_OAI21X1_232 gnd vdd FILL
XFILL_1_OAI21X1_243 gnd vdd FILL
XNAND2X1_721 BUFX2_833/A BUFX4_344/Y gnd NAND2X1_721/Y vdd NAND2X1
XFILL_1_DFFPOSX1_871 gnd vdd FILL
XDFFPOSX1_695 BUFX2_332/A CLKBUF1_40/Y OAI21X1_939/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_893 gnd vdd FILL
XFILL_1_OAI21X1_221 gnd vdd FILL
XFILL_2_OAI21X1_414 gnd vdd FILL
XFILL_2_OAI21X1_403 gnd vdd FILL
XFILL_0_NOR2X1_4 gnd vdd FILL
XFILL_1_OAI21X1_254 gnd vdd FILL
XNAND2X1_732 BUFX2_786/A BUFX4_385/Y gnd NAND2X1_732/Y vdd NAND2X1
XFILL_1_OAI21X1_276 gnd vdd FILL
XFILL_1_OAI21X1_287 gnd vdd FILL
XNAND2X1_754 BUFX2_810/A BUFX4_375/Y gnd NAND2X1_754/Y vdd NAND2X1
XFILL_2_OAI21X1_458 gnd vdd FILL
XNAND2X1_743 BUFX2_798/A BUFX4_343/Y gnd NAND2X1_743/Y vdd NAND2X1
XFILL_1_OAI21X1_265 gnd vdd FILL
XFILL_2_OAI21X1_425 gnd vdd FILL
XNAND2X1_765 BUFX2_823/A BUFX4_359/Y gnd NAND2X1_765/Y vdd NAND2X1
XFILL_1_OAI21X1_298 gnd vdd FILL
XBUFX2_108 BUFX2_108/A gnd addr2_o[15] vdd BUFX2
XFILL_29_5_1 gnd vdd FILL
XFILL_28_0_0 gnd vdd FILL
XFILL_2_XNOR2X1_38 gnd vdd FILL
XFILL_2_XNOR2X1_16 gnd vdd FILL
XFILL_2_XNOR2X1_27 gnd vdd FILL
XFILL_4_5_1 gnd vdd FILL
XBUFX2_119 BUFX2_119/A gnd addr2_o[5] vdd BUFX2
XFILL_2_XNOR2X1_49 gnd vdd FILL
XFILL_3_0_0 gnd vdd FILL
XFILL_0_DFFPOSX1_450 gnd vdd FILL
XFILL_1_NAND2X1_260 gnd vdd FILL
XFILL_1_NAND2X1_271 gnd vdd FILL
XFILL_0_DFFPOSX1_483 gnd vdd FILL
XFILL_26_14_0 gnd vdd FILL
XINVX8_2 INVX8_2/A gnd INVX8_2/Y vdd INVX8
XFILL_0_DFFPOSX1_461 gnd vdd FILL
XFILL_12_4_1 gnd vdd FILL
XFILL_2_DFFPOSX1_3 gnd vdd FILL
XFILL_0_DFFPOSX1_494 gnd vdd FILL
XFILL_0_DFFPOSX1_472 gnd vdd FILL
XFILL_3_DFFPOSX1_932 gnd vdd FILL
XFILL_3_DFFPOSX1_921 gnd vdd FILL
XFILL_3_DFFPOSX1_910 gnd vdd FILL
XFILL_3_DFFPOSX1_954 gnd vdd FILL
XFILL_3_DFFPOSX1_943 gnd vdd FILL
XFILL_3_DFFPOSX1_965 gnd vdd FILL
XFILL_3_DFFPOSX1_998 gnd vdd FILL
XFILL_3_DFFPOSX1_987 gnd vdd FILL
XFILL_3_DFFPOSX1_976 gnd vdd FILL
XBUFX4_11 BUFX4_11/A gnd BUFX4_11/Y vdd BUFX4
XBUFX4_44 BUFX4_82/A gnd BUFX4_44/Y vdd BUFX4
XBUFX4_22 BUFX4_26/A gnd BUFX4_22/Y vdd BUFX4
XBUFX4_33 BUFX4_82/A gnd BUFX4_33/Y vdd BUFX4
XBUFX4_55 BUFX4_55/A gnd BUFX4_55/Y vdd BUFX4
XBUFX4_77 BUFX4_82/A gnd BUFX4_77/Y vdd BUFX4
XBUFX4_66 BUFX4_66/A gnd BUFX4_66/Y vdd BUFX4
XBUFX2_620 BUFX2_620/A gnd majID4_o[23] vdd BUFX2
XFILL_19_0_0 gnd vdd FILL
XBUFX4_99 BUFX4_6/A gnd BUFX4_99/Y vdd BUFX4
XBUFX4_88 clock_i gnd BUFX4_88/Y vdd BUFX4
XFILL_2_DFFPOSX1_500 gnd vdd FILL
XFILL_2_DFFPOSX1_522 gnd vdd FILL
XFILL_2_DFFPOSX1_511 gnd vdd FILL
XBUFX2_664 BUFX2_664/A gnd pid1_o[9] vdd BUFX2
XFILL_2_DFFPOSX1_544 gnd vdd FILL
XBUFX2_631 BUFX2_631/A gnd majID4_o[13] vdd BUFX2
XFILL_2_DFFPOSX1_555 gnd vdd FILL
XBUFX2_653 BUFX2_653/A gnd pid1_o[19] vdd BUFX2
XFILL_2_DFFPOSX1_533 gnd vdd FILL
XFILL_1_15_0 gnd vdd FILL
XBUFX2_642 BUFX2_642/A gnd majID4_o[3] vdd BUFX2
XBUFX2_697 BUFX2_697/A gnd pid2_o[8] vdd BUFX2
XFILL_2_DFFPOSX1_599 gnd vdd FILL
XFILL_2_DFFPOSX1_588 gnd vdd FILL
XFILL_2_DFFPOSX1_566 gnd vdd FILL
XBUFX2_675 BUFX2_675/A gnd pid1_o[27] vdd BUFX2
XFILL_2_DFFPOSX1_577 gnd vdd FILL
XBUFX2_686 BUFX2_686/A gnd pid2_o[18] vdd BUFX2
XOR2X2_14 OR2X2_14/A bundleStartMajId_i[0] gnd OR2X2_14/Y vdd OR2X2
XFILL_1_DFFPOSX1_112 gnd vdd FILL
XFILL_1_DFFPOSX1_101 gnd vdd FILL
XINVX2_160 bundleTid_i[49] gnd INVX2_160/Y vdd INVX2
XINVX2_193 bundleTid_i[16] gnd INVX2_193/Y vdd INVX2
XFILL_1_DFFPOSX1_134 gnd vdd FILL
XFILL_1_DFFPOSX1_156 gnd vdd FILL
XINVX2_171 bundleTid_i[38] gnd INVX2_171/Y vdd INVX2
XFILL_1_DFFPOSX1_145 gnd vdd FILL
XINVX2_182 bundleTid_i[27] gnd INVX2_182/Y vdd INVX2
XFILL_1_DFFPOSX1_123 gnd vdd FILL
XFILL_2_AOI21X1_27 gnd vdd FILL
XFILL_0_BUFX2_382 gnd vdd FILL
XOR2X2_7 OR2X2_7/A bundleStartMajId_i[31] gnd OR2X2_7/Y vdd OR2X2
XFILL_0_BUFX2_393 gnd vdd FILL
XFILL_0_BUFX2_360 gnd vdd FILL
XFILL_0_BUFX2_371 gnd vdd FILL
XFILL_1_DFFPOSX1_178 gnd vdd FILL
XFILL_1_DFFPOSX1_189 gnd vdd FILL
XXNOR2X1_9 XNOR2X1_9/A INVX4_9/Y gnd XNOR2X1_9/Y vdd XNOR2X1
XFILL_1_DFFPOSX1_167 gnd vdd FILL
XFILL_4_DFFPOSX1_627 gnd vdd FILL
XFILL_4_DFFPOSX1_605 gnd vdd FILL
XFILL_4_DFFPOSX1_616 gnd vdd FILL
XFILL_6_14_0 gnd vdd FILL
XFILL_4_DFFPOSX1_649 gnd vdd FILL
XFILL_4_DFFPOSX1_638 gnd vdd FILL
XFILL_10_12_1 gnd vdd FILL
XFILL_1_BUFX2_517 gnd vdd FILL
XFILL_1_BUFX2_528 gnd vdd FILL
XFILL_1_BUFX2_539 gnd vdd FILL
XOAI21X1_501 BUFX4_176/Y INVX4_1/Y OAI21X1_501/C gnd OAI21X1_501/Y vdd OAI21X1
XOAI21X1_523 BUFX4_7/A BUFX4_388/Y BUFX2_583/A gnd OAI21X1_524/C vdd OAI21X1
XOAI21X1_512 OAI21X1_512/A BUFX4_163/Y OAI21X1_512/C gnd OAI21X1_512/Y vdd OAI21X1
XINVX1_9 OR2X2_1/A gnd INVX1_9/Y vdd INVX1
XFILL_3_DFFPOSX1_217 gnd vdd FILL
XFILL_3_DFFPOSX1_228 gnd vdd FILL
XOAI21X1_556 OAI21X1_556/A BUFX4_175/Y OAI21X1_556/C gnd OAI21X1_556/Y vdd OAI21X1
XOAI21X1_534 OAI21X1_534/A BUFX4_122/Y OAI21X1_534/C gnd OAI21X1_534/Y vdd OAI21X1
XOAI21X1_545 XNOR2X1_27/A INVX4_6/Y INVX2_17/Y gnd OAI21X1_545/Y vdd OAI21X1
XFILL_3_DFFPOSX1_206 gnd vdd FILL
XFILL_3_DFFPOSX1_239 gnd vdd FILL
XOAI21X1_567 XNOR2X1_32/Y BUFX4_147/Y OAI21X1_567/C gnd OAI21X1_567/Y vdd OAI21X1
XOAI21X1_578 XNOR2X1_33/Y BUFX4_174/Y OAI21X1_578/C gnd OAI21X1_578/Y vdd OAI21X1
XOAI21X1_589 BUFX4_9/Y BUFX4_335/Y BUFX2_549/A gnd OAI21X1_590/C vdd OAI21X1
XDFFPOSX1_470 BUFX2_503/A CLKBUF1_100/Y OAI21X1_477/Y gnd vdd DFFPOSX1
XDFFPOSX1_481 BUFX2_515/A CLKBUF1_19/Y OAI21X1_496/Y gnd vdd DFFPOSX1
XDFFPOSX1_492 BUFX2_583/A CLKBUF1_46/Y OAI21X1_524/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_690 gnd vdd FILL
XFILL_2_OAI21X1_233 gnd vdd FILL
XFILL_2_OAI21X1_266 gnd vdd FILL
XNAND2X1_551 BUFX2_103/A BUFX4_202/Y gnd NAND2X1_551/Y vdd NAND2X1
XNAND2X1_562 BUFX2_109/A BUFX4_187/Y gnd NAND2X1_562/Y vdd NAND2X1
XNAND2X1_540 bundleAddress_i[28] bundleAddress_i[27] gnd INVX1_208/A vdd NAND2X1
XNAND2X1_595 bundleAddress_i[49] NOR2X1_183/Y gnd NOR2X1_184/B vdd NAND2X1
XNAND2X1_584 BUFX2_122/A BUFX4_187/Y gnd NAND2X1_584/Y vdd NAND2X1
XFILL_15_11_1 gnd vdd FILL
XNAND2X1_573 BUFX2_114/A BUFX4_201/Y gnd NAND2X1_573/Y vdd NAND2X1
XFILL_0_AND2X2_30 gnd vdd FILL
XFILL_1_DFFPOSX1_1019 gnd vdd FILL
XFILL_1_DFFPOSX1_1008 gnd vdd FILL
XFILL_0_DFFPOSX1_291 gnd vdd FILL
XFILL_0_DFFPOSX1_280 gnd vdd FILL
XOAI21X1_1808 BUFX4_316/Y INVX2_180/Y NAND2X1_749/Y gnd OAI21X1_1808/Y vdd OAI21X1
XOAI21X1_1819 BUFX4_316/Y INVX2_191/Y NAND2X1_760/Y gnd OAI21X1_1819/Y vdd OAI21X1
XFILL_3_DFFPOSX1_740 gnd vdd FILL
XFILL_3_DFFPOSX1_751 gnd vdd FILL
XFILL_3_DFFPOSX1_773 gnd vdd FILL
XFILL_3_DFFPOSX1_762 gnd vdd FILL
XFILL_3_CLKBUF1_50 gnd vdd FILL
XFILL_3_CLKBUF1_61 gnd vdd FILL
XFILL_0_OAI21X1_808 gnd vdd FILL
XFILL_3_CLKBUF1_72 gnd vdd FILL
XFILL_3_CLKBUF1_83 gnd vdd FILL
XFILL_0_OAI21X1_819 gnd vdd FILL
XFILL_3_CLKBUF1_94 gnd vdd FILL
XFILL_3_DFFPOSX1_784 gnd vdd FILL
XFILL_3_DFFPOSX1_795 gnd vdd FILL
XFILL_33_12_1 gnd vdd FILL
XFILL_2_DFFPOSX1_330 gnd vdd FILL
XFILL_0_OAI21X1_1607 gnd vdd FILL
XFILL_0_OAI21X1_1629 gnd vdd FILL
XFILL_35_3_1 gnd vdd FILL
XFILL_2_DFFPOSX1_341 gnd vdd FILL
XBUFX2_450 BUFX2_450/A gnd majID1_o[3] vdd BUFX2
XFILL_2_DFFPOSX1_374 gnd vdd FILL
XFILL_0_OAI21X1_1618 gnd vdd FILL
XFILL_2_DFFPOSX1_352 gnd vdd FILL
XBUFX2_472 BUFX2_472/A gnd majID2_o[41] vdd BUFX2
XBUFX2_461 BUFX2_461/A gnd majID2_o[51] vdd BUFX2
XFILL_2_DFFPOSX1_363 gnd vdd FILL
XBUFX2_494 BUFX2_494/A gnd majID2_o[21] vdd BUFX2
XFILL_2_DFFPOSX1_396 gnd vdd FILL
XFILL_2_DFFPOSX1_385 gnd vdd FILL
XBUFX2_483 BUFX2_483/A gnd majID2_o[31] vdd BUFX2
XFILL_5_DFFPOSX1_812 gnd vdd FILL
XFILL_5_DFFPOSX1_801 gnd vdd FILL
XFILL_5_DFFPOSX1_823 gnd vdd FILL
XFILL_5_DFFPOSX1_834 gnd vdd FILL
XFILL_5_DFFPOSX1_845 gnd vdd FILL
XFILL_5_DFFPOSX1_889 gnd vdd FILL
XFILL_5_DFFPOSX1_878 gnd vdd FILL
XFILL_5_DFFPOSX1_856 gnd vdd FILL
XFILL_5_DFFPOSX1_867 gnd vdd FILL
XFILL_1_XNOR2X1_13 gnd vdd FILL
XFILL_1_XNOR2X1_46 gnd vdd FILL
XFILL_1_XNOR2X1_35 gnd vdd FILL
XFILL_1_XNOR2X1_24 gnd vdd FILL
XFILL_1_XNOR2X1_57 gnd vdd FILL
XFILL_1_XNOR2X1_79 gnd vdd FILL
XFILL_1_XNOR2X1_68 gnd vdd FILL
XFILL_2_OAI21X1_90 gnd vdd FILL
XFILL_0_BUFX2_190 gnd vdd FILL
XFILL_38_11_1 gnd vdd FILL
XFILL_4_DFFPOSX1_402 gnd vdd FILL
XFILL_4_DFFPOSX1_413 gnd vdd FILL
XFILL_4_DFFPOSX1_424 gnd vdd FILL
XFILL_4_DFFPOSX1_435 gnd vdd FILL
XFILL_4_DFFPOSX1_446 gnd vdd FILL
XFILL_4_DFFPOSX1_479 gnd vdd FILL
XFILL_4_DFFPOSX1_468 gnd vdd FILL
XFILL_4_DFFPOSX1_457 gnd vdd FILL
XFILL_26_3_1 gnd vdd FILL
XFILL_1_3_1 gnd vdd FILL
XFILL_1_BUFX2_325 gnd vdd FILL
XFILL_1_BUFX2_336 gnd vdd FILL
XFILL_1_BUFX2_314 gnd vdd FILL
XFILL_1_BUFX2_369 gnd vdd FILL
XOAI21X1_320 BUFX4_174/Y BUFX4_79/Y BUFX2_1026/A gnd OAI21X1_321/C vdd OAI21X1
XOAI21X1_331 BUFX4_321/Y INVX2_10/Y NAND2X1_75/Y gnd OAI21X1_331/Y vdd OAI21X1
XOAI21X1_364 BUFX4_351/Y INVX4_17/Y OAI21X1_364/C gnd OAI21X1_364/Y vdd OAI21X1
XOAI21X1_353 BUFX4_378/Y INVX4_11/Y NAND2X1_97/Y gnd OAI21X1_353/Y vdd OAI21X1
XOAI21X1_342 BUFX4_335/Y NOR2X1_9/A NAND2X1_86/Y gnd OAI21X1_342/Y vdd OAI21X1
XOAI21X1_386 BUFX4_328/Y INVX4_26/Y OAI21X1_386/C gnd OAI21X1_386/Y vdd OAI21X1
XOAI21X1_375 BUFX4_362/Y INVX2_32/Y OAI21X1_375/C gnd OAI21X1_375/Y vdd OAI21X1
XOAI21X1_397 INVX1_24/A INVX4_1/Y INVX2_10/Y gnd OAI21X1_398/C vdd OAI21X1
XAND2X2_9 NOR3X1_2/Y bundleStartMajId_i[18] gnd AND2X2_9/Y vdd AND2X2
XFILL_6_DFFPOSX1_507 gnd vdd FILL
XFILL_6_DFFPOSX1_518 gnd vdd FILL
XFILL_6_DFFPOSX1_529 gnd vdd FILL
XFILL_9_4_1 gnd vdd FILL
XNAND2X1_370 BUFX2_293/A BUFX4_180/Y gnd OAI21X1_876/C vdd NAND2X1
XNAND2X1_381 BUFX2_296/A BUFX4_232/Y gnd OAI21X1_887/C vdd NAND2X1
XNAND2X1_392 BUFX2_308/A BUFX4_220/Y gnd OAI21X1_898/C vdd NAND2X1
XFILL_4_DFFPOSX1_980 gnd vdd FILL
XFILL_0_INVX1_102 gnd vdd FILL
XFILL_0_INVX1_113 gnd vdd FILL
XFILL_4_DFFPOSX1_991 gnd vdd FILL
XFILL_1_AOI21X1_24 gnd vdd FILL
XFILL_1_AOI21X1_13 gnd vdd FILL
XFILL_17_3_1 gnd vdd FILL
XFILL_0_INVX1_124 gnd vdd FILL
XFILL_0_INVX1_146 gnd vdd FILL
XFILL_0_INVX1_135 gnd vdd FILL
XFILL_1_AOI21X1_46 gnd vdd FILL
XFILL_1_AOI21X1_35 gnd vdd FILL
XFILL_0_INVX1_179 gnd vdd FILL
XFILL_0_INVX1_157 gnd vdd FILL
XFILL_1_AOI21X1_57 gnd vdd FILL
XFILL_0_INVX1_168 gnd vdd FILL
XFILL_5_DFFPOSX1_108 gnd vdd FILL
XFILL_5_DFFPOSX1_119 gnd vdd FILL
XFILL_1_INVX2_70 gnd vdd FILL
XFILL_1_BUFX2_881 gnd vdd FILL
XFILL_1_BUFX2_892 gnd vdd FILL
XFILL_2_NOR3X1_1 gnd vdd FILL
XOAI21X1_1605 OAI21X1_4/A INVX2_141/Y NAND2X1_674/Y gnd OAI21X1_1605/Y vdd OAI21X1
XOAI21X1_1616 INVX2_119/Y BUFX4_227/Y NAND2X1_684/Y gnd DFFPOSX1_6/D vdd OAI21X1
XFILL_1_OAI21X1_1825 gnd vdd FILL
XOAI21X1_1627 INVX2_130/Y INVX8_1/A NAND2X1_695/Y gnd DFFPOSX1_17/D vdd OAI21X1
XFILL_1_OAI21X1_1803 gnd vdd FILL
XOAI21X1_1638 INVX2_141/Y BUFX4_192/Y NAND2X1_706/Y gnd DFFPOSX1_28/D vdd OAI21X1
XFILL_1_OAI21X1_1814 gnd vdd FILL
XOAI21X1_1649 BUFX4_150/Y INVX2_118/Y OAI21X1_1649/C gnd DFFPOSX1_37/D vdd OAI21X1
XFILL_0_OAI21X1_605 gnd vdd FILL
XFILL_3_DFFPOSX1_592 gnd vdd FILL
XFILL_3_DFFPOSX1_570 gnd vdd FILL
XFILL_3_DFFPOSX1_581 gnd vdd FILL
XFILL_1_OAI21X1_809 gnd vdd FILL
XFILL_0_OAI21X1_627 gnd vdd FILL
XFILL_0_OAI21X1_638 gnd vdd FILL
XFILL_0_OAI21X1_616 gnd vdd FILL
XFILL_0_OAI21X1_649 gnd vdd FILL
XFILL_1_AND2X2_17 gnd vdd FILL
XFILL_1_AND2X2_28 gnd vdd FILL
XFILL_0_NAND2X1_600 gnd vdd FILL
XFILL_0_NAND2X1_611 gnd vdd FILL
XFILL_0_OAI21X1_1415 gnd vdd FILL
XFILL_0_OAI21X1_1404 gnd vdd FILL
XFILL_0_NAND2X1_633 gnd vdd FILL
XFILL_0_NAND2X1_622 gnd vdd FILL
XFILL_0_NAND2X1_644 gnd vdd FILL
XFILL_0_NAND2X1_666 gnd vdd FILL
XFILL_0_NAND2X1_677 gnd vdd FILL
XFILL_0_OAI21X1_1437 gnd vdd FILL
XFILL_0_OAI21X1_1426 gnd vdd FILL
XFILL_2_DFFPOSX1_171 gnd vdd FILL
XFILL_2_DFFPOSX1_182 gnd vdd FILL
XBUFX2_280 INVX1_71/A gnd instr1_o[5] vdd BUFX2
XFILL_0_OAI21X1_1448 gnd vdd FILL
XFILL_2_DFFPOSX1_160 gnd vdd FILL
XFILL_0_NAND2X1_655 gnd vdd FILL
XFILL_0_NAND2X1_699 gnd vdd FILL
XBUFX2_291 INVX1_53/A gnd instr1_o[23] vdd BUFX2
XFILL_0_OAI21X1_1459 gnd vdd FILL
XFILL_2_DFFPOSX1_193 gnd vdd FILL
XFILL_0_NAND2X1_688 gnd vdd FILL
XFILL_5_DFFPOSX1_620 gnd vdd FILL
XFILL_5_DFFPOSX1_664 gnd vdd FILL
XFILL_5_DFFPOSX1_642 gnd vdd FILL
XFILL_5_DFFPOSX1_631 gnd vdd FILL
XFILL_5_DFFPOSX1_653 gnd vdd FILL
XFILL_24_17_1 gnd vdd FILL
XFILL_5_DFFPOSX1_675 gnd vdd FILL
XFILL_5_DFFPOSX1_697 gnd vdd FILL
XFILL_5_DFFPOSX1_686 gnd vdd FILL
XFILL_4_DFFPOSX1_221 gnd vdd FILL
XFILL_4_DFFPOSX1_210 gnd vdd FILL
XFILL_4_DFFPOSX1_232 gnd vdd FILL
XFILL_4_DFFPOSX1_254 gnd vdd FILL
XFILL_4_DFFPOSX1_243 gnd vdd FILL
XFILL_2_OAI21X1_1509 gnd vdd FILL
XFILL_4_DFFPOSX1_276 gnd vdd FILL
XFILL_4_DFFPOSX1_265 gnd vdd FILL
XFILL_4_DFFPOSX1_287 gnd vdd FILL
XFILL_4_DFFPOSX1_298 gnd vdd FILL
XFILL_2_CLKBUF1_91 gnd vdd FILL
XFILL_2_CLKBUF1_80 gnd vdd FILL
XFILL_29_16_1 gnd vdd FILL
XFILL_1_BUFX2_133 gnd vdd FILL
XFILL_1_BUFX2_122 gnd vdd FILL
XFILL_1_BUFX2_166 gnd vdd FILL
XFILL_1_BUFX2_177 gnd vdd FILL
XFILL_0_BUFX2_915 gnd vdd FILL
XOAI21X1_172 BUFX4_10/Y BUFX4_385/Y BUFX2_951/A gnd OAI21X1_173/C vdd OAI21X1
XOAI21X1_161 BUFX4_148/Y INVX2_190/Y OAI21X1_161/C gnd OAI21X1_161/Y vdd OAI21X1
XFILL_0_BUFX2_904 gnd vdd FILL
XFILL_23_12_0 gnd vdd FILL
XFILL_1_BUFX2_188 gnd vdd FILL
XOAI21X1_150 BUFX4_1/A BUFX4_330/Y BUFX2_938/A gnd OAI21X1_151/C vdd OAI21X1
XOAI21X1_183 BUFX4_134/Y INVX2_201/Y OAI21X1_183/C gnd OAI21X1_183/Y vdd OAI21X1
XFILL_0_BUFX2_937 gnd vdd FILL
XFILL_0_BUFX2_948 gnd vdd FILL
XOAI21X1_194 BUFX4_106/Y BUFX4_311/Y BUFX2_963/A gnd OAI21X1_195/C vdd OAI21X1
XINVX1_225 INVX1_225/A gnd INVX1_225/Y vdd INVX1
XINVX1_203 OR2X2_17/Y gnd INVX1_203/Y vdd INVX1
XINVX1_214 INVX1_214/A gnd INVX1_214/Y vdd INVX1
XFILL_0_BUFX2_926 gnd vdd FILL
XFILL_0_BUFX2_959 gnd vdd FILL
XFILL_6_DFFPOSX1_304 gnd vdd FILL
XFILL_6_DFFPOSX1_315 gnd vdd FILL
XNAND2X1_25 BUFX2_850/A BUFX4_216/Y gnd OAI21X1_25/C vdd NAND2X1
XNAND2X1_14 BUFX2_897/A BUFX4_219/Y gnd OAI21X1_14/C vdd NAND2X1
XNAND2X1_58 BUFX2_887/A BUFX4_218/Y gnd OAI21X1_58/C vdd NAND2X1
XFILL_0_XNOR2X1_21 gnd vdd FILL
XFILL_2_INVX8_4 gnd vdd FILL
XNAND2X1_47 BUFX2_874/A BUFX4_188/Y gnd OAI21X1_47/C vdd NAND2X1
XFILL_0_XNOR2X1_10 gnd vdd FILL
XNAND2X1_36 BUFX2_862/A BUFX4_196/Y gnd OAI21X1_36/C vdd NAND2X1
XNAND2X1_69 BUFX2_899/A BUFX4_230/Y gnd OAI21X1_69/C vdd NAND2X1
XFILL_0_XNOR2X1_32 gnd vdd FILL
XFILL_0_XNOR2X1_43 gnd vdd FILL
XFILL_0_XNOR2X1_54 gnd vdd FILL
XFILL_4_17_1 gnd vdd FILL
XFILL_0_XNOR2X1_76 gnd vdd FILL
XFILL_0_XNOR2X1_65 gnd vdd FILL
XFILL_0_XNOR2X1_87 gnd vdd FILL
XFILL_0_XNOR2X1_98 gnd vdd FILL
XFILL_32_1_1 gnd vdd FILL
XFILL_28_11_0 gnd vdd FILL
XOAI21X1_1413 INVX4_50/Y INVX2_94/Y INVX2_63/Y gnd NAND2X1_625/A vdd OAI21X1
XOAI21X1_1402 INVX4_50/Y INVX2_59/Y INVX2_60/Y gnd OAI21X1_1403/C vdd OAI21X1
XFILL_0_BUFX4_230 gnd vdd FILL
XFILL_0_BUFX4_241 gnd vdd FILL
XFILL_1_OAI21X1_1600 gnd vdd FILL
XFILL_1_OAI21X1_1622 gnd vdd FILL
XOAI21X1_1424 OAI21X1_1424/A BUFX4_289/Y OAI21X1_1424/C gnd OAI21X1_1424/Y vdd OAI21X1
XOAI21X1_1435 XNOR2X1_93/Y BUFX4_291/Y OAI21X1_1435/C gnd OAI21X1_1435/Y vdd OAI21X1
XOAI21X1_1457 XNOR2X1_97/Y BUFX4_292/Y OAI21X1_1457/C gnd OAI21X1_1457/Y vdd OAI21X1
XFILL_0_BUFX4_263 gnd vdd FILL
XFILL_0_BUFX4_252 gnd vdd FILL
XFILL_0_BUFX4_274 gnd vdd FILL
XFILL_0_BUFX4_285 gnd vdd FILL
XNOR3X1_2 NOR3X1_2/A NOR3X1_2/B NOR3X1_2/C gnd NOR3X1_2/Y vdd NOR3X1
XOAI21X1_1446 BUFX4_169/Y BUFX4_80/A BUFX2_207/A gnd OAI21X1_1447/C vdd OAI21X1
XFILL_1_OAI21X1_1633 gnd vdd FILL
XFILL_1_OAI21X1_1611 gnd vdd FILL
XFILL_1_OAI21X1_1666 gnd vdd FILL
XOAI21X1_1479 OAI21X1_1479/A BUFX4_301/Y OAI21X1_1479/C gnd OAI21X1_1479/Y vdd OAI21X1
XFILL_0_BUFX4_296 gnd vdd FILL
XOAI21X1_1468 NOR2X1_145/A INVX2_109/Y OAI21X1_1468/C gnd OAI21X1_1470/A vdd OAI21X1
XFILL_1_OAI21X1_1655 gnd vdd FILL
XFILL_1_OAI21X1_1644 gnd vdd FILL
XFILL_0_OAI21X1_413 gnd vdd FILL
XFILL_0_OAI21X1_402 gnd vdd FILL
XFILL_1_OAI21X1_1688 gnd vdd FILL
XFILL_1_OAI21X1_1677 gnd vdd FILL
XFILL_1_OAI21X1_1699 gnd vdd FILL
XFILL_1_OAI21X1_606 gnd vdd FILL
XFILL_0_OAI21X1_446 gnd vdd FILL
XFILL_1_OAI21X1_617 gnd vdd FILL
XFILL_0_OAI21X1_424 gnd vdd FILL
XFILL_0_OAI21X1_435 gnd vdd FILL
XFILL_1_OAI21X1_628 gnd vdd FILL
XFILL_0_OAI21X1_457 gnd vdd FILL
XFILL_1_OAI21X1_639 gnd vdd FILL
XFILL_0_OAI21X1_479 gnd vdd FILL
XFILL_9_16_1 gnd vdd FILL
XFILL_0_OAI21X1_468 gnd vdd FILL
XFILL_3_DFFPOSX1_1032 gnd vdd FILL
XFILL_3_DFFPOSX1_1021 gnd vdd FILL
XFILL_6_DFFPOSX1_882 gnd vdd FILL
XFILL_6_DFFPOSX1_871 gnd vdd FILL
XFILL_3_DFFPOSX1_1010 gnd vdd FILL
XFILL_6_DFFPOSX1_893 gnd vdd FILL
XFILL_1_XNOR2X1_1 gnd vdd FILL
XFILL_3_12_0 gnd vdd FILL
XFILL_0_OAI21X1_1212 gnd vdd FILL
XFILL_0_OAI21X1_1223 gnd vdd FILL
XFILL_0_NAND2X1_430 gnd vdd FILL
XFILL_1_NAND2X1_623 gnd vdd FILL
XFILL_0_OAI21X1_1201 gnd vdd FILL
XFILL_1_NAND2X1_612 gnd vdd FILL
XFILL_0_NAND2X1_441 gnd vdd FILL
XFILL_0_NAND2X1_452 gnd vdd FILL
XFILL_0_NAND2X1_474 gnd vdd FILL
XFILL_0_DFFPOSX1_813 gnd vdd FILL
XFILL_0_OAI21X1_1256 gnd vdd FILL
XFILL_0_NAND2X1_485 gnd vdd FILL
XFILL_0_OAI21X1_1234 gnd vdd FILL
XFILL_0_DFFPOSX1_824 gnd vdd FILL
XFILL_0_NAND2X1_496 gnd vdd FILL
XFILL_0_OAI21X1_1245 gnd vdd FILL
XFILL_1_NAND2X1_634 gnd vdd FILL
XFILL_0_DFFPOSX1_802 gnd vdd FILL
XFILL_1_NAND2X1_645 gnd vdd FILL
XFILL_0_NAND2X1_463 gnd vdd FILL
XFILL_1_NAND2X1_656 gnd vdd FILL
XFILL_1_NAND2X1_689 gnd vdd FILL
XFILL_1_NAND2X1_678 gnd vdd FILL
XFILL_0_DFFPOSX1_835 gnd vdd FILL
XFILL_23_1_1 gnd vdd FILL
XFILL_0_OAI21X1_1289 gnd vdd FILL
XFILL_0_DFFPOSX1_868 gnd vdd FILL
XFILL_0_OAI21X1_1278 gnd vdd FILL
XFILL_0_DFFPOSX1_857 gnd vdd FILL
XFILL_0_OAI21X1_1267 gnd vdd FILL
XFILL_0_DFFPOSX1_846 gnd vdd FILL
XFILL_0_DFFPOSX1_879 gnd vdd FILL
XDFFPOSX1_1009 BUFX2_676/A CLKBUF1_58/Y OAI21X1_1586/Y gnd vdd DFFPOSX1
XFILL_5_DFFPOSX1_450 gnd vdd FILL
XFILL_5_DFFPOSX1_461 gnd vdd FILL
XFILL_5_DFFPOSX1_472 gnd vdd FILL
XFILL_5_DFFPOSX1_483 gnd vdd FILL
XFILL_5_DFFPOSX1_494 gnd vdd FILL
XFILL_0_AOI21X1_21 gnd vdd FILL
XFILL_0_AOI21X1_10 gnd vdd FILL
XFILL_0_AOI21X1_32 gnd vdd FILL
XFILL_2_CLKBUF1_1 gnd vdd FILL
XFILL_0_AOI21X1_54 gnd vdd FILL
XFILL_0_AOI21X1_65 gnd vdd FILL
XFILL_0_AOI21X1_43 gnd vdd FILL
XFILL_0_OAI21X1_991 gnd vdd FILL
XFILL_0_OAI21X1_980 gnd vdd FILL
XFILL_8_11_0 gnd vdd FILL
XFILL_6_2_1 gnd vdd FILL
XFILL_2_DFFPOSX1_918 gnd vdd FILL
XFILL_2_DFFPOSX1_929 gnd vdd FILL
XFILL_2_DFFPOSX1_907 gnd vdd FILL
XFILL_2_BUFX4_150 gnd vdd FILL
XFILL_6_DFFPOSX1_1014 gnd vdd FILL
XFILL_6_DFFPOSX1_1025 gnd vdd FILL
XFILL_2_BUFX4_183 gnd vdd FILL
XFILL_14_1_1 gnd vdd FILL
XFILL_0_OAI21X1_1790 gnd vdd FILL
XFILL_0_BUFX2_712 gnd vdd FILL
XFILL_0_BUFX2_723 gnd vdd FILL
XFILL_0_NOR2X1_41 gnd vdd FILL
XFILL_0_NOR2X1_30 gnd vdd FILL
XFILL_0_BUFX2_701 gnd vdd FILL
XFILL_0_BUFX2_745 gnd vdd FILL
XFILL_0_BUFX2_734 gnd vdd FILL
XFILL_0_BUFX2_756 gnd vdd FILL
XFILL_0_NOR2X1_52 gnd vdd FILL
XFILL_0_BUFX2_767 gnd vdd FILL
XFILL_0_NOR2X1_85 gnd vdd FILL
XFILL_0_NOR2X1_74 gnd vdd FILL
XFILL_0_NOR2X1_63 gnd vdd FILL
XFILL_1_DFFPOSX1_519 gnd vdd FILL
XFILL_1_DFFPOSX1_508 gnd vdd FILL
XFILL_0_NOR2X1_96 gnd vdd FILL
XFILL_0_BUFX2_778 gnd vdd FILL
XFILL_0_BUFX2_789 gnd vdd FILL
XFILL_6_DFFPOSX1_156 gnd vdd FILL
XFILL_3_DFFPOSX1_7 gnd vdd FILL
XFILL_6_DFFPOSX1_167 gnd vdd FILL
XFILL_6_DFFPOSX1_178 gnd vdd FILL
XFILL_6_DFFPOSX1_189 gnd vdd FILL
XFILL_14_17_0 gnd vdd FILL
XBUFX4_331 BUFX4_384/A gnd NAND2X1_7/B vdd BUFX4
XBUFX4_320 BUFX4_388/A gnd BUFX4_320/Y vdd BUFX4
XBUFX4_353 BUFX4_386/A gnd BUFX4_353/Y vdd BUFX4
XFILL_30_10_1 gnd vdd FILL
XBUFX4_342 BUFX4_381/A gnd BUFX4_342/Y vdd BUFX4
XBUFX4_364 BUFX4_384/A gnd BUFX4_364/Y vdd BUFX4
XBUFX4_386 BUFX4_386/A gnd BUFX4_386/Y vdd BUFX4
XBUFX4_375 BUFX4_381/A gnd BUFX4_375/Y vdd BUFX4
XFILL_34_9_0 gnd vdd FILL
XFILL_0_DFFPOSX1_109 gnd vdd FILL
XFILL_26_1 gnd vdd FILL
XOAI21X1_908 BUFX4_112/Y BUFX4_382/Y BUFX2_325/A gnd OAI21X1_909/C vdd OAI21X1
XFILL_0_NAND2X1_7 gnd vdd FILL
XOAI21X1_919 BUFX4_139/Y INVX1_114/Y OAI21X1_919/C gnd OAI21X1_919/Y vdd OAI21X1
XOAI21X1_1221 INVX1_183/A INVX2_58/Y INVX2_59/Y gnd OAI21X1_1222/C vdd OAI21X1
XOAI21X1_1210 BUFX4_98/Y BUFX4_366/Y BUFX2_130/A gnd OAI21X1_1211/C vdd OAI21X1
XOAI21X1_1232 BUFX4_251/Y BUFX4_312/Y BUFX2_192/A gnd OAI21X1_1233/C vdd OAI21X1
XDFFPOSX1_822 BUFX2_71/A CLKBUF1_70/Y OAI21X1_1128/Y gnd vdd DFFPOSX1
XOAI21X1_1254 BUFX4_97/Y BUFX4_359/Y BUFX2_137/A gnd OAI21X1_1255/C vdd OAI21X1
XFILL_1_OAI21X1_1430 gnd vdd FILL
XOAI21X1_1243 NOR2X1_183/A INVX1_201/A OAI21X1_1243/C gnd OAI21X1_1245/A vdd OAI21X1
XDFFPOSX1_811 BUFX2_88/A CLKBUF1_7/Y OAI21X1_1103/Y gnd vdd DFFPOSX1
XDFFPOSX1_833 BUFX2_83/A CLKBUF1_16/Y OAI21X1_1144/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1441 gnd vdd FILL
XOAI21X1_1265 OR2X2_18/A NOR3X1_18/C OAI21X1_1265/C gnd OAI21X1_1267/A vdd OAI21X1
XDFFPOSX1_800 BUFX2_53/A CLKBUF1_71/Y OAI21X1_1092/Y gnd vdd DFFPOSX1
XDFFPOSX1_855 BUFX2_107/A CLKBUF1_21/Y OAI21X1_1176/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1474 gnd vdd FILL
XFILL_1_OAI21X1_1463 gnd vdd FILL
XOAI21X1_1287 AOI21X1_47/Y OAI21X1_1287/B OAI21X1_1287/C gnd OAI21X1_1287/Y vdd OAI21X1
XOAI21X1_1298 AND2X2_30/A INVX2_75/Y MUX2X1_2/S gnd OAI21X1_1299/B vdd OAI21X1
XDFFPOSX1_866 BUFX2_119/A CLKBUF1_36/Y OAI21X1_1197/Y gnd vdd DFFPOSX1
XOAI21X1_1276 BUFX4_4/A OAI21X1_5/A BUFX2_146/A gnd OAI21X1_1277/C vdd OAI21X1
XFILL_0_OAI21X1_221 gnd vdd FILL
XFILL_1_OAI21X1_1452 gnd vdd FILL
XDFFPOSX1_844 BUFX2_95/A CLKBUF1_62/Y OAI21X1_1160/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_210 gnd vdd FILL
XFILL_0_OAI21X1_254 gnd vdd FILL
XDFFPOSX1_888 BUFX2_137/A CLKBUF1_23/Y OAI21X1_1255/Y gnd vdd DFFPOSX1
XDFFPOSX1_877 BUFX2_174/A CLKBUF1_31/Y OAI21X1_1220/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_232 gnd vdd FILL
XFILL_0_OAI21X1_243 gnd vdd FILL
XDFFPOSX1_899 BUFX2_149/A CLKBUF1_49/Y OAI21X1_1284/Y gnd vdd DFFPOSX1
XINVX2_27 bundleStartMajId_i[25] gnd NOR3X1_6/A vdd INVX2
XFILL_1_OAI21X1_1496 gnd vdd FILL
XFILL_1_OAI21X1_1485 gnd vdd FILL
XFILL_1_OAI21X1_414 gnd vdd FILL
XINVX2_16 bundleStartMajId_i[49] gnd NOR2X1_9/A vdd INVX2
XFILL_1_OAI21X1_403 gnd vdd FILL
XFILL_1_OAI21X1_436 gnd vdd FILL
XFILL_1_OAI21X1_425 gnd vdd FILL
XFILL_0_OAI21X1_276 gnd vdd FILL
XFILL_0_OAI21X1_298 gnd vdd FILL
XFILL_0_OAI21X1_287 gnd vdd FILL
XINVX2_38 bundleStartMajId_i[3] gnd INVX2_38/Y vdd INVX2
XFILL_19_16_0 gnd vdd FILL
XFILL_1_OAI21X1_458 gnd vdd FILL
XINVX2_49 INVX2_49/A gnd INVX2_49/Y vdd INVX2
XFILL_1_OAI21X1_447 gnd vdd FILL
XFILL_1_OAI21X1_469 gnd vdd FILL
XFILL_0_OAI21X1_265 gnd vdd FILL
XFILL_32_18_0 gnd vdd FILL
XFILL_0_OAI21X1_1031 gnd vdd FILL
XFILL_0_OAI21X1_1020 gnd vdd FILL
XFILL_1_INVX4_38 gnd vdd FILL
XFILL_25_9_0 gnd vdd FILL
XFILL_1_NAND2X1_420 gnd vdd FILL
XFILL_0_NAND2X1_260 gnd vdd FILL
XFILL_1_INVX4_49 gnd vdd FILL
XFILL_0_9_0 gnd vdd FILL
XFILL_1_NAND2X1_442 gnd vdd FILL
XFILL_0_OAI21X1_1053 gnd vdd FILL
XFILL_0_OAI21X1_1042 gnd vdd FILL
XFILL_0_DFFPOSX1_632 gnd vdd FILL
XFILL_0_OAI21X1_1064 gnd vdd FILL
XFILL_0_DFFPOSX1_621 gnd vdd FILL
XFILL_0_DFFPOSX1_610 gnd vdd FILL
XFILL_0_NAND2X1_282 gnd vdd FILL
XFILL_0_NAND2X1_293 gnd vdd FILL
XFILL_0_DFFPOSX1_643 gnd vdd FILL
XFILL_1_BUFX4_206 gnd vdd FILL
XFILL_0_OAI21X1_1075 gnd vdd FILL
XFILL_1_BUFX4_228 gnd vdd FILL
XFILL_0_NAND2X1_271 gnd vdd FILL
XFILL_1_NAND2X1_453 gnd vdd FILL
XFILL_1_BUFX4_217 gnd vdd FILL
XFILL_0_DFFPOSX1_654 gnd vdd FILL
XFILL_1_NAND2X1_486 gnd vdd FILL
XFILL_1_BUFX4_239 gnd vdd FILL
XFILL_0_OAI21X1_1097 gnd vdd FILL
XFILL_0_DFFPOSX1_665 gnd vdd FILL
XFILL_0_DFFPOSX1_676 gnd vdd FILL
XFILL_0_OAI21X1_1086 gnd vdd FILL
XFILL_0_DFFPOSX1_698 gnd vdd FILL
XFILL_0_DFFPOSX1_687 gnd vdd FILL
XFILL_5_DFFPOSX1_280 gnd vdd FILL
XFILL_5_DFFPOSX1_291 gnd vdd FILL
XFILL_37_17_0 gnd vdd FILL
XFILL_2_BUFX4_33 gnd vdd FILL
XFILL_1_OAI21X1_970 gnd vdd FILL
XFILL_1_OAI21X1_981 gnd vdd FILL
XFILL_2_BUFX4_66 gnd vdd FILL
XFILL_1_OAI21X1_992 gnd vdd FILL
XFILL_2_DFFPOSX1_704 gnd vdd FILL
XBUFX2_802 BUFX2_802/A gnd tid1_o[32] vdd BUFX2
XBUFX2_813 BUFX2_813/A gnd tid1_o[22] vdd BUFX2
XFILL_2_DFFPOSX1_715 gnd vdd FILL
XFILL_2_DFFPOSX1_737 gnd vdd FILL
XFILL_2_DFFPOSX1_748 gnd vdd FILL
XBUFX2_824 BUFX2_824/A gnd tid1_o[12] vdd BUFX2
XFILL_2_DFFPOSX1_726 gnd vdd FILL
XBUFX2_846 BUFX2_846/A gnd tid2_o[50] vdd BUFX2
XBUFX2_835 NAND2X1_5/A gnd tid1_o[2] vdd BUFX2
XBUFX2_868 BUFX2_868/A gnd tid2_o[30] vdd BUFX2
XFILL_2_DFFPOSX1_759 gnd vdd FILL
XBUFX2_879 BUFX2_879/A gnd tid2_o[20] vdd BUFX2
XBUFX2_857 BUFX2_857/A gnd tid2_o[40] vdd BUFX2
XFILL_16_9_0 gnd vdd FILL
XFILL_2_NAND3X1_60 gnd vdd FILL
XFILL_0_NOR2X1_219 gnd vdd FILL
XFILL_0_NOR2X1_208 gnd vdd FILL
XDFFPOSX1_118 BUFX2_787/A CLKBUF1_89/Y OAI21X1_1792/Y gnd vdd DFFPOSX1
XDFFPOSX1_107 BUFX2_838/A CLKBUF1_26/Y OAI21X1_1781/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_542 gnd vdd FILL
XFILL_0_BUFX2_520 gnd vdd FILL
XFILL_1_DFFPOSX1_305 gnd vdd FILL
XFILL_0_BUFX2_531 gnd vdd FILL
XFILL_1_DFFPOSX1_316 gnd vdd FILL
XFILL_0_BUFX2_575 gnd vdd FILL
XCLKBUF1_1 BUFX4_91/Y gnd CLKBUF1_1/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_327 gnd vdd FILL
XFILL_1_DFFPOSX1_338 gnd vdd FILL
XDFFPOSX1_129 BUFX2_799/A CLKBUF1_62/Y OAI21X1_1803/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_553 gnd vdd FILL
XFILL_0_BUFX2_564 gnd vdd FILL
XFILL_1_DFFPOSX1_349 gnd vdd FILL
XFILL_0_BUFX2_597 gnd vdd FILL
XFILL_0_BUFX2_586 gnd vdd FILL
XFILL_4_DFFPOSX1_809 gnd vdd FILL
XFILL_37_0_1 gnd vdd FILL
XFILL_4_CLKBUF1_32 gnd vdd FILL
XBUFX4_172 BUFX4_14/Y gnd BUFX4_172/Y vdd BUFX4
XBUFX4_150 BUFX4_17/Y gnd BUFX4_150/Y vdd BUFX4
XFILL_0_INVX1_61 gnd vdd FILL
XFILL_4_CLKBUF1_21 gnd vdd FILL
XBUFX4_161 BUFX4_17/Y gnd BUFX4_161/Y vdd BUFX4
XFILL_0_INVX1_50 gnd vdd FILL
XFILL_2_OAI21X1_1692 gnd vdd FILL
XFILL_4_CLKBUF1_65 gnd vdd FILL
XBUFX4_183 BUFX4_24/Y gnd BUFX4_183/Y vdd BUFX4
XNOR2X1_232 bundleAddress_i[4] INVX2_112/Y gnd NOR2X1_232/Y vdd NOR2X1
XNOR2X1_221 INVX2_97/Y INVX4_51/Y gnd NOR2X1_221/Y vdd NOR2X1
XNOR2X1_210 INVX1_197/A NOR2X1_210/B gnd INVX1_216/A vdd NOR2X1
XFILL_0_INVX1_83 gnd vdd FILL
XFILL_0_INVX1_72 gnd vdd FILL
XFILL_0_INVX1_94 gnd vdd FILL
XFILL_4_CLKBUF1_54 gnd vdd FILL
XBUFX4_194 BUFX4_22/Y gnd BUFX4_194/Y vdd BUFX4
XFILL_4_CLKBUF1_76 gnd vdd FILL
XFILL_0_BUFX2_25 gnd vdd FILL
XFILL_4_CLKBUF1_98 gnd vdd FILL
XFILL_4_CLKBUF1_87 gnd vdd FILL
XFILL_0_BUFX2_36 gnd vdd FILL
XFILL_0_BUFX2_14 gnd vdd FILL
XFILL_0_BUFX2_69 gnd vdd FILL
XFILL_0_BUFX2_58 gnd vdd FILL
XFILL_1_NOR2X1_28 gnd vdd FILL
XFILL_0_BUFX2_47 gnd vdd FILL
XFILL_1_NOR2X1_39 gnd vdd FILL
XOAI21X1_705 BUFX4_131/Y BUFX4_61/Y BUFX2_593/A gnd OAI21X1_706/C vdd OAI21X1
XOAI21X1_738 XNOR2X1_46/Y BUFX4_295/Y OAI21X1_738/C gnd OAI21X1_738/Y vdd OAI21X1
XOAI21X1_749 BUFX4_155/Y BUFX4_61/Y BUFX2_611/A gnd OAI21X1_750/C vdd OAI21X1
XOAI21X1_716 NOR2X1_106/Y bundleStartMajId_i[43] BUFX4_287/Y gnd OAI21X1_718/B vdd
+ OAI21X1
XOAI21X1_727 NOR3X1_9/A NOR2X1_30/A INVX4_10/Y gnd OAI21X1_727/Y vdd OAI21X1
XOAI21X1_1040 BUFX4_347/Y INVX2_57/Y NAND2X1_406/Y gnd OAI21X1_1040/Y vdd OAI21X1
XFILL_21_15_1 gnd vdd FILL
XOAI21X1_1051 BUFX4_385/Y INVX2_67/Y NAND2X1_417/Y gnd OAI21X1_1051/Y vdd OAI21X1
XDFFPOSX1_630 INVX1_59/A CLKBUF1_61/Y OAI21X1_858/Y gnd vdd DFFPOSX1
XOAI21X1_1062 BUFX4_317/Y INVX2_71/Y NAND2X1_428/Y gnd OAI21X1_1062/Y vdd OAI21X1
XOAI21X1_1073 BUFX4_370/Y INVX4_41/Y NAND2X1_439/Y gnd OAI21X1_1073/Y vdd OAI21X1
XDFFPOSX1_641 INVX1_70/A CLKBUF1_82/Y OAI21X1_869/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1260 gnd vdd FILL
XFILL_1_OAI21X1_200 gnd vdd FILL
XFILL_1_OAI21X1_1293 gnd vdd FILL
XFILL_1_OAI21X1_1282 gnd vdd FILL
XOAI21X1_1084 BUFX4_375/Y INVX1_179/Y NAND2X1_450/Y gnd OAI21X1_1084/Y vdd OAI21X1
XOAI21X1_1095 BUFX4_360/Y INVX2_90/Y NAND2X1_461/Y gnd OAI21X1_1095/Y vdd OAI21X1
XFILL_1_DFFPOSX1_850 gnd vdd FILL
XFILL_1_OAI21X1_1271 gnd vdd FILL
XDFFPOSX1_652 BUFX2_319/A CLKBUF1_41/Y OAI21X1_880/Y gnd vdd DFFPOSX1
XDFFPOSX1_663 BUFX2_300/A CLKBUF1_82/Y OAI21X1_891/Y gnd vdd DFFPOSX1
XDFFPOSX1_674 BUFX2_312/A CLKBUF1_54/Y OAI21X1_902/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_861 gnd vdd FILL
XFILL_1_DFFPOSX1_883 gnd vdd FILL
XFILL_1_DFFPOSX1_872 gnd vdd FILL
XFILL_1_OAI21X1_222 gnd vdd FILL
XFILL_1_OAI21X1_233 gnd vdd FILL
XNAND2X1_700 BUFX2_691/A BUFX4_230/Y gnd NAND2X1_700/Y vdd NAND2X1
XFILL_1_OAI21X1_244 gnd vdd FILL
XFILL_1_DFFPOSX1_894 gnd vdd FILL
XDFFPOSX1_696 BUFX2_333/A CLKBUF1_40/Y OAI21X1_941/Y gnd vdd DFFPOSX1
XNAND2X1_711 BUFX2_703/A BUFX4_188/Y gnd NAND2X1_711/Y vdd NAND2X1
XFILL_1_OAI21X1_211 gnd vdd FILL
XDFFPOSX1_685 BUFX2_352/A CLKBUF1_58/Y OAI21X1_919/Y gnd vdd DFFPOSX1
XFILL_0_NOR2X1_5 gnd vdd FILL
XFILL_1_OAI21X1_255 gnd vdd FILL
XFILL_1_OAI21X1_277 gnd vdd FILL
XNAND2X1_733 BUFX2_787/A BUFX4_318/Y gnd NAND2X1_733/Y vdd NAND2X1
XFILL_1_OAI21X1_266 gnd vdd FILL
XNAND2X1_722 BUFX2_838/A BUFX4_348/Y gnd NAND2X1_722/Y vdd NAND2X1
XNAND2X1_744 BUFX2_799/A BUFX4_384/Y gnd NAND2X1_744/Y vdd NAND2X1
XNAND2X1_755 BUFX2_812/A BUFX4_354/Y gnd NAND2X1_755/Y vdd NAND2X1
XFILL_1_OAI21X1_299 gnd vdd FILL
XFILL_1_OAI21X1_288 gnd vdd FILL
XNAND2X1_766 BUFX2_824/A BUFX4_348/Y gnd NAND2X1_766/Y vdd NAND2X1
XFILL_2_XNOR2X1_17 gnd vdd FILL
XFILL_2_XNOR2X1_28 gnd vdd FILL
XFILL_28_0_1 gnd vdd FILL
XFILL_2_XNOR2X1_39 gnd vdd FILL
XBUFX2_109 BUFX2_109/A gnd addr2_o[14] vdd BUFX2
XFILL_3_0_1 gnd vdd FILL
XFILL_1_NAND2X1_250 gnd vdd FILL
XFILL_1_NAND2X1_261 gnd vdd FILL
XFILL_0_DFFPOSX1_451 gnd vdd FILL
XFILL_1_NAND2X1_283 gnd vdd FILL
XFILL_0_DFFPOSX1_440 gnd vdd FILL
XFILL_1_NAND2X1_272 gnd vdd FILL
XFILL_2_DFFPOSX1_4 gnd vdd FILL
XFILL_26_14_1 gnd vdd FILL
XFILL_0_DFFPOSX1_484 gnd vdd FILL
XFILL_0_DFFPOSX1_462 gnd vdd FILL
XFILL_1_NAND2X1_294 gnd vdd FILL
XFILL_0_DFFPOSX1_473 gnd vdd FILL
XINVX8_3 bundleAddress_i[24] gnd INVX8_3/Y vdd INVX8
XFILL_0_DFFPOSX1_495 gnd vdd FILL
XFILL_3_DFFPOSX1_900 gnd vdd FILL
XFILL_3_DFFPOSX1_922 gnd vdd FILL
XFILL_3_DFFPOSX1_911 gnd vdd FILL
XFILL_3_DFFPOSX1_944 gnd vdd FILL
XFILL_3_DFFPOSX1_966 gnd vdd FILL
XFILL_3_DFFPOSX1_955 gnd vdd FILL
XFILL_3_DFFPOSX1_933 gnd vdd FILL
XFILL_3_DFFPOSX1_999 gnd vdd FILL
XFILL_20_10_0 gnd vdd FILL
XFILL_3_DFFPOSX1_977 gnd vdd FILL
XFILL_3_DFFPOSX1_988 gnd vdd FILL
XBUFX4_34 BUFX4_60/A gnd BUFX4_34/Y vdd BUFX4
XBUFX4_23 BUFX4_26/A gnd BUFX4_23/Y vdd BUFX4
XBUFX4_12 BUFX4_1/A gnd BUFX4_12/Y vdd BUFX4
XBUFX4_67 BUFX4_67/A gnd BUFX4_67/Y vdd BUFX4
XBUFX4_45 BUFX4_51/A gnd BUFX4_45/Y vdd BUFX4
XBUFX4_56 BUFX4_71/A gnd BUFX4_56/Y vdd BUFX4
XBUFX4_78 BUFX4_80/A gnd BUFX4_78/Y vdd BUFX4
XFILL_19_0_1 gnd vdd FILL
XFILL_2_DFFPOSX1_512 gnd vdd FILL
XBUFX4_89 clock_i gnd BUFX4_89/Y vdd BUFX4
XBUFX2_621 BUFX2_621/A gnd majID4_o[22] vdd BUFX2
XFILL_2_DFFPOSX1_501 gnd vdd FILL
XFILL_2_DFFPOSX1_523 gnd vdd FILL
XBUFX2_610 INVX1_39/A gnd majID4_o[32] vdd BUFX2
XBUFX2_654 BUFX2_654/A gnd pid1_o[18] vdd BUFX2
XFILL_2_DFFPOSX1_545 gnd vdd FILL
XBUFX2_643 BUFX2_643/A gnd majID4_o[2] vdd BUFX2
XBUFX2_632 BUFX2_632/A gnd majID4_o[12] vdd BUFX2
XFILL_2_DFFPOSX1_534 gnd vdd FILL
XFILL_1_15_1 gnd vdd FILL
XFILL_2_DFFPOSX1_556 gnd vdd FILL
XBUFX2_665 BUFX2_665/A gnd pid1_o[8] vdd BUFX2
XBUFX2_687 BUFX2_687/A gnd pid2_o[17] vdd BUFX2
XFILL_2_DFFPOSX1_578 gnd vdd FILL
XFILL_2_DFFPOSX1_567 gnd vdd FILL
XFILL_2_DFFPOSX1_589 gnd vdd FILL
XBUFX2_676 BUFX2_676/A gnd pid1_o[26] vdd BUFX2
XBUFX2_698 BUFX2_698/A gnd pid2_o[7] vdd BUFX2
XFILL_31_7_0 gnd vdd FILL
XOR2X2_15 OR2X2_15/A OR2X2_15/B gnd OR2X2_15/Y vdd OR2X2
XINVX2_150 bundleTid_i[59] gnd INVX2_150/Y vdd INVX2
XFILL_0_BUFX2_350 gnd vdd FILL
XFILL_1_DFFPOSX1_102 gnd vdd FILL
XFILL_1_DFFPOSX1_113 gnd vdd FILL
XINVX2_172 bundleTid_i[37] gnd INVX2_172/Y vdd INVX2
XINVX2_161 bundleTid_i[48] gnd INVX2_161/Y vdd INVX2
XFILL_1_DFFPOSX1_124 gnd vdd FILL
XINVX2_183 bundleTid_i[26] gnd INVX2_183/Y vdd INVX2
XFILL_0_BUFX2_383 gnd vdd FILL
XFILL_1_DFFPOSX1_135 gnd vdd FILL
XOR2X2_8 OR2X2_8/A OR2X2_8/B gnd OR2X2_9/B vdd OR2X2
XFILL_1_DFFPOSX1_146 gnd vdd FILL
XFILL_0_BUFX2_372 gnd vdd FILL
XFILL_0_BUFX2_361 gnd vdd FILL
XINVX2_194 bundleTid_i[15] gnd INVX2_194/Y vdd INVX2
XFILL_1_DFFPOSX1_157 gnd vdd FILL
XFILL_1_DFFPOSX1_179 gnd vdd FILL
XFILL_1_DFFPOSX1_168 gnd vdd FILL
XFILL_0_BUFX2_394 gnd vdd FILL
XFILL_4_DFFPOSX1_606 gnd vdd FILL
XFILL_4_DFFPOSX1_617 gnd vdd FILL
XFILL_4_DFFPOSX1_628 gnd vdd FILL
XFILL_4_DFFPOSX1_639 gnd vdd FILL
XFILL_6_14_1 gnd vdd FILL
XFILL_0_10_0 gnd vdd FILL
XFILL_22_7_0 gnd vdd FILL
XFILL_1_BUFX2_518 gnd vdd FILL
XFILL_1_BUFX2_507 gnd vdd FILL
XOAI21X1_502 BUFX4_9/Y BUFX4_365/Y BUFX2_522/A gnd OAI21X1_503/C vdd OAI21X1
XOAI21X1_513 NOR2X1_59/Y bundleStartMajId_i[58] NOR2X1_89/B gnd OAI21X1_515/B vdd
+ OAI21X1
XFILL_3_DFFPOSX1_218 gnd vdd FILL
XFILL_3_DFFPOSX1_207 gnd vdd FILL
XOAI21X1_557 OR2X2_10/B OR2X2_2/Y INVX8_6/A gnd NOR2X1_65/B vdd OAI21X1
XOAI21X1_535 BUFX4_107/Y BUFX4_345/Y BUFX2_525/A gnd OAI21X1_536/C vdd OAI21X1
XOAI21X1_546 OAI21X1_546/A BUFX4_122/Y OAI21X1_546/C gnd OAI21X1_546/Y vdd OAI21X1
XOAI21X1_524 OAI21X1_524/A BUFX4_167/Y OAI21X1_524/C gnd OAI21X1_524/Y vdd OAI21X1
XFILL_3_DFFPOSX1_229 gnd vdd FILL
XOAI21X1_568 BUFX4_10/A BUFX4_334/Y BUFX2_540/A gnd OAI21X1_571/C vdd OAI21X1
XOAI21X1_579 BUFX4_104/Y BUFX4_378/Y BUFX2_545/A gnd OAI21X1_581/C vdd OAI21X1
XDFFPOSX1_471 BUFX2_504/A CLKBUF1_91/Y OAI21X1_478/Y gnd vdd DFFPOSX1
XDFFPOSX1_482 BUFX2_516/A CLKBUF1_19/Y OAI21X1_498/Y gnd vdd DFFPOSX1
XDFFPOSX1_460 BUFX2_492/A CLKBUF1_84/Y OAI21X1_459/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1090 gnd vdd FILL
XFILL_1_DFFPOSX1_691 gnd vdd FILL
XFILL_1_DFFPOSX1_680 gnd vdd FILL
XFILL_2_OAI21X1_201 gnd vdd FILL
XNAND2X1_530 BUFX2_89/A BUFX4_202/Y gnd NAND2X1_530/Y vdd NAND2X1
XDFFPOSX1_493 BUFX2_584/A CLKBUF1_100/Y OAI21X1_526/Y gnd vdd DFFPOSX1
XNAND2X1_552 BUFX2_104/A BUFX4_203/Y gnd NAND2X1_552/Y vdd NAND2X1
XNAND2X1_563 bundleAddress_i[17] bundleAddress_i[14] gnd NOR2X1_165/B vdd NAND2X1
XNAND2X1_541 bundleAddress_i[29] bundleAddress_i[26] gnd NOR2X1_155/B vdd NAND2X1
XNAND2X1_596 bundleAddress_i[46] NOR2X1_184/Y gnd NAND2X1_597/B vdd NAND2X1
XNAND2X1_585 BUFX2_123/A BUFX4_187/Y gnd NAND2X1_585/Y vdd NAND2X1
XNAND2X1_574 bundleAddress_i[13] INVX2_103/A gnd INVX1_196/A vdd NAND2X1
XFILL_5_8_0 gnd vdd FILL
XFILL_0_AND2X2_31 gnd vdd FILL
XFILL_0_AND2X2_20 gnd vdd FILL
XFILL_1_DFFPOSX1_1009 gnd vdd FILL
XFILL_13_7_0 gnd vdd FILL
XFILL_0_DFFPOSX1_281 gnd vdd FILL
XFILL_0_DFFPOSX1_292 gnd vdd FILL
XFILL_0_DFFPOSX1_270 gnd vdd FILL
XFILL_3_DFFPOSX1_741 gnd vdd FILL
XOAI21X1_1809 BUFX4_376/Y INVX2_181/Y NAND2X1_750/Y gnd OAI21X1_1809/Y vdd OAI21X1
XFILL_3_DFFPOSX1_730 gnd vdd FILL
XFILL_3_DFFPOSX1_752 gnd vdd FILL
XFILL_3_DFFPOSX1_774 gnd vdd FILL
XFILL_3_DFFPOSX1_763 gnd vdd FILL
XFILL_3_CLKBUF1_40 gnd vdd FILL
XFILL_3_CLKBUF1_51 gnd vdd FILL
XFILL_0_OAI21X1_809 gnd vdd FILL
XFILL_3_CLKBUF1_73 gnd vdd FILL
XFILL_3_CLKBUF1_84 gnd vdd FILL
XFILL_3_DFFPOSX1_785 gnd vdd FILL
XFILL_3_CLKBUF1_62 gnd vdd FILL
XFILL_3_DFFPOSX1_796 gnd vdd FILL
XFILL_3_CLKBUF1_95 gnd vdd FILL
XFILL_1_NOR2X1_191 gnd vdd FILL
XFILL_2_DFFPOSX1_331 gnd vdd FILL
XFILL_11_15_0 gnd vdd FILL
XFILL_2_DFFPOSX1_320 gnd vdd FILL
XFILL_2_DFFPOSX1_342 gnd vdd FILL
XFILL_0_OAI21X1_1608 gnd vdd FILL
XBUFX2_440 BUFX2_440/A gnd majID1_o[12] vdd BUFX2
XFILL_2_DFFPOSX1_353 gnd vdd FILL
XFILL_2_DFFPOSX1_364 gnd vdd FILL
XBUFX2_451 BUFX2_451/A gnd majID1_o[2] vdd BUFX2
XBUFX2_462 BUFX2_462/A gnd majID2_o[50] vdd BUFX2
XFILL_0_OAI21X1_1619 gnd vdd FILL
XFILL_2_DFFPOSX1_375 gnd vdd FILL
XBUFX2_495 BUFX2_495/A gnd majID2_o[20] vdd BUFX2
XFILL_2_DFFPOSX1_397 gnd vdd FILL
XFILL_2_DFFPOSX1_386 gnd vdd FILL
XBUFX2_473 BUFX2_473/A gnd majID2_o[40] vdd BUFX2
XBUFX2_484 BUFX2_484/A gnd majID2_o[30] vdd BUFX2
XFILL_5_DFFPOSX1_813 gnd vdd FILL
XFILL_5_DFFPOSX1_802 gnd vdd FILL
XFILL_5_DFFPOSX1_835 gnd vdd FILL
XFILL_5_DFFPOSX1_824 gnd vdd FILL
XFILL_5_DFFPOSX1_846 gnd vdd FILL
XFILL_5_DFFPOSX1_879 gnd vdd FILL
XFILL_5_DFFPOSX1_868 gnd vdd FILL
XFILL_5_DFFPOSX1_857 gnd vdd FILL
XFILL_1_XNOR2X1_36 gnd vdd FILL
XFILL_1_XNOR2X1_25 gnd vdd FILL
XFILL_1_XNOR2X1_14 gnd vdd FILL
XFILL_1_XNOR2X1_58 gnd vdd FILL
XFILL_1_XNOR2X1_47 gnd vdd FILL
XFILL_1_XNOR2X1_69 gnd vdd FILL
XFILL_0_BUFX2_191 gnd vdd FILL
XFILL_0_BUFX2_180 gnd vdd FILL
XFILL_1_DFFPOSX1_1 gnd vdd FILL
XFILL_4_DFFPOSX1_403 gnd vdd FILL
XFILL_4_DFFPOSX1_414 gnd vdd FILL
XFILL_16_14_0 gnd vdd FILL
XFILL_4_DFFPOSX1_425 gnd vdd FILL
XFILL_4_DFFPOSX1_436 gnd vdd FILL
XFILL_4_DFFPOSX1_458 gnd vdd FILL
XFILL_4_DFFPOSX1_469 gnd vdd FILL
XFILL_4_DFFPOSX1_447 gnd vdd FILL
XFILL_1_BUFX2_315 gnd vdd FILL
XFILL_1_BUFX2_304 gnd vdd FILL
XFILL_1_BUFX2_348 gnd vdd FILL
XFILL_1_BUFX2_359 gnd vdd FILL
XOAI21X1_310 BUFX4_134/Y BUFX4_42/Y BUFX2_1020/A gnd OAI21X1_311/C vdd OAI21X1
XOAI21X1_321 INVX2_4/Y INVX8_2/A OAI21X1_321/C gnd OAI21X1_321/Y vdd OAI21X1
XOAI21X1_332 BUFX4_320/Y INVX2_11/Y NAND2X1_76/Y gnd OAI21X1_332/Y vdd OAI21X1
XOAI21X1_354 BUFX4_378/Y INVX2_22/Y NAND2X1_98/Y gnd OAI21X1_354/Y vdd OAI21X1
XOAI21X1_365 BUFX4_319/Y INVX2_26/Y OAI21X1_365/C gnd OAI21X1_365/Y vdd OAI21X1
XOAI21X1_343 BUFX4_388/Y INVX4_6/Y NAND2X1_87/Y gnd OAI21X1_343/Y vdd OAI21X1
XOAI21X1_387 BUFX4_316/Y INVX1_4/Y OAI21X1_387/C gnd OAI21X1_387/Y vdd OAI21X1
XOAI21X1_398 INVX1_7/A NOR2X1_3/B OAI21X1_398/C gnd OAI21X1_399/A vdd OAI21X1
XOAI21X1_376 BUFX4_345/Y INVX4_22/Y OAI21X1_376/C gnd OAI21X1_376/Y vdd OAI21X1
XDFFPOSX1_290 BUFX2_964/A CLKBUF1_4/Y OAI21X1_197/Y gnd vdd DFFPOSX1
XFILL_3_NOR3X1_10 gnd vdd FILL
XFILL_34_15_0 gnd vdd FILL
XNAND2X1_371 BUFX2_294/A BUFX4_211/Y gnd OAI21X1_877/C vdd NAND2X1
XNAND2X1_360 BUFX4_261/Y bundle_i[9] gnd OAI21X1_866/C vdd NAND2X1
XNAND2X1_382 BUFX2_297/A BUFX4_193/Y gnd OAI21X1_888/C vdd NAND2X1
XNAND2X1_393 BUFX2_309/A BUFX4_237/Y gnd OAI21X1_899/C vdd NAND2X1
XFILL_4_DFFPOSX1_981 gnd vdd FILL
XFILL_4_DFFPOSX1_970 gnd vdd FILL
XFILL_4_DFFPOSX1_992 gnd vdd FILL
XFILL_0_INVX1_103 gnd vdd FILL
XFILL_1_AOI21X1_14 gnd vdd FILL
XFILL_0_INVX1_125 gnd vdd FILL
XFILL_0_INVX1_136 gnd vdd FILL
XFILL_0_INVX1_114 gnd vdd FILL
XFILL_0_INVX1_147 gnd vdd FILL
XFILL_0_INVX1_169 gnd vdd FILL
XFILL_1_AOI21X1_25 gnd vdd FILL
XFILL_1_AOI21X1_36 gnd vdd FILL
XFILL_0_INVX1_158 gnd vdd FILL
XFILL_1_AOI21X1_47 gnd vdd FILL
XFILL_1_AOI21X1_58 gnd vdd FILL
XFILL_5_DFFPOSX1_109 gnd vdd FILL
XFILL_1_BUFX2_860 gnd vdd FILL
XFILL_1_BUFX2_871 gnd vdd FILL
XFILL_2_NOR3X1_2 gnd vdd FILL
XFILL_1_BUFX2_882 gnd vdd FILL
XFILL_1_OAI21X1_1804 gnd vdd FILL
XOAI21X1_1628 INVX2_131/Y BUFX4_203/Y NAND2X1_696/Y gnd DFFPOSX1_18/D vdd OAI21X1
XOAI21X1_1639 INVX2_142/Y BUFX4_209/Y NAND2X1_707/Y gnd DFFPOSX1_29/D vdd OAI21X1
XOAI21X1_1606 BUFX4_326/Y INVX2_142/Y NAND2X1_675/Y gnd OAI21X1_1606/Y vdd OAI21X1
XOAI21X1_1617 INVX2_120/Y BUFX4_192/Y NAND2X1_685/Y gnd DFFPOSX1_7/D vdd OAI21X1
XFILL_1_OAI21X1_1815 gnd vdd FILL
XFILL_3_DFFPOSX1_582 gnd vdd FILL
XFILL_3_DFFPOSX1_560 gnd vdd FILL
XFILL_1_OAI21X1_1826 gnd vdd FILL
XFILL_3_DFFPOSX1_571 gnd vdd FILL
XFILL_0_OAI21X1_628 gnd vdd FILL
XFILL_0_OAI21X1_606 gnd vdd FILL
XFILL_3_DFFPOSX1_593 gnd vdd FILL
XFILL_0_OAI21X1_617 gnd vdd FILL
XFILL_0_OAI21X1_639 gnd vdd FILL
XFILL_1_AND2X2_29 gnd vdd FILL
XFILL_1_AND2X2_18 gnd vdd FILL
XFILL_0_NAND2X1_601 gnd vdd FILL
XFILL_36_6_0 gnd vdd FILL
XFILL_0_OAI21X1_1405 gnd vdd FILL
XFILL_0_NAND2X1_634 gnd vdd FILL
XFILL_0_NAND2X1_623 gnd vdd FILL
XFILL_0_NAND2X1_645 gnd vdd FILL
XFILL_0_NAND2X1_612 gnd vdd FILL
XFILL_0_NAND2X1_667 gnd vdd FILL
XFILL_2_DFFPOSX1_150 gnd vdd FILL
XFILL_0_NAND2X1_678 gnd vdd FILL
XBUFX2_270 INVX1_62/A gnd instr1_o[14] vdd BUFX2
XFILL_0_OAI21X1_1427 gnd vdd FILL
XFILL_0_OAI21X1_1416 gnd vdd FILL
XFILL_0_OAI21X1_1438 gnd vdd FILL
XFILL_2_DFFPOSX1_161 gnd vdd FILL
XFILL_0_OAI21X1_1449 gnd vdd FILL
XFILL_2_DFFPOSX1_172 gnd vdd FILL
XBUFX2_281 INVX1_72/A gnd instr1_o[4] vdd BUFX2
XFILL_0_NAND2X1_656 gnd vdd FILL
XFILL_0_NAND2X1_689 gnd vdd FILL
XFILL_2_DFFPOSX1_194 gnd vdd FILL
XFILL_2_DFFPOSX1_183 gnd vdd FILL
XBUFX2_292 INVX1_54/A gnd instr1_o[22] vdd BUFX2
XFILL_5_DFFPOSX1_621 gnd vdd FILL
XFILL_5_DFFPOSX1_610 gnd vdd FILL
XFILL_5_DFFPOSX1_654 gnd vdd FILL
XFILL_5_DFFPOSX1_632 gnd vdd FILL
XFILL_5_DFFPOSX1_643 gnd vdd FILL
XFILL_5_DFFPOSX1_687 gnd vdd FILL
XFILL_5_DFFPOSX1_665 gnd vdd FILL
XFILL_5_DFFPOSX1_676 gnd vdd FILL
XFILL_5_DFFPOSX1_698 gnd vdd FILL
XFILL_4_DFFPOSX1_211 gnd vdd FILL
XFILL_4_DFFPOSX1_200 gnd vdd FILL
XFILL_4_DFFPOSX1_244 gnd vdd FILL
XFILL_4_DFFPOSX1_222 gnd vdd FILL
XFILL_4_DFFPOSX1_233 gnd vdd FILL
XFILL_4_DFFPOSX1_255 gnd vdd FILL
XFILL_4_DFFPOSX1_266 gnd vdd FILL
XFILL_4_DFFPOSX1_277 gnd vdd FILL
XFILL_4_DFFPOSX1_288 gnd vdd FILL
XFILL_27_6_0 gnd vdd FILL
XFILL_4_DFFPOSX1_299 gnd vdd FILL
XFILL_2_6_0 gnd vdd FILL
XFILL_2_BUFX4_343 gnd vdd FILL
XFILL_2_CLKBUF1_70 gnd vdd FILL
XFILL_2_BUFX4_376 gnd vdd FILL
XFILL_2_CLKBUF1_81 gnd vdd FILL
XFILL_2_CLKBUF1_92 gnd vdd FILL
XFILL_1_BUFX2_101 gnd vdd FILL
XFILL_1_BUFX2_123 gnd vdd FILL
XFILL_1_BUFX2_112 gnd vdd FILL
XOAI21X1_140 BUFX4_94/Y BUFX4_386/Y BUFX2_933/A gnd OAI21X1_141/C vdd OAI21X1
XFILL_1_BUFX2_156 gnd vdd FILL
XFILL_1_BUFX2_167 gnd vdd FILL
XFILL_10_5_0 gnd vdd FILL
XFILL_1_BUFX2_145 gnd vdd FILL
XOAI21X1_162 BUFX4_110/Y OAI21X1_1/A BUFX2_945/A gnd OAI21X1_163/C vdd OAI21X1
XFILL_0_BUFX2_916 gnd vdd FILL
XOAI21X1_173 BUFX4_164/Y INVX2_196/Y OAI21X1_173/C gnd OAI21X1_173/Y vdd OAI21X1
XFILL_0_BUFX2_905 gnd vdd FILL
XFILL_23_12_1 gnd vdd FILL
XOAI21X1_151 BUFX4_141/Y INVX2_185/Y OAI21X1_151/C gnd OAI21X1_151/Y vdd OAI21X1
XOAI21X1_184 BUFX4_10/A BUFX4_359/Y BUFX2_957/A gnd OAI21X1_185/C vdd OAI21X1
XOAI21X1_195 BUFX4_159/Y INVX2_5/Y OAI21X1_195/C gnd OAI21X1_195/Y vdd OAI21X1
XINVX1_204 OR2X2_19/A gnd INVX1_204/Y vdd INVX1
XFILL_0_BUFX2_938 gnd vdd FILL
XINVX1_215 INVX1_215/A gnd INVX1_215/Y vdd INVX1
XFILL_0_BUFX2_949 gnd vdd FILL
XFILL_0_BUFX2_927 gnd vdd FILL
XINVX1_226 INVX1_226/A gnd INVX1_226/Y vdd INVX1
XFILL_6_DFFPOSX1_349 gnd vdd FILL
XFILL_6_DFFPOSX1_338 gnd vdd FILL
XNAND2X1_15 BUFX2_902/A BUFX4_219/Y gnd OAI21X1_15/C vdd NAND2X1
XFILL_2_INVX8_5 gnd vdd FILL
XNAND2X1_59 BUFX2_888/A BUFX4_219/Y gnd OAI21X1_59/C vdd NAND2X1
XNAND2X1_26 BUFX2_851/A BUFX4_219/Y gnd OAI21X1_26/C vdd NAND2X1
XNAND2X1_48 BUFX2_876/A BUFX4_190/Y gnd OAI21X1_48/C vdd NAND2X1
XNAND2X1_37 BUFX2_863/A BUFX4_189/Y gnd OAI21X1_37/C vdd NAND2X1
XFILL_0_XNOR2X1_11 gnd vdd FILL
XFILL_0_XNOR2X1_33 gnd vdd FILL
XFILL_0_XNOR2X1_44 gnd vdd FILL
XFILL_0_XNOR2X1_22 gnd vdd FILL
XNAND2X1_190 OAI21X1_438/Y NAND3X1_2/Y gnd OAI21X1_439/A vdd NAND2X1
XFILL_0_XNOR2X1_77 gnd vdd FILL
XFILL_0_XNOR2X1_66 gnd vdd FILL
XFILL_0_XNOR2X1_55 gnd vdd FILL
XFILL_18_6_0 gnd vdd FILL
XFILL_0_XNOR2X1_88 gnd vdd FILL
XFILL_0_XNOR2X1_99 gnd vdd FILL
XFILL_28_11_1 gnd vdd FILL
XFILL_0_BUFX4_220 gnd vdd FILL
XFILL_0_BUFX4_231 gnd vdd FILL
XOAI21X1_1414 BUFX4_146/Y BUFX4_70/Y BUFX2_195/A gnd OAI21X1_1415/C vdd OAI21X1
XOAI21X1_1403 NOR2X1_216/A INVX4_50/Y OAI21X1_1403/C gnd OAI21X1_1405/A vdd OAI21X1
XFILL_0_BUFX4_242 gnd vdd FILL
XFILL_1_OAI21X1_1623 gnd vdd FILL
XFILL_1_OAI21X1_1601 gnd vdd FILL
XOAI21X1_1425 INVX1_220/Y bundleAddress_i[49] BUFX4_288/Y gnd OAI21X1_1427/A vdd OAI21X1
XFILL_0_BUFX4_253 gnd vdd FILL
XOAI21X1_1436 NOR2X1_220/B NOR2X1_220/A INVX2_69/Y gnd NAND2X1_628/A vdd OAI21X1
XFILL_0_BUFX4_275 gnd vdd FILL
XOAI21X1_1447 XNOR2X1_94/Y INVX8_2/A OAI21X1_1447/C gnd OAI21X1_1447/Y vdd OAI21X1
XFILL_0_BUFX4_264 gnd vdd FILL
XFILL_1_OAI21X1_1612 gnd vdd FILL
XFILL_1_OAI21X1_1667 gnd vdd FILL
XFILL_1_OAI21X1_1634 gnd vdd FILL
XOAI21X1_1458 INVX4_51/Y INVX1_189/A INVX2_71/Y gnd NAND2X1_633/A vdd OAI21X1
XOAI21X1_1469 BUFX4_157/Y BUFX4_53/Y BUFX2_215/A gnd OAI21X1_1470/C vdd OAI21X1
XFILL_0_BUFX4_297 gnd vdd FILL
XFILL_0_BUFX4_286 gnd vdd FILL
XNOR3X1_3 NOR3X1_3/A NOR3X1_3/B NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XFILL_1_OAI21X1_1656 gnd vdd FILL
XFILL_3_DFFPOSX1_390 gnd vdd FILL
XFILL_1_OAI21X1_1645 gnd vdd FILL
XFILL_0_OAI21X1_403 gnd vdd FILL
XFILL_1_OAI21X1_1678 gnd vdd FILL
XFILL_1_OAI21X1_1689 gnd vdd FILL
XFILL_1_OAI21X1_607 gnd vdd FILL
XFILL_1_OAI21X1_618 gnd vdd FILL
XFILL_0_OAI21X1_447 gnd vdd FILL
XFILL_0_OAI21X1_414 gnd vdd FILL
XFILL_0_OAI21X1_436 gnd vdd FILL
XFILL_0_OAI21X1_425 gnd vdd FILL
XFILL_1_OAI21X1_629 gnd vdd FILL
XFILL_0_OAI21X1_458 gnd vdd FILL
XFILL_0_OAI21X1_469 gnd vdd FILL
XFILL_3_DFFPOSX1_1011 gnd vdd FILL
XFILL_0_INVX4_50 gnd vdd FILL
XFILL_3_DFFPOSX1_1000 gnd vdd FILL
XFILL_3_DFFPOSX1_1022 gnd vdd FILL
XFILL_6_DFFPOSX1_850 gnd vdd FILL
XFILL_6_DFFPOSX1_861 gnd vdd FILL
XXNOR2X1_90 INVX4_50/A bundleAddress_i[57] gnd XNOR2X1_90/Y vdd XNOR2X1
XFILL_3_12_1 gnd vdd FILL
XFILL_1_XNOR2X1_2 gnd vdd FILL
XFILL_0_OAI21X1_1213 gnd vdd FILL
XFILL_0_OAI21X1_1224 gnd vdd FILL
XFILL_0_NAND2X1_431 gnd vdd FILL
XFILL_1_NAND2X1_624 gnd vdd FILL
XFILL_0_NAND2X1_420 gnd vdd FILL
XFILL_0_OAI21X1_1202 gnd vdd FILL
XFILL_1_NAND2X1_602 gnd vdd FILL
XFILL_0_NAND2X1_442 gnd vdd FILL
XFILL_0_NAND2X1_453 gnd vdd FILL
XFILL_0_NAND2X1_475 gnd vdd FILL
XFILL_0_DFFPOSX1_814 gnd vdd FILL
XFILL_1_NAND2X1_657 gnd vdd FILL
XFILL_0_OAI21X1_1257 gnd vdd FILL
XFILL_0_NAND2X1_486 gnd vdd FILL
XFILL_0_OAI21X1_1235 gnd vdd FILL
XFILL_0_OAI21X1_1246 gnd vdd FILL
XFILL_0_DFFPOSX1_825 gnd vdd FILL
XFILL_0_NAND2X1_464 gnd vdd FILL
XFILL_0_DFFPOSX1_803 gnd vdd FILL
XFILL_1_NAND2X1_646 gnd vdd FILL
XFILL_0_NAND2X1_497 gnd vdd FILL
XFILL_0_DFFPOSX1_836 gnd vdd FILL
XFILL_0_OAI21X1_1279 gnd vdd FILL
XFILL_0_DFFPOSX1_858 gnd vdd FILL
XFILL_0_OAI21X1_1268 gnd vdd FILL
XFILL_0_DFFPOSX1_847 gnd vdd FILL
XFILL_0_DFFPOSX1_869 gnd vdd FILL
XFILL_5_DFFPOSX1_462 gnd vdd FILL
XFILL_5_DFFPOSX1_451 gnd vdd FILL
XFILL_5_DFFPOSX1_440 gnd vdd FILL
XFILL_5_DFFPOSX1_484 gnd vdd FILL
XFILL_5_DFFPOSX1_495 gnd vdd FILL
XFILL_5_DFFPOSX1_473 gnd vdd FILL
XFILL_0_AOI21X1_22 gnd vdd FILL
XFILL_0_AOI21X1_11 gnd vdd FILL
XFILL_0_AOI21X1_66 gnd vdd FILL
XFILL_0_AOI21X1_44 gnd vdd FILL
XFILL_0_AOI21X1_33 gnd vdd FILL
XFILL_0_AOI21X1_55 gnd vdd FILL
XFILL_2_CLKBUF1_2 gnd vdd FILL
XFILL_0_OAI21X1_970 gnd vdd FILL
XFILL_0_OAI21X1_992 gnd vdd FILL
XFILL_0_OAI21X1_981 gnd vdd FILL
XFILL_8_11_1 gnd vdd FILL
XFILL_2_OAI21X1_1318 gnd vdd FILL
XFILL_2_DFFPOSX1_919 gnd vdd FILL
XFILL_2_DFFPOSX1_908 gnd vdd FILL
XFILL_6_DFFPOSX1_1004 gnd vdd FILL
XFILL_0_OAI21X1_1791 gnd vdd FILL
XFILL_0_OAI21X1_1780 gnd vdd FILL
XFILL_0_BUFX2_702 gnd vdd FILL
XFILL_0_BUFX2_713 gnd vdd FILL
XFILL_0_NOR2X1_42 gnd vdd FILL
XFILL_0_BUFX2_724 gnd vdd FILL
XFILL_0_NOR2X1_20 gnd vdd FILL
XFILL_0_NOR2X1_31 gnd vdd FILL
XFILL_0_BUFX2_746 gnd vdd FILL
XFILL_0_BUFX2_757 gnd vdd FILL
XFILL_0_NOR2X1_53 gnd vdd FILL
XFILL_1_DFFPOSX1_509 gnd vdd FILL
XFILL_0_NOR2X1_64 gnd vdd FILL
XFILL_0_NOR2X1_75 gnd vdd FILL
XFILL_0_BUFX2_735 gnd vdd FILL
XFILL_0_BUFX2_768 gnd vdd FILL
XFILL_0_NOR2X1_97 gnd vdd FILL
XFILL_0_NOR2X1_86 gnd vdd FILL
XFILL_0_BUFX2_779 gnd vdd FILL
XFILL_6_DFFPOSX1_124 gnd vdd FILL
XFILL_6_DFFPOSX1_135 gnd vdd FILL
XFILL_6_DFFPOSX1_102 gnd vdd FILL
XFILL_6_DFFPOSX1_113 gnd vdd FILL
XFILL_3_DFFPOSX1_8 gnd vdd FILL
XFILL_6_DFFPOSX1_146 gnd vdd FILL
XBUFX4_310 BUFX4_310/A gnd BUFX4_310/Y vdd BUFX4
XBUFX4_321 BUFX4_376/A gnd BUFX4_321/Y vdd BUFX4
XFILL_14_17_1 gnd vdd FILL
XFILL_2_OAI21X1_1830 gnd vdd FILL
XBUFX4_332 BUFX4_380/A gnd BUFX4_332/Y vdd BUFX4
XBUFX4_343 BUFX4_384/A gnd BUFX4_343/Y vdd BUFX4
XBUFX4_354 BUFX4_378/A gnd BUFX4_354/Y vdd BUFX4
XBUFX4_376 BUFX4_376/A gnd BUFX4_376/Y vdd BUFX4
XBUFX4_365 BUFX4_388/A gnd BUFX4_365/Y vdd BUFX4
XBUFX4_387 BUFX4_388/A gnd BUFX4_387/Y vdd BUFX4
XFILL_34_9_1 gnd vdd FILL
XFILL_33_4_0 gnd vdd FILL
XFILL_26_2 gnd vdd FILL
XFILL_19_1 gnd vdd FILL
XOAI21X1_909 BUFX4_126/Y INVX1_109/Y OAI21X1_909/C gnd OAI21X1_909/Y vdd OAI21X1
XFILL_0_NAND2X1_8 gnd vdd FILL
XOAI21X1_1222 INVX1_183/A NOR2X1_124/B OAI21X1_1222/C gnd OAI21X1_1224/A vdd OAI21X1
XOAI21X1_1211 BUFX4_125/Y INVX2_55/Y OAI21X1_1211/C gnd OAI21X1_1211/Y vdd OAI21X1
XOAI21X1_1200 NAND3X1_51/Y INVX1_199/Y BUFX4_242/Y gnd OAI21X1_1201/A vdd OAI21X1
XDFFPOSX1_812 BUFX2_99/A CLKBUF1_101/Y OAI21X1_1106/Y gnd vdd DFFPOSX1
XOAI21X1_1233 XNOR2X1_74/Y BUFX4_132/Y OAI21X1_1233/C gnd OAI21X1_1233/Y vdd OAI21X1
XOAI21X1_1255 OAI21X1_1255/A BUFX4_127/Y OAI21X1_1255/C gnd OAI21X1_1255/Y vdd OAI21X1
XFILL_1_OAI21X1_1431 gnd vdd FILL
XFILL_1_OAI21X1_1420 gnd vdd FILL
XDFFPOSX1_823 BUFX2_72/A CLKBUF1_59/Y OAI21X1_1129/Y gnd vdd DFFPOSX1
XOAI21X1_1244 BUFX4_109/Y BUFX4_334/Y BUFX2_134/A gnd OAI21X1_1245/C vdd OAI21X1
XFILL_1_OAI21X1_1442 gnd vdd FILL
XDFFPOSX1_801 BUFX2_54/A CLKBUF1_71/Y OAI21X1_1093/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_222 gnd vdd FILL
XFILL_0_OAI21X1_200 gnd vdd FILL
XFILL_1_OAI21X1_1475 gnd vdd FILL
XDFFPOSX1_856 BUFX2_108/A CLKBUF1_21/Y OAI21X1_1178/Y gnd vdd DFFPOSX1
XDFFPOSX1_834 BUFX2_84/A CLKBUF1_55/Y OAI21X1_1146/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1464 gnd vdd FILL
XOAI21X1_1288 BUFX4_109/Y BUFX4_317/Y BUFX2_151/A gnd OAI21X1_1290/C vdd OAI21X1
XOAI21X1_1277 NAND2X1_601/Y BUFX4_174/Y OAI21X1_1277/C gnd OAI21X1_1277/Y vdd OAI21X1
XDFFPOSX1_845 BUFX2_96/A CLKBUF1_28/Y OAI21X1_1161/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1453 gnd vdd FILL
XOAI21X1_1266 BUFX4_4/Y BUFX4_324/Y BUFX2_142/A gnd OAI21X1_1267/C vdd OAI21X1
XFILL_0_OAI21X1_211 gnd vdd FILL
XFILL_0_OAI21X1_255 gnd vdd FILL
XDFFPOSX1_889 BUFX2_138/A CLKBUF1_59/Y OAI21X1_1258/Y gnd vdd DFFPOSX1
XDFFPOSX1_878 BUFX2_185/A CLKBUF1_31/Y OAI21X1_1224/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_233 gnd vdd FILL
XOAI21X1_1299 AND2X2_30/Y OAI21X1_1299/B OAI21X1_1299/C gnd OAI21X1_1299/Y vdd OAI21X1
XFILL_0_OAI21X1_244 gnd vdd FILL
XDFFPOSX1_867 BUFX2_120/A CLKBUF1_69/Y OAI21X1_1199/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_426 gnd vdd FILL
XFILL_1_OAI21X1_1486 gnd vdd FILL
XFILL_1_OAI21X1_1497 gnd vdd FILL
XINVX2_17 bundleStartMajId_i[47] gnd INVX2_17/Y vdd INVX2
XFILL_1_OAI21X1_415 gnd vdd FILL
XFILL_1_OAI21X1_404 gnd vdd FILL
XFILL_0_OAI21X1_277 gnd vdd FILL
XFILL_0_OAI21X1_288 gnd vdd FILL
XFILL_0_OAI21X1_266 gnd vdd FILL
XINVX2_39 bundleStartMajId_i[0] gnd INVX2_39/Y vdd INVX2
XFILL_1_OAI21X1_437 gnd vdd FILL
XFILL_19_16_1 gnd vdd FILL
XFILL_1_OAI21X1_459 gnd vdd FILL
XINVX2_28 bundleStartMajId_i[21] gnd INVX2_28/Y vdd INVX2
XFILL_1_OAI21X1_448 gnd vdd FILL
XFILL_0_OAI21X1_299 gnd vdd FILL
XFILL_32_18_1 gnd vdd FILL
XFILL_13_12_0 gnd vdd FILL
XFILL_1_INVX4_28 gnd vdd FILL
XFILL_1_INVX4_17 gnd vdd FILL
XFILL_0_OAI21X1_1032 gnd vdd FILL
XFILL_1_NAND2X1_432 gnd vdd FILL
XFILL_0_OAI21X1_1021 gnd vdd FILL
XFILL_0_DFFPOSX1_600 gnd vdd FILL
XFILL_25_9_1 gnd vdd FILL
XFILL_1_INVX4_39 gnd vdd FILL
XFILL_0_NAND2X1_261 gnd vdd FILL
XFILL_0_NAND2X1_250 gnd vdd FILL
XFILL_1_NAND2X1_421 gnd vdd FILL
XFILL_0_9_1 gnd vdd FILL
XFILL_0_OAI21X1_1010 gnd vdd FILL
XFILL_1_BUFX4_207 gnd vdd FILL
XFILL_0_OAI21X1_1043 gnd vdd FILL
XFILL_1_BUFX4_218 gnd vdd FILL
XFILL_0_DFFPOSX1_633 gnd vdd FILL
XFILL_0_OAI21X1_1065 gnd vdd FILL
XFILL_24_4_0 gnd vdd FILL
XFILL_0_OAI21X1_1054 gnd vdd FILL
XFILL_1_NAND2X1_465 gnd vdd FILL
XFILL_0_DFFPOSX1_611 gnd vdd FILL
XFILL_0_NAND2X1_294 gnd vdd FILL
XFILL_0_NAND2X1_283 gnd vdd FILL
XFILL_0_DFFPOSX1_622 gnd vdd FILL
XFILL_1_NAND2X1_443 gnd vdd FILL
XFILL_0_NAND2X1_272 gnd vdd FILL
XFILL_0_DFFPOSX1_655 gnd vdd FILL
XFILL_1_BUFX4_229 gnd vdd FILL
XFILL_1_NAND2X1_498 gnd vdd FILL
XFILL_0_OAI21X1_1098 gnd vdd FILL
XFILL_0_DFFPOSX1_644 gnd vdd FILL
XFILL_0_DFFPOSX1_666 gnd vdd FILL
XFILL_0_OAI21X1_1076 gnd vdd FILL
XFILL_0_OAI21X1_1087 gnd vdd FILL
XFILL_0_DFFPOSX1_688 gnd vdd FILL
XFILL_0_DFFPOSX1_677 gnd vdd FILL
XFILL_0_DFFPOSX1_699 gnd vdd FILL
XFILL_5_DFFPOSX1_281 gnd vdd FILL
XFILL_5_DFFPOSX1_270 gnd vdd FILL
XFILL_5_DFFPOSX1_292 gnd vdd FILL
XFILL_37_17_1 gnd vdd FILL
XFILL_1_OAI21X1_971 gnd vdd FILL
XFILL_18_11_0 gnd vdd FILL
XFILL_1_OAI21X1_960 gnd vdd FILL
XFILL_1_OR2X2_1 gnd vdd FILL
XFILL_1_OAI21X1_982 gnd vdd FILL
XFILL_7_5_0 gnd vdd FILL
XFILL_1_OAI21X1_993 gnd vdd FILL
XFILL_31_13_0 gnd vdd FILL
XFILL_2_OAI21X1_1115 gnd vdd FILL
XBUFX2_803 BUFX2_803/A gnd tid1_o[31] vdd BUFX2
XFILL_2_DFFPOSX1_705 gnd vdd FILL
XFILL_2_DFFPOSX1_716 gnd vdd FILL
XFILL_2_DFFPOSX1_727 gnd vdd FILL
XBUFX2_836 NAND2X1_6/A gnd tid1_o[1] vdd BUFX2
XBUFX2_814 BUFX2_814/A gnd tid1_o[21] vdd BUFX2
XBUFX2_825 BUFX2_825/A gnd tid1_o[11] vdd BUFX2
XFILL_2_OAI21X1_1159 gnd vdd FILL
XFILL_2_DFFPOSX1_738 gnd vdd FILL
XBUFX2_869 BUFX2_869/A gnd tid2_o[29] vdd BUFX2
XBUFX2_847 BUFX2_847/A gnd tid2_o[49] vdd BUFX2
XBUFX2_858 BUFX2_858/A gnd tid2_o[39] vdd BUFX2
XFILL_2_DFFPOSX1_749 gnd vdd FILL
XFILL_2_NAND3X1_50 gnd vdd FILL
XFILL_16_9_1 gnd vdd FILL
XFILL_15_4_0 gnd vdd FILL
XFILL_0_NOR2X1_209 gnd vdd FILL
XMUX2X1_1 MUX2X1_1/A MUX2X1_1/B INVX8_6/A gnd MUX2X1_1/Y vdd MUX2X1
XDFFPOSX1_119 BUFX2_788/A CLKBUF1_12/Y OAI21X1_1793/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_532 gnd vdd FILL
XFILL_0_BUFX2_521 gnd vdd FILL
XDFFPOSX1_108 BUFX2_839/A CLKBUF1_56/Y OAI21X1_1782/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_510 gnd vdd FILL
XFILL_1_DFFPOSX1_306 gnd vdd FILL
XFILL_1_DFFPOSX1_328 gnd vdd FILL
XFILL_1_DFFPOSX1_317 gnd vdd FILL
XFILL_0_BUFX2_565 gnd vdd FILL
XFILL_0_BUFX2_543 gnd vdd FILL
XFILL_0_BUFX2_554 gnd vdd FILL
XCLKBUF1_2 BUFX4_88/Y gnd CLKBUF1_2/Y vdd CLKBUF1
XFILL_0_BUFX2_576 gnd vdd FILL
XFILL_1_DFFPOSX1_339 gnd vdd FILL
XFILL_0_BUFX2_598 gnd vdd FILL
XFILL_0_BUFX2_587 gnd vdd FILL
XFILL_36_12_0 gnd vdd FILL
XFILL_2_OAI21X1_1660 gnd vdd FILL
XFILL_4_CLKBUF1_11 gnd vdd FILL
XBUFX4_140 BUFX4_14/Y gnd BUFX4_140/Y vdd BUFX4
XBUFX4_151 BUFX4_18/Y gnd BUFX4_151/Y vdd BUFX4
XFILL_4_CLKBUF1_22 gnd vdd FILL
XBUFX4_162 BUFX4_14/Y gnd BUFX4_162/Y vdd BUFX4
XFILL_0_INVX1_40 gnd vdd FILL
XNOR2X1_200 INVX1_208/A NOR2X1_200/B gnd AND2X2_31/B vdd NOR2X1
XFILL_4_CLKBUF1_33 gnd vdd FILL
XFILL_0_INVX1_51 gnd vdd FILL
XBUFX4_173 BUFX4_13/Y gnd BUFX4_173/Y vdd BUFX4
XFILL_0_INVX1_84 gnd vdd FILL
XBUFX4_184 BUFX4_24/Y gnd BUFX4_184/Y vdd BUFX4
XFILL_0_INVX1_62 gnd vdd FILL
XBUFX4_195 BUFX4_23/Y gnd BUFX4_195/Y vdd BUFX4
XNOR2X1_233 BUFX4_11/Y BUFX4_344/Y gnd BUFX4_310/A vdd NOR2X1
XFILL_4_CLKBUF1_55 gnd vdd FILL
XNOR2X1_211 INVX1_216/Y NOR2X1_211/B gnd XNOR2X1_88/A vdd NOR2X1
XFILL_4_CLKBUF1_77 gnd vdd FILL
XNOR2X1_222 OR2X2_17/Y NOR2X1_222/B gnd XNOR2X1_95/A vdd NOR2X1
XFILL_4_CLKBUF1_44 gnd vdd FILL
XFILL_0_INVX1_73 gnd vdd FILL
XFILL_0_INVX1_95 gnd vdd FILL
XFILL_4_CLKBUF1_66 gnd vdd FILL
XFILL_4_CLKBUF1_99 gnd vdd FILL
XFILL_0_BUFX2_26 gnd vdd FILL
XFILL_0_BUFX2_15 gnd vdd FILL
XFILL_0_BUFX2_59 gnd vdd FILL
XFILL_0_BUFX2_37 gnd vdd FILL
XFILL_0_BUFX2_48 gnd vdd FILL
XOAI21X1_706 OAI21X1_706/A BUFX4_299/Y OAI21X1_706/C gnd OAI21X1_706/Y vdd OAI21X1
XOAI21X1_717 BUFX4_142/Y BUFX4_43/Y BUFX2_598/A gnd OAI21X1_718/C vdd OAI21X1
XOAI21X1_728 BUFX4_133/Y BUFX4_27/Y BUFX2_602/A gnd OAI21X1_729/C vdd OAI21X1
XOAI21X1_739 XNOR2X1_46/A INVX4_12/Y INVX4_13/Y gnd OAI21X1_739/Y vdd OAI21X1
XOAI21X1_1030 BUFX4_137/Y BUFX4_60/Y BUFX2_379/A gnd OAI21X1_1031/C vdd OAI21X1
XFILL_1_OAI21X1_1250 gnd vdd FILL
XOAI21X1_1041 BUFX4_347/Y INVX2_58/Y NAND2X1_407/Y gnd OAI21X1_1041/Y vdd OAI21X1
XOAI21X1_1052 BUFX4_356/Y INVX4_34/Y NAND2X1_418/Y gnd OAI21X1_1052/Y vdd OAI21X1
XOAI21X1_1063 BUFX4_317/Y INVX2_72/Y NAND2X1_429/Y gnd OAI21X1_1063/Y vdd OAI21X1
XDFFPOSX1_620 INVX1_49/A CLKBUF1_54/Y OAI21X1_848/Y gnd vdd DFFPOSX1
XDFFPOSX1_631 INVX1_60/A CLKBUF1_10/Y OAI21X1_859/Y gnd vdd DFFPOSX1
XDFFPOSX1_664 BUFX2_301/A CLKBUF1_96/Y OAI21X1_892/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_840 gnd vdd FILL
XFILL_1_OAI21X1_1261 gnd vdd FILL
XFILL_1_OAI21X1_201 gnd vdd FILL
XFILL_1_DFFPOSX1_851 gnd vdd FILL
XDFFPOSX1_642 INVX1_71/A CLKBUF1_82/Y OAI21X1_870/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1283 gnd vdd FILL
XOAI21X1_1085 BUFX4_342/Y INVX2_83/Y NAND2X1_451/Y gnd OAI21X1_1085/Y vdd OAI21X1
XOAI21X1_1096 BUFX4_357/Y INVX1_181/Y NAND2X1_462/Y gnd OAI21X1_1096/Y vdd OAI21X1
XFILL_1_OAI21X1_1272 gnd vdd FILL
XDFFPOSX1_675 BUFX2_313/A CLKBUF1_13/Y OAI21X1_903/Y gnd vdd DFFPOSX1
XDFFPOSX1_653 BUFX2_320/A CLKBUF1_82/Y OAI21X1_881/Y gnd vdd DFFPOSX1
XOAI21X1_1074 BUFX4_384/Y INVX2_78/Y NAND2X1_440/Y gnd OAI21X1_1074/Y vdd OAI21X1
XFILL_1_OAI21X1_234 gnd vdd FILL
XFILL_1_DFFPOSX1_884 gnd vdd FILL
XFILL_1_OAI21X1_223 gnd vdd FILL
XFILL_1_OAI21X1_1294 gnd vdd FILL
XFILL_1_DFFPOSX1_873 gnd vdd FILL
XFILL_1_OAI21X1_212 gnd vdd FILL
XNAND2X1_701 BUFX2_692/A BUFX4_233/Y gnd NAND2X1_701/Y vdd NAND2X1
XNAND2X1_712 BUFX2_705/A BUFX4_225/Y gnd NAND2X1_712/Y vdd NAND2X1
XDFFPOSX1_697 BUFX2_334/A CLKBUF1_52/Y OAI21X1_943/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_862 gnd vdd FILL
XDFFPOSX1_686 BUFX2_353/A CLKBUF1_37/Y OAI21X1_921/Y gnd vdd DFFPOSX1
XNAND2X1_734 BUFX2_788/A BUFX4_353/Y gnd NAND2X1_734/Y vdd NAND2X1
XNAND2X1_745 BUFX2_801/A BUFX4_336/Y gnd NAND2X1_745/Y vdd NAND2X1
XFILL_1_OAI21X1_267 gnd vdd FILL
XFILL_1_OAI21X1_278 gnd vdd FILL
XFILL_1_OAI21X1_245 gnd vdd FILL
XFILL_1_DFFPOSX1_895 gnd vdd FILL
XFILL_2_OAI21X1_416 gnd vdd FILL
XFILL_1_OAI21X1_256 gnd vdd FILL
XNAND2X1_723 BUFX2_839/A BUFX4_315/Y gnd NAND2X1_723/Y vdd NAND2X1
XFILL_0_NOR2X1_6 gnd vdd FILL
XFILL_1_OAI21X1_289 gnd vdd FILL
XNAND2X1_767 BUFX2_825/A OAI21X1_2/A gnd NAND2X1_767/Y vdd NAND2X1
XNAND2X1_756 BUFX2_813/A BUFX4_343/Y gnd NAND2X1_756/Y vdd NAND2X1
XFILL_2_XNOR2X1_18 gnd vdd FILL
XFILL_2_XNOR2X1_29 gnd vdd FILL
XFILL_1_NAND2X1_240 gnd vdd FILL
XFILL_1_NAND2X1_284 gnd vdd FILL
XFILL_1_NAND2X1_273 gnd vdd FILL
XFILL_0_DFFPOSX1_430 gnd vdd FILL
XFILL_0_DFFPOSX1_441 gnd vdd FILL
XFILL_2_DFFPOSX1_5 gnd vdd FILL
XFILL_0_DFFPOSX1_463 gnd vdd FILL
XFILL_1_NAND2X1_295 gnd vdd FILL
XFILL_0_DFFPOSX1_485 gnd vdd FILL
XFILL_0_DFFPOSX1_452 gnd vdd FILL
XFILL_0_DFFPOSX1_474 gnd vdd FILL
XINVX8_4 INVX8_4/A gnd INVX8_4/Y vdd INVX8
XFILL_0_DFFPOSX1_496 gnd vdd FILL
XFILL_3_DFFPOSX1_901 gnd vdd FILL
XFILL_3_DFFPOSX1_923 gnd vdd FILL
XFILL_3_DFFPOSX1_912 gnd vdd FILL
XFILL_3_DFFPOSX1_945 gnd vdd FILL
XFILL_3_DFFPOSX1_934 gnd vdd FILL
XFILL_3_DFFPOSX1_956 gnd vdd FILL
XFILL_3_DFFPOSX1_967 gnd vdd FILL
XFILL_20_10_1 gnd vdd FILL
XFILL_3_DFFPOSX1_978 gnd vdd FILL
XFILL_3_DFFPOSX1_989 gnd vdd FILL
XDFFPOSX1_90 BUFX2_760/A CLKBUF1_16/Y DFFPOSX1_90/D gnd vdd DFFPOSX1
XBUFX4_35 BUFX4_55/A gnd BUFX4_35/Y vdd BUFX4
XBUFX4_24 BUFX4_26/A gnd BUFX4_24/Y vdd BUFX4
XBUFX4_13 INVX8_6/Y gnd BUFX4_13/Y vdd BUFX4
XFILL_1_OAI21X1_790 gnd vdd FILL
XBUFX4_57 BUFX4_82/A gnd BUFX4_57/Y vdd BUFX4
XBUFX4_46 BUFX4_81/A gnd BUFX4_46/Y vdd BUFX4
XBUFX4_68 BUFX4_73/A gnd BUFX4_68/Y vdd BUFX4
XBUFX2_611 BUFX2_611/A gnd majID4_o[31] vdd BUFX2
XBUFX4_79 BUFX4_79/A gnd BUFX4_79/Y vdd BUFX4
XFILL_2_DFFPOSX1_513 gnd vdd FILL
XFILL_2_DFFPOSX1_502 gnd vdd FILL
XBUFX2_600 BUFX2_600/A gnd majID4_o[41] vdd BUFX2
XBUFX2_644 BUFX2_644/A gnd majID4_o[1] vdd BUFX2
XBUFX2_655 BUFX2_655/A gnd pid1_o[17] vdd BUFX2
XFILL_2_DFFPOSX1_546 gnd vdd FILL
XBUFX2_633 BUFX2_633/A gnd majID4_o[11] vdd BUFX2
XFILL_2_DFFPOSX1_535 gnd vdd FILL
XBUFX2_622 BUFX2_622/A gnd majID4_o[21] vdd BUFX2
XFILL_2_DFFPOSX1_524 gnd vdd FILL
XBUFX2_688 BUFX2_688/A gnd pid2_o[16] vdd BUFX2
XFILL_2_DFFPOSX1_568 gnd vdd FILL
XFILL_2_DFFPOSX1_579 gnd vdd FILL
XBUFX2_666 BUFX2_666/A gnd pid1_o[7] vdd BUFX2
XFILL_2_DFFPOSX1_557 gnd vdd FILL
XBUFX2_677 BUFX2_677/A gnd pid1_o[25] vdd BUFX2
XBUFX2_699 BUFX2_699/A gnd pid2_o[6] vdd BUFX2
XFILL_31_7_1 gnd vdd FILL
XFILL_30_2_0 gnd vdd FILL
XFILL_22_18_0 gnd vdd FILL
XINVX2_140 bundlePid_i[8] gnd INVX2_140/Y vdd INVX2
XOR2X2_16 OR2X2_16/A OR2X2_16/B gnd OR2X2_16/Y vdd OR2X2
XFILL_0_BUFX2_340 gnd vdd FILL
XFILL_1_DFFPOSX1_103 gnd vdd FILL
XINVX2_173 bundleTid_i[36] gnd INVX2_173/Y vdd INVX2
XFILL_1_DFFPOSX1_114 gnd vdd FILL
XFILL_1_DFFPOSX1_125 gnd vdd FILL
XINVX2_162 bundleTid_i[47] gnd INVX2_162/Y vdd INVX2
XFILL_0_BUFX2_362 gnd vdd FILL
XFILL_1_DFFPOSX1_147 gnd vdd FILL
XINVX2_184 bundleTid_i[25] gnd INVX2_184/Y vdd INVX2
XFILL_1_DFFPOSX1_136 gnd vdd FILL
XFILL_0_BUFX2_373 gnd vdd FILL
XOR2X2_9 OR2X2_9/A OR2X2_9/B gnd OR2X2_9/Y vdd OR2X2
XFILL_0_BUFX2_384 gnd vdd FILL
XINVX2_151 bundleTid_i[58] gnd INVX2_151/Y vdd INVX2
XFILL_0_BUFX2_351 gnd vdd FILL
XINVX2_195 bundleTid_i[14] gnd INVX2_195/Y vdd INVX2
XFILL_0_BUFX2_395 gnd vdd FILL
XFILL_1_DFFPOSX1_158 gnd vdd FILL
XFILL_1_DFFPOSX1_169 gnd vdd FILL
XFILL_4_DFFPOSX1_607 gnd vdd FILL
XFILL_4_DFFPOSX1_618 gnd vdd FILL
XFILL_4_DFFPOSX1_629 gnd vdd FILL
XFILL_38_3_0 gnd vdd FILL
XFILL_0_10_1 gnd vdd FILL
XFILL_27_17_0 gnd vdd FILL
XFILL_22_7_1 gnd vdd FILL
XFILL_21_2_0 gnd vdd FILL
XOAI21X1_503 BUFX4_135/Y bundleStartMajId_i[62] OAI21X1_503/C gnd OAI21X1_503/Y vdd
+ OAI21X1
XOAI21X1_514 BUFX4_7/A BUFX4_365/Y BUFX2_566/A gnd OAI21X1_515/C vdd OAI21X1
XFILL_3_DFFPOSX1_208 gnd vdd FILL
XOAI21X1_525 BUFX4_2/A BUFX4_323/Y BUFX2_584/A gnd OAI21X1_526/C vdd OAI21X1
XFILL_3_DFFPOSX1_219 gnd vdd FILL
XOAI21X1_547 BUFX4_7/Y BUFX4_358/Y BUFX2_530/A gnd OAI21X1_548/C vdd OAI21X1
XOAI21X1_536 XNOR2X1_26/Y BUFX4_122/Y OAI21X1_536/C gnd OAI21X1_536/Y vdd OAI21X1
XOAI21X1_569 NOR2X1_70/B INVX4_11/Y INVX2_22/Y gnd OAI21X1_570/C vdd OAI21X1
XOAI21X1_558 BUFX4_10/A BUFX4_319/Y BUFX2_534/A gnd OAI21X1_559/C vdd OAI21X1
XDFFPOSX1_483 BUFX2_517/A CLKBUF1_65/Y NAND2X1_265/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1080 gnd vdd FILL
XDFFPOSX1_450 BUFX2_481/A CLKBUF1_50/Y OAI21X1_445/Y gnd vdd DFFPOSX1
XDFFPOSX1_461 BUFX2_493/A CLKBUF1_84/Y OAI21X1_461/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1091 gnd vdd FILL
XDFFPOSX1_472 BUFX2_505/A CLKBUF1_48/Y OAI21X1_480/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_670 gnd vdd FILL
XFILL_1_DFFPOSX1_692 gnd vdd FILL
XFILL_1_DFFPOSX1_681 gnd vdd FILL
XNAND2X1_520 INVX1_189/Y INVX1_188/A gnd INVX1_190/A vdd NAND2X1
XDFFPOSX1_494 BUFX2_523/A CLKBUF1_75/Y OAI21X1_530/Y gnd vdd DFFPOSX1
XFILL_2_OAI21X1_246 gnd vdd FILL
XNAND2X1_531 BUFX2_91/A BUFX4_202/Y gnd NAND2X1_531/Y vdd NAND2X1
XNAND2X1_553 bundleAddress_i[20] bundleAddress_i[19] gnd NOR2X1_204/A vdd NAND2X1
XNAND2X1_542 bundleAddress_i[25] NOR2X1_156/Y gnd INVX1_193/A vdd NAND2X1
XNAND2X1_597 NAND2X1_597/A NAND2X1_597/B gnd NAND2X1_597/Y vdd NAND2X1
XFILL_2_OAI21X1_279 gnd vdd FILL
XNAND2X1_564 INVX2_111/A NOR2X1_165/Y gnd NOR2X1_166/A vdd NAND2X1
XNAND2X1_586 bundleAddress_i[5] INVX1_199/A gnd NOR2X1_176/B vdd NAND2X1
XNAND2X1_575 BUFX4_242/Y NAND2X1_575/B gnd NAND2X1_575/Y vdd NAND2X1
XFILL_5_8_1 gnd vdd FILL
XFILL_29_3_0 gnd vdd FILL
XFILL_4_3_0 gnd vdd FILL
XFILL_0_AND2X2_10 gnd vdd FILL
XFILL_2_18_0 gnd vdd FILL
XFILL_0_AND2X2_32 gnd vdd FILL
XFILL_0_AND2X2_21 gnd vdd FILL
XFILL_13_7_1 gnd vdd FILL
XFILL_0_DFFPOSX1_282 gnd vdd FILL
XFILL_0_DFFPOSX1_271 gnd vdd FILL
XFILL_12_2_0 gnd vdd FILL
XFILL_0_DFFPOSX1_260 gnd vdd FILL
XFILL_0_DFFPOSX1_293 gnd vdd FILL
XFILL_3_DFFPOSX1_720 gnd vdd FILL
XFILL_3_DFFPOSX1_731 gnd vdd FILL
XFILL_3_DFFPOSX1_742 gnd vdd FILL
XFILL_3_DFFPOSX1_753 gnd vdd FILL
XFILL_3_CLKBUF1_30 gnd vdd FILL
XFILL_3_CLKBUF1_41 gnd vdd FILL
XFILL_3_DFFPOSX1_764 gnd vdd FILL
XFILL_3_CLKBUF1_74 gnd vdd FILL
XFILL_3_DFFPOSX1_775 gnd vdd FILL
XFILL_3_CLKBUF1_63 gnd vdd FILL
XFILL_3_DFFPOSX1_786 gnd vdd FILL
XFILL_3_CLKBUF1_85 gnd vdd FILL
XFILL_3_DFFPOSX1_797 gnd vdd FILL
XFILL_3_CLKBUF1_52 gnd vdd FILL
XFILL_3_CLKBUF1_96 gnd vdd FILL
XFILL_1_NOR2X1_181 gnd vdd FILL
XFILL_1_NOR2X1_192 gnd vdd FILL
XFILL_1_NOR2X1_170 gnd vdd FILL
XFILL_7_17_0 gnd vdd FILL
XFILL_2_NAND3X1_1 gnd vdd FILL
XFILL_2_DFFPOSX1_321 gnd vdd FILL
XBUFX2_430 BUFX2_430/A gnd majID1_o[21] vdd BUFX2
XFILL_2_DFFPOSX1_310 gnd vdd FILL
XFILL_11_15_1 gnd vdd FILL
XFILL_0_OAI21X1_1609 gnd vdd FILL
XBUFX2_452 BUFX2_452/A gnd majID1_o[1] vdd BUFX2
XFILL_2_DFFPOSX1_343 gnd vdd FILL
XBUFX2_441 BUFX2_441/A gnd majID1_o[11] vdd BUFX2
XFILL_2_DFFPOSX1_354 gnd vdd FILL
XFILL_2_DFFPOSX1_332 gnd vdd FILL
XBUFX2_463 BUFX2_463/A gnd majID2_o[49] vdd BUFX2
XFILL_2_DFFPOSX1_365 gnd vdd FILL
XFILL_2_DFFPOSX1_398 gnd vdd FILL
XBUFX2_485 BUFX2_485/A gnd majID2_o[29] vdd BUFX2
XFILL_2_DFFPOSX1_376 gnd vdd FILL
XBUFX2_474 BUFX2_474/A gnd majID2_o[39] vdd BUFX2
XBUFX2_496 BUFX2_496/A gnd majID2_o[19] vdd BUFX2
XFILL_2_DFFPOSX1_387 gnd vdd FILL
XFILL_5_DFFPOSX1_803 gnd vdd FILL
XFILL_5_DFFPOSX1_814 gnd vdd FILL
XFILL_5_DFFPOSX1_825 gnd vdd FILL
XFILL_5_DFFPOSX1_836 gnd vdd FILL
XFILL_5_DFFPOSX1_869 gnd vdd FILL
XFILL_5_DFFPOSX1_858 gnd vdd FILL
XFILL_5_DFFPOSX1_847 gnd vdd FILL
XFILL_1_XNOR2X1_15 gnd vdd FILL
XFILL_1_XNOR2X1_37 gnd vdd FILL
XFILL_1_XNOR2X1_26 gnd vdd FILL
XFILL_1_XNOR2X1_59 gnd vdd FILL
XFILL_1_XNOR2X1_48 gnd vdd FILL
XFILL_0_BUFX2_192 gnd vdd FILL
XFILL_0_BUFX2_170 gnd vdd FILL
XFILL_0_BUFX2_181 gnd vdd FILL
XFILL_1_DFFPOSX1_2 gnd vdd FILL
XFILL_4_DFFPOSX1_415 gnd vdd FILL
XFILL_16_14_1 gnd vdd FILL
XFILL_4_DFFPOSX1_404 gnd vdd FILL
XFILL_4_DFFPOSX1_426 gnd vdd FILL
XFILL_4_DFFPOSX1_437 gnd vdd FILL
XFILL_4_DFFPOSX1_459 gnd vdd FILL
XFILL_4_DFFPOSX1_448 gnd vdd FILL
XFILL_10_10_0 gnd vdd FILL
XFILL_1_BUFX2_327 gnd vdd FILL
XFILL_1_BUFX2_305 gnd vdd FILL
XOAI21X1_300 BUFX4_165/Y BUFX4_60/Y BUFX2_1015/A gnd OAI21X1_301/C vdd OAI21X1
XFILL_1_BUFX2_338 gnd vdd FILL
XOAI21X1_322 BUFX4_179/Y BUFX4_75/Y BUFX2_1027/A gnd OAI21X1_323/C vdd OAI21X1
XFILL_1_BUFX2_349 gnd vdd FILL
XOAI21X1_311 INVX2_201/Y BUFX4_302/Y OAI21X1_311/C gnd OAI21X1_311/Y vdd OAI21X1
XOAI21X1_355 BUFX4_319/Y INVX4_12/Y NAND2X1_99/Y gnd OAI21X1_355/Y vdd OAI21X1
XOAI21X1_333 BUFX4_355/Y INVX2_12/Y NAND2X1_77/Y gnd OAI21X1_333/Y vdd OAI21X1
XOAI21X1_344 BUFX4_355/Y INVX2_17/Y NAND2X1_88/Y gnd OAI21X1_344/Y vdd OAI21X1
XOAI21X1_366 BUFX4_351/Y NOR3X1_6/A OAI21X1_366/C gnd OAI21X1_366/Y vdd OAI21X1
XOAI21X1_388 BUFX4_351/Y INVX2_38/Y OAI21X1_388/C gnd OAI21X1_388/Y vdd OAI21X1
XOAI21X1_377 BUFX4_323/Y INVX4_23/Y OAI21X1_377/C gnd OAI21X1_377/Y vdd OAI21X1
XOAI21X1_399 OAI21X1_399/A BUFX4_222/Y OAI21X1_399/C gnd OAI21X1_399/Y vdd OAI21X1
XDFFPOSX1_291 BUFX2_965/A CLKBUF1_69/Y OAI21X1_199/Y gnd vdd DFFPOSX1
XDFFPOSX1_280 BUFX2_953/A CLKBUF1_15/Y OAI21X1_177/Y gnd vdd DFFPOSX1
XFILL_3_NOR3X1_11 gnd vdd FILL
XNAND2X1_361 BUFX4_263/Y bundle_i[8] gnd OAI21X1_867/C vdd NAND2X1
XFILL_34_15_1 gnd vdd FILL
XNAND2X1_372 BUFX2_305/A BUFX4_211/Y gnd OAI21X1_878/C vdd NAND2X1
XNAND2X1_350 BUFX4_264/Y bundle_i[19] gnd OAI21X1_856/C vdd NAND2X1
XNAND2X1_394 BUFX2_310/A BUFX4_197/Y gnd OAI21X1_900/C vdd NAND2X1
XNAND2X1_383 BUFX2_298/A BUFX4_205/Y gnd OAI21X1_889/C vdd NAND2X1
XFILL_4_DFFPOSX1_982 gnd vdd FILL
XFILL_4_DFFPOSX1_960 gnd vdd FILL
XFILL_0_INVX1_104 gnd vdd FILL
XFILL_4_DFFPOSX1_971 gnd vdd FILL
XFILL_1_AOI21X1_15 gnd vdd FILL
XFILL_4_DFFPOSX1_993 gnd vdd FILL
XFILL_0_INVX1_115 gnd vdd FILL
XFILL_0_INVX1_126 gnd vdd FILL
XFILL_0_INVX1_137 gnd vdd FILL
XFILL_1_AOI21X1_26 gnd vdd FILL
XFILL_1_AOI21X1_37 gnd vdd FILL
XFILL_1_AOI21X1_48 gnd vdd FILL
XFILL_0_INVX1_148 gnd vdd FILL
XFILL_0_INVX1_159 gnd vdd FILL
XFILL_1_AOI21X1_59 gnd vdd FILL
XFILL_1_INVX2_61 gnd vdd FILL
XFILL_1_BUFX2_861 gnd vdd FILL
XFILL_1_BUFX2_850 gnd vdd FILL
XFILL_2_NOR3X1_3 gnd vdd FILL
XOAI21X1_1629 INVX2_132/Y BUFX4_218/Y NAND2X1_697/Y gnd DFFPOSX1_19/D vdd OAI21X1
XOAI21X1_1607 BUFX4_349/Y INVX2_143/Y NAND2X1_676/Y gnd OAI21X1_1607/Y vdd OAI21X1
XFILL_1_BUFX2_894 gnd vdd FILL
XFILL_1_OAI21X1_1805 gnd vdd FILL
XOAI21X1_1618 INVX2_121/Y BUFX4_180/Y NAND2X1_686/Y gnd DFFPOSX1_8/D vdd OAI21X1
XFILL_1_OAI21X1_1816 gnd vdd FILL
XFILL_1_OAI21X1_1827 gnd vdd FILL
XFILL_3_DFFPOSX1_583 gnd vdd FILL
XFILL_3_DFFPOSX1_550 gnd vdd FILL
XFILL_3_DFFPOSX1_572 gnd vdd FILL
XFILL_3_DFFPOSX1_561 gnd vdd FILL
XFILL_0_OAI21X1_629 gnd vdd FILL
XFILL_0_OAI21X1_607 gnd vdd FILL
XFILL_3_DFFPOSX1_594 gnd vdd FILL
XFILL_0_OAI21X1_618 gnd vdd FILL
XFILL_7_1 gnd vdd FILL
XFILL_1_AND2X2_19 gnd vdd FILL
XFILL_33_10_0 gnd vdd FILL
XFILL_0_NAND2X1_602 gnd vdd FILL
XFILL_36_6_1 gnd vdd FILL
XFILL_0_NAND2X1_624 gnd vdd FILL
XFILL_0_OAI21X1_1406 gnd vdd FILL
XFILL_0_NAND2X1_635 gnd vdd FILL
XFILL_0_NAND2X1_613 gnd vdd FILL
XFILL_2_DFFPOSX1_140 gnd vdd FILL
XBUFX2_271 INVX1_63/A gnd instr1_o[13] vdd BUFX2
XFILL_0_NAND2X1_657 gnd vdd FILL
XFILL_35_1_0 gnd vdd FILL
XFILL_0_OAI21X1_1417 gnd vdd FILL
XFILL_0_OAI21X1_1428 gnd vdd FILL
XBUFX2_260 BUFX2_260/A gnd enable4_o vdd BUFX2
XFILL_2_DFFPOSX1_173 gnd vdd FILL
XFILL_0_NAND2X1_668 gnd vdd FILL
XFILL_2_DFFPOSX1_151 gnd vdd FILL
XFILL_0_OAI21X1_1439 gnd vdd FILL
XFILL_0_NAND2X1_646 gnd vdd FILL
XFILL_2_DFFPOSX1_162 gnd vdd FILL
XFILL_2_DFFPOSX1_195 gnd vdd FILL
XBUFX2_293 BUFX2_293/A gnd instr2_o[31] vdd BUFX2
XFILL_0_NAND2X1_679 gnd vdd FILL
XFILL_2_DFFPOSX1_184 gnd vdd FILL
XBUFX2_282 INVX1_73/A gnd instr1_o[3] vdd BUFX2
XFILL_5_DFFPOSX1_600 gnd vdd FILL
XFILL_5_DFFPOSX1_611 gnd vdd FILL
XFILL_5_DFFPOSX1_655 gnd vdd FILL
XFILL_5_DFFPOSX1_633 gnd vdd FILL
XFILL_5_DFFPOSX1_622 gnd vdd FILL
XFILL_5_DFFPOSX1_644 gnd vdd FILL
XFILL_5_DFFPOSX1_688 gnd vdd FILL
XFILL_5_DFFPOSX1_677 gnd vdd FILL
XFILL_5_DFFPOSX1_666 gnd vdd FILL
XFILL_5_DFFPOSX1_699 gnd vdd FILL
XFILL_4_DFFPOSX1_212 gnd vdd FILL
XFILL_4_DFFPOSX1_201 gnd vdd FILL
XNAND3X1_1 NOR2X1_7/Y NOR2X1_8/Y AND2X2_1/Y gnd NOR2X1_9/B vdd NAND3X1
XFILL_4_DFFPOSX1_245 gnd vdd FILL
XFILL_4_DFFPOSX1_234 gnd vdd FILL
XFILL_4_DFFPOSX1_223 gnd vdd FILL
XFILL_4_DFFPOSX1_278 gnd vdd FILL
XFILL_4_DFFPOSX1_267 gnd vdd FILL
XFILL_4_DFFPOSX1_256 gnd vdd FILL
XFILL_27_6_1 gnd vdd FILL
XFILL_4_DFFPOSX1_289 gnd vdd FILL
XFILL_2_BUFX4_311 gnd vdd FILL
XFILL_2_6_1 gnd vdd FILL
XFILL_2_CLKBUF1_93 gnd vdd FILL
XFILL_26_1_0 gnd vdd FILL
XFILL_2_CLKBUF1_60 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XFILL_2_CLKBUF1_82 gnd vdd FILL
XFILL_2_CLKBUF1_71 gnd vdd FILL
XFILL_1_BUFX2_102 gnd vdd FILL
XFILL_1_BUFX2_135 gnd vdd FILL
XFILL_1_BUFX2_146 gnd vdd FILL
XFILL_10_5_1 gnd vdd FILL
XOAI21X1_130 BUFX4_6/A BUFX4_370/Y BUFX2_927/A gnd OAI21X1_131/C vdd OAI21X1
XOAI21X1_163 BUFX4_164/Y INVX2_191/Y OAI21X1_163/C gnd OAI21X1_163/Y vdd OAI21X1
XOAI21X1_141 BUFX4_146/Y INVX2_180/Y OAI21X1_141/C gnd OAI21X1_141/Y vdd OAI21X1
XFILL_0_DFFPOSX1_1030 gnd vdd FILL
XFILL_0_BUFX2_906 gnd vdd FILL
XOAI21X1_174 BUFX4_6/Y NAND2X1_7/B BUFX2_952/A gnd OAI21X1_175/C vdd OAI21X1
XOAI21X1_152 BUFX4_4/A OAI21X1_2/A BUFX2_940/A gnd OAI21X1_153/C vdd OAI21X1
XFILL_1_BUFX2_179 gnd vdd FILL
XFILL_0_BUFX2_939 gnd vdd FILL
XOAI21X1_185 BUFX4_149/Y INVX2_202/Y OAI21X1_185/C gnd OAI21X1_185/Y vdd OAI21X1
XINVX1_205 INVX1_205/A gnd INVX1_205/Y vdd INVX1
XINVX1_216 INVX1_216/A gnd INVX1_216/Y vdd INVX1
XFILL_0_BUFX2_928 gnd vdd FILL
XOAI21X1_196 BUFX4_102/Y BUFX4_367/Y BUFX2_964/A gnd OAI21X1_197/C vdd OAI21X1
XFILL_0_BUFX2_917 gnd vdd FILL
XINVX1_227 INVX1_227/A gnd INVX1_227/Y vdd INVX1
XFILL_6_DFFPOSX1_306 gnd vdd FILL
XFILL_6_DFFPOSX1_317 gnd vdd FILL
XFILL_6_DFFPOSX1_328 gnd vdd FILL
XFILL_9_2_0 gnd vdd FILL
XNAND2X1_16 BUFX2_903/A BUFX4_237/Y gnd OAI21X1_16/C vdd NAND2X1
XNAND2X1_38 BUFX2_865/A OAI21X1_8/B gnd OAI21X1_38/C vdd NAND2X1
XNAND2X1_27 BUFX2_852/A BUFX4_208/Y gnd OAI21X1_27/C vdd NAND2X1
XFILL_0_XNOR2X1_12 gnd vdd FILL
XNAND2X1_49 BUFX2_877/A BUFX4_188/Y gnd OAI21X1_49/C vdd NAND2X1
XNAND2X1_180 BUFX2_471/A BUFX4_236/Y gnd OAI21X1_432/C vdd NAND2X1
XFILL_0_XNOR2X1_23 gnd vdd FILL
XNAND2X1_191 BUFX2_476/A BUFX4_214/Y gnd OAI21X1_439/C vdd NAND2X1
XFILL_0_XNOR2X1_45 gnd vdd FILL
XFILL_0_XNOR2X1_34 gnd vdd FILL
XFILL_0_XNOR2X1_56 gnd vdd FILL
XFILL_4_DFFPOSX1_790 gnd vdd FILL
XFILL_18_6_1 gnd vdd FILL
XFILL_0_XNOR2X1_78 gnd vdd FILL
XFILL_0_XNOR2X1_67 gnd vdd FILL
XFILL_0_XNOR2X1_89 gnd vdd FILL
XFILL_17_1_0 gnd vdd FILL
XFILL_0_BUFX4_210 gnd vdd FILL
XOAI21X1_1404 BUFX4_146/Y BUFX4_82/Y BUFX2_254/A gnd OAI21X1_1405/C vdd OAI21X1
XFILL_1_BUFX2_691 gnd vdd FILL
XFILL_0_BUFX4_221 gnd vdd FILL
XFILL_0_BUFX4_232 gnd vdd FILL
XOAI21X1_1415 NAND2X1_625/Y BUFX4_289/Y OAI21X1_1415/C gnd OAI21X1_1415/Y vdd OAI21X1
XFILL_1_OAI21X1_1613 gnd vdd FILL
XOAI21X1_1437 BUFX4_168/Y BUFX4_36/Y BUFX2_203/A gnd OAI21X1_1438/C vdd OAI21X1
XFILL_1_OAI21X1_1602 gnd vdd FILL
XFILL_1_OAI21X1_1624 gnd vdd FILL
XOAI21X1_1426 BUFX4_171/Y BUFX4_52/Y BUFX2_199/A gnd OAI21X1_1427/C vdd OAI21X1
XFILL_0_BUFX4_265 gnd vdd FILL
XFILL_0_BUFX4_243 gnd vdd FILL
XFILL_0_BUFX4_254 gnd vdd FILL
XFILL_0_BUFX4_276 gnd vdd FILL
XFILL_1_OAI21X1_1646 gnd vdd FILL
XOAI21X1_1459 BUFX4_159/Y BUFX4_65/Y BUFX2_212/A gnd OAI21X1_1460/C vdd OAI21X1
XFILL_1_OAI21X1_1635 gnd vdd FILL
XNOR3X1_4 NOR3X1_4/A NOR3X1_4/B NOR3X1_4/C gnd NOR3X1_4/Y vdd NOR3X1
XFILL_0_BUFX4_298 gnd vdd FILL
XFILL_0_BUFX4_287 gnd vdd FILL
XOAI21X1_1448 INVX1_222/A OR2X2_18/B INVX2_70/Y gnd OAI21X1_1449/C vdd OAI21X1
XFILL_3_DFFPOSX1_391 gnd vdd FILL
XFILL_3_DFFPOSX1_380 gnd vdd FILL
XFILL_1_OAI21X1_1657 gnd vdd FILL
XFILL_0_OAI21X1_404 gnd vdd FILL
XFILL_1_OAI21X1_1679 gnd vdd FILL
XFILL_1_OAI21X1_1668 gnd vdd FILL
XFILL_0_OAI21X1_437 gnd vdd FILL
XFILL_1_OAI21X1_608 gnd vdd FILL
XFILL_0_OAI21X1_426 gnd vdd FILL
XFILL_0_OAI21X1_415 gnd vdd FILL
XFILL_0_OAI21X1_459 gnd vdd FILL
XFILL_1_OAI21X1_619 gnd vdd FILL
XFILL_0_OAI21X1_448 gnd vdd FILL
XFILL_3_DFFPOSX1_1012 gnd vdd FILL
XFILL_3_DFFPOSX1_1001 gnd vdd FILL
XFILL_0_INVX4_51 gnd vdd FILL
XFILL_3_DFFPOSX1_1023 gnd vdd FILL
XFILL_0_INVX4_40 gnd vdd FILL
XFILL_6_DFFPOSX1_884 gnd vdd FILL
XFILL_6_DFFPOSX1_895 gnd vdd FILL
XXNOR2X1_91 INVX2_108/A bundleAddress_i[52] gnd XNOR2X1_91/Y vdd XNOR2X1
XXNOR2X1_80 AND2X2_29/A bundleAddress_i[36] gnd XNOR2X1_80/Y vdd XNOR2X1
XFILL_0_NAND2X1_410 gnd vdd FILL
XFILL_1_XNOR2X1_3 gnd vdd FILL
XFILL_0_OAI21X1_1214 gnd vdd FILL
XFILL_0_NAND2X1_432 gnd vdd FILL
XFILL_0_OAI21X1_1203 gnd vdd FILL
XFILL_0_NAND2X1_421 gnd vdd FILL
XFILL_0_NAND2X1_443 gnd vdd FILL
XFILL_0_DFFPOSX1_815 gnd vdd FILL
XFILL_0_OAI21X1_1236 gnd vdd FILL
XFILL_0_OAI21X1_1225 gnd vdd FILL
XFILL_1_NAND2X1_658 gnd vdd FILL
XFILL_0_NAND2X1_487 gnd vdd FILL
XFILL_0_OAI21X1_1247 gnd vdd FILL
XFILL_1_NAND2X1_625 gnd vdd FILL
XFILL_0_NAND2X1_476 gnd vdd FILL
XBUFX2_90 BUFX2_90/A gnd addr2_o[32] vdd BUFX2
XFILL_0_NAND2X1_465 gnd vdd FILL
XFILL_0_DFFPOSX1_804 gnd vdd FILL
XFILL_0_NAND2X1_454 gnd vdd FILL
XFILL_0_OAI21X1_1258 gnd vdd FILL
XFILL_0_DFFPOSX1_837 gnd vdd FILL
XFILL_0_NAND2X1_498 gnd vdd FILL
XFILL_1_NAND2X1_669 gnd vdd FILL
XFILL_0_OAI21X1_1269 gnd vdd FILL
XFILL_0_DFFPOSX1_848 gnd vdd FILL
XFILL_0_DFFPOSX1_826 gnd vdd FILL
XFILL_0_DFFPOSX1_859 gnd vdd FILL
XFILL_5_DFFPOSX1_430 gnd vdd FILL
XFILL_5_DFFPOSX1_463 gnd vdd FILL
XFILL_5_DFFPOSX1_452 gnd vdd FILL
XFILL_5_DFFPOSX1_441 gnd vdd FILL
XFILL_24_15_0 gnd vdd FILL
XFILL_5_DFFPOSX1_485 gnd vdd FILL
XFILL_5_DFFPOSX1_496 gnd vdd FILL
XFILL_5_DFFPOSX1_474 gnd vdd FILL
XFILL_1_BUFX4_90 gnd vdd FILL
XFILL_0_AOI21X1_23 gnd vdd FILL
XFILL_0_AOI21X1_12 gnd vdd FILL
XFILL_0_AOI21X1_45 gnd vdd FILL
XFILL_0_AOI21X1_34 gnd vdd FILL
XFILL_0_AOI21X1_56 gnd vdd FILL
XFILL_2_CLKBUF1_3 gnd vdd FILL
XFILL_0_OAI21X1_960 gnd vdd FILL
XFILL_0_OAI21X1_971 gnd vdd FILL
XFILL_0_OAI21X1_993 gnd vdd FILL
XFILL_0_OAI21X1_982 gnd vdd FILL
XFILL_2_DFFPOSX1_909 gnd vdd FILL
XFILL_2_BUFX4_163 gnd vdd FILL
XFILL_2_MUX2X1_1 gnd vdd FILL
XFILL_6_DFFPOSX1_1027 gnd vdd FILL
XFILL_29_14_0 gnd vdd FILL
XFILL_2_BUFX4_196 gnd vdd FILL
XFILL_0_OAI21X1_1770 gnd vdd FILL
XFILL_0_OAI21X1_1792 gnd vdd FILL
XFILL_0_OAI21X1_1781 gnd vdd FILL
XFILL_0_BUFX2_714 gnd vdd FILL
XFILL_0_NOR2X1_32 gnd vdd FILL
XFILL_0_NOR2X1_21 gnd vdd FILL
XFILL_0_BUFX2_703 gnd vdd FILL
XFILL_0_NOR2X1_10 gnd vdd FILL
XFILL_0_BUFX2_736 gnd vdd FILL
XFILL_0_BUFX2_725 gnd vdd FILL
XFILL_0_BUFX2_747 gnd vdd FILL
XFILL_0_NOR2X1_54 gnd vdd FILL
XFILL_0_NOR2X1_43 gnd vdd FILL
XFILL_0_NOR2X1_76 gnd vdd FILL
XFILL_0_NOR2X1_65 gnd vdd FILL
XFILL_0_BUFX2_758 gnd vdd FILL
XFILL_0_NOR2X1_98 gnd vdd FILL
XFILL_0_NOR2X1_87 gnd vdd FILL
XFILL_0_BUFX2_769 gnd vdd FILL
XFILL_3_DFFPOSX1_9 gnd vdd FILL
XFILL_6_DFFPOSX1_169 gnd vdd FILL
XBUFX4_322 BUFX4_380/A gnd BUFX4_322/Y vdd BUFX4
XBUFX4_311 BUFX4_378/A gnd BUFX4_311/Y vdd BUFX4
XBUFX4_300 BUFX4_303/A gnd BUFX4_300/Y vdd BUFX4
XBUFX4_344 BUFX4_381/A gnd BUFX4_344/Y vdd BUFX4
XBUFX4_333 BUFX4_378/A gnd OAI21X1_2/A vdd BUFX4
XFILL_4_15_0 gnd vdd FILL
XBUFX4_355 BUFX4_388/A gnd BUFX4_355/Y vdd BUFX4
XBUFX4_377 BUFX4_380/A gnd BUFX4_377/Y vdd BUFX4
XBUFX4_366 BUFX4_376/A gnd BUFX4_366/Y vdd BUFX4
XBUFX4_388 BUFX4_388/A gnd BUFX4_388/Y vdd BUFX4
XFILL_33_4_1 gnd vdd FILL
XFILL_19_2 gnd vdd FILL
XFILL_0_NAND2X1_9 gnd vdd FILL
XOAI21X1_1212 BUFX4_94/Y BUFX4_312/Y BUFX2_141/A gnd OAI21X1_1213/C vdd OAI21X1
XOAI21X1_1201 OAI21X1_1201/A AOI21X1_44/Y NAND2X1_584/Y gnd OAI21X1_1201/Y vdd OAI21X1
XOAI21X1_1223 BUFX4_8/A BUFX4_382/Y BUFX2_185/A gnd OAI21X1_1224/C vdd OAI21X1
XDFFPOSX1_813 BUFX2_110/A CLKBUF1_12/Y OAI21X1_1108/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1432 gnd vdd FILL
XOAI21X1_1256 NOR2X1_184/B INVX2_105/Y INVX2_68/Y gnd NAND2X1_597/A vdd OAI21X1
XOAI21X1_1234 BUFX4_2/A BUFX4_382/Y BUFX2_131/A gnd OAI21X1_1235/C vdd OAI21X1
XDFFPOSX1_824 BUFX2_73/A CLKBUF1_23/Y OAI21X1_1130/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1421 gnd vdd FILL
XFILL_1_OAI21X1_1410 gnd vdd FILL
XOAI21X1_1245 OAI21X1_1245/A BUFX4_127/Y OAI21X1_1245/C gnd OAI21X1_1245/Y vdd OAI21X1
XDFFPOSX1_802 BUFX2_55/A CLKBUF1_97/Y OAI21X1_1094/Y gnd vdd DFFPOSX1
XDFFPOSX1_835 BUFX2_85/A CLKBUF1_7/Y OAI21X1_1147/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_201 gnd vdd FILL
XFILL_1_OAI21X1_1465 gnd vdd FILL
XOAI21X1_1289 NAND2X1_606/Y INVX4_38/Y MUX2X1_2/S gnd OAI21X1_1290/A vdd OAI21X1
XFILL_1_OAI21X1_1454 gnd vdd FILL
XOAI21X1_1278 BUFX4_4/A OAI21X1_5/A BUFX2_147/A gnd OAI21X1_1280/C vdd OAI21X1
XFILL_0_OAI21X1_212 gnd vdd FILL
XFILL_1_CLKBUF1_90 gnd vdd FILL
XDFFPOSX1_857 BUFX2_109/A CLKBUF1_36/Y OAI21X1_1179/Y gnd vdd DFFPOSX1
XOAI21X1_1267 OAI21X1_1267/A BUFX4_157/Y OAI21X1_1267/C gnd OAI21X1_1267/Y vdd OAI21X1
XFILL_1_OAI21X1_1443 gnd vdd FILL
XDFFPOSX1_846 BUFX2_97/A CLKBUF1_28/Y OAI21X1_1163/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_234 gnd vdd FILL
XDFFPOSX1_879 BUFX2_190/A CLKBUF1_31/Y OAI21X1_1227/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_223 gnd vdd FILL
XFILL_1_OAI21X1_1476 gnd vdd FILL
XFILL_0_OAI21X1_245 gnd vdd FILL
XDFFPOSX1_868 BUFX2_122/A CLKBUF1_69/Y OAI21X1_1201/Y gnd vdd DFFPOSX1
XINVX2_18 bundleStartMajId_i[45] gnd INVX2_18/Y vdd INVX2
XFILL_1_OAI21X1_427 gnd vdd FILL
XFILL_1_OAI21X1_416 gnd vdd FILL
XFILL_1_OAI21X1_1487 gnd vdd FILL
XFILL_1_OAI21X1_405 gnd vdd FILL
XFILL_1_OAI21X1_1498 gnd vdd FILL
XFILL_0_OAI21X1_289 gnd vdd FILL
XFILL_0_OAI21X1_267 gnd vdd FILL
XFILL_0_OAI21X1_278 gnd vdd FILL
XINVX2_29 bundleStartMajId_i[19] gnd NOR3X1_2/A vdd INVX2
XFILL_1_OAI21X1_438 gnd vdd FILL
XFILL_0_OAI21X1_256 gnd vdd FILL
XFILL_1_OAI21X1_449 gnd vdd FILL
XFILL_9_14_0 gnd vdd FILL
XFILL_6_DFFPOSX1_670 gnd vdd FILL
XFILL_6_DFFPOSX1_681 gnd vdd FILL
XFILL_6_DFFPOSX1_692 gnd vdd FILL
XFILL_13_12_1 gnd vdd FILL
XFILL_1_INVX4_18 gnd vdd FILL
XFILL_1_NAND2X1_411 gnd vdd FILL
XFILL_0_OAI21X1_1022 gnd vdd FILL
XFILL_0_NAND2X1_240 gnd vdd FILL
XFILL_0_NAND2X1_251 gnd vdd FILL
XFILL_1_INVX4_29 gnd vdd FILL
XFILL_1_NAND2X1_400 gnd vdd FILL
XFILL_0_OAI21X1_1000 gnd vdd FILL
XFILL_0_OAI21X1_1011 gnd vdd FILL
XFILL_1_NAND2X1_422 gnd vdd FILL
XFILL_1_NAND2X1_466 gnd vdd FILL
XFILL_0_OAI21X1_1033 gnd vdd FILL
XFILL_1_BUFX4_208 gnd vdd FILL
XFILL_0_OAI21X1_1044 gnd vdd FILL
XFILL_0_OAI21X1_1066 gnd vdd FILL
XFILL_1_BUFX4_219 gnd vdd FILL
XFILL_24_4_1 gnd vdd FILL
XFILL_0_NAND2X1_262 gnd vdd FILL
XFILL_1_NAND2X1_444 gnd vdd FILL
XFILL_0_OAI21X1_1055 gnd vdd FILL
XFILL_0_NAND2X1_284 gnd vdd FILL
XFILL_0_NAND2X1_295 gnd vdd FILL
XFILL_0_DFFPOSX1_601 gnd vdd FILL
XFILL_0_NAND2X1_273 gnd vdd FILL
XFILL_0_DFFPOSX1_612 gnd vdd FILL
XFILL_0_DFFPOSX1_623 gnd vdd FILL
XFILL_0_DFFPOSX1_645 gnd vdd FILL
XFILL_0_DFFPOSX1_634 gnd vdd FILL
XFILL_0_DFFPOSX1_656 gnd vdd FILL
XFILL_1_NAND2X1_488 gnd vdd FILL
XFILL_1_NAND2X1_477 gnd vdd FILL
XFILL_1_NAND2X1_499 gnd vdd FILL
XFILL_0_OAI21X1_1099 gnd vdd FILL
XFILL_0_OAI21X1_1088 gnd vdd FILL
XFILL_0_DFFPOSX1_667 gnd vdd FILL
XFILL_0_OAI21X1_1077 gnd vdd FILL
XFILL_0_DFFPOSX1_678 gnd vdd FILL
XFILL_0_DFFPOSX1_689 gnd vdd FILL
XFILL_5_DFFPOSX1_271 gnd vdd FILL
XFILL_5_DFFPOSX1_260 gnd vdd FILL
XFILL_5_DFFPOSX1_282 gnd vdd FILL
XFILL_5_DFFPOSX1_293 gnd vdd FILL
XOAI21X1_1790 BUFX4_334/Y INVX2_162/Y NAND2X1_731/Y gnd OAI21X1_1790/Y vdd OAI21X1
XFILL_1_OAI21X1_950 gnd vdd FILL
XFILL_2_BUFX4_46 gnd vdd FILL
XFILL_18_11_1 gnd vdd FILL
XFILL_2_BUFX4_79 gnd vdd FILL
XFILL_0_OAI21X1_790 gnd vdd FILL
XFILL_1_OR2X2_2 gnd vdd FILL
XFILL_1_OAI21X1_961 gnd vdd FILL
XFILL_1_OAI21X1_972 gnd vdd FILL
XFILL_7_5_1 gnd vdd FILL
XFILL_1_OAI21X1_983 gnd vdd FILL
XFILL_1_OAI21X1_994 gnd vdd FILL
XFILL_6_0_0 gnd vdd FILL
XBUFX2_804 BUFX2_804/A gnd tid1_o[30] vdd BUFX2
XFILL_31_13_1 gnd vdd FILL
XFILL_2_OAI21X1_1138 gnd vdd FILL
XBUFX2_826 BUFX2_826/A gnd tid1_o[10] vdd BUFX2
XBUFX2_815 BUFX2_815/A gnd tid1_o[20] vdd BUFX2
XFILL_2_DFFPOSX1_728 gnd vdd FILL
XFILL_2_DFFPOSX1_706 gnd vdd FILL
XFILL_2_DFFPOSX1_717 gnd vdd FILL
XFILL_2_DFFPOSX1_739 gnd vdd FILL
XBUFX2_837 NAND2X1_7/A gnd tid1_o[0] vdd BUFX2
XBUFX2_848 BUFX2_848/A gnd tid2_o[48] vdd BUFX2
XBUFX2_859 BUFX2_859/A gnd tid2_o[38] vdd BUFX2
XFILL_15_4_1 gnd vdd FILL
XMUX2X1_2 MUX2X1_2/A MUX2X1_2/B MUX2X1_2/S gnd MUX2X1_2/Y vdd MUX2X1
XFILL_2_OR2X2_16 gnd vdd FILL
XFILL_0_BUFX2_511 gnd vdd FILL
XFILL_0_BUFX2_500 gnd vdd FILL
XDFFPOSX1_109 BUFX2_840/A CLKBUF1_1/Y OAI21X1_1783/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_533 gnd vdd FILL
XFILL_0_BUFX2_522 gnd vdd FILL
XFILL_1_DFFPOSX1_318 gnd vdd FILL
XFILL_1_DFFPOSX1_307 gnd vdd FILL
XFILL_1_DFFPOSX1_329 gnd vdd FILL
XCLKBUF1_3 BUFX4_86/Y gnd CLKBUF1_3/Y vdd CLKBUF1
XFILL_0_BUFX2_555 gnd vdd FILL
XFILL_0_BUFX2_544 gnd vdd FILL
XFILL_0_BUFX2_566 gnd vdd FILL
XFILL_0_BUFX2_588 gnd vdd FILL
XFILL_0_BUFX2_599 gnd vdd FILL
XFILL_0_BUFX2_577 gnd vdd FILL
XFILL_36_12_1 gnd vdd FILL
XBUFX4_130 BUFX4_19/Y gnd BUFX4_130/Y vdd BUFX4
XFILL_4_CLKBUF1_12 gnd vdd FILL
XFILL_0_INVX1_41 gnd vdd FILL
XBUFX4_141 BUFX4_16/Y gnd BUFX4_141/Y vdd BUFX4
XFILL_0_INVX1_30 gnd vdd FILL
XFILL_4_CLKBUF1_34 gnd vdd FILL
XFILL_0_INVX1_52 gnd vdd FILL
XBUFX4_152 BUFX4_16/Y gnd BUFX4_152/Y vdd BUFX4
XBUFX4_163 BUFX4_13/Y gnd BUFX4_163/Y vdd BUFX4
XFILL_0_INVX1_85 gnd vdd FILL
XFILL_0_INVX1_74 gnd vdd FILL
XFILL_0_INVX1_63 gnd vdd FILL
XFILL_4_CLKBUF1_67 gnd vdd FILL
XNOR2X1_223 INVX1_202/A NOR2X1_223/B gnd XNOR2X1_96/A vdd NOR2X1
XFILL_4_CLKBUF1_45 gnd vdd FILL
XBUFX4_174 BUFX4_15/Y gnd BUFX4_174/Y vdd BUFX4
XNOR2X1_212 bundleAddress_i[2] INVX1_217/Y gnd NOR2X1_212/Y vdd NOR2X1
XNOR2X1_201 NOR3X1_16/B NOR2X1_201/B gnd NOR2X1_201/Y vdd NOR2X1
XBUFX4_185 BUFX4_21/Y gnd OAI21X1_9/B vdd BUFX4
XBUFX4_196 BUFX4_21/Y gnd BUFX4_196/Y vdd BUFX4
XFILL_31_1 gnd vdd FILL
XFILL_0_BUFX2_27 gnd vdd FILL
XFILL_4_CLKBUF1_89 gnd vdd FILL
XFILL_4_CLKBUF1_78 gnd vdd FILL
XFILL_0_INVX1_96 gnd vdd FILL
XFILL_0_BUFX2_16 gnd vdd FILL
XFILL_0_BUFX2_38 gnd vdd FILL
XFILL_0_BUFX2_49 gnd vdd FILL
XOAI21X1_718 INVX1_37/Y OAI21X1_718/B OAI21X1_718/C gnd OAI21X1_718/Y vdd OAI21X1
XOAI21X1_707 BUFX4_175/Y BUFX4_56/Y BUFX2_594/A gnd OAI21X1_708/C vdd OAI21X1
XOAI21X1_729 OAI21X1_729/A BUFX4_295/Y OAI21X1_729/C gnd OAI21X1_729/Y vdd OAI21X1
XOAI21X1_1031 BUFX4_293/Y INVX1_170/Y OAI21X1_1031/C gnd OAI21X1_1031/Y vdd OAI21X1
XOAI21X1_1020 BUFX4_136/Y BUFX4_81/Y BUFX2_374/A gnd OAI21X1_1021/C vdd OAI21X1
XFILL_1_OAI21X1_1240 gnd vdd FILL
XOAI21X1_1053 BUFX4_385/Y INVX2_68/Y NAND2X1_419/Y gnd OAI21X1_1053/Y vdd OAI21X1
XOAI21X1_1042 BUFX4_347/Y INVX2_59/Y NAND2X1_408/Y gnd OAI21X1_1042/Y vdd OAI21X1
XDFFPOSX1_632 INVX1_61/A CLKBUF1_61/Y OAI21X1_860/Y gnd vdd DFFPOSX1
XOAI21X1_1064 BUFX4_317/Y INVX1_176/Y NAND2X1_430/Y gnd OAI21X1_1064/Y vdd OAI21X1
XDFFPOSX1_621 INVX1_50/A CLKBUF1_78/Y OAI21X1_849/Y gnd vdd DFFPOSX1
XDFFPOSX1_610 BUFX2_644/A CLKBUF1_29/Y OAI21X1_840/Y gnd vdd DFFPOSX1
XDFFPOSX1_654 BUFX2_321/A CLKBUF1_32/Y OAI21X1_882/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1251 gnd vdd FILL
XFILL_1_DFFPOSX1_841 gnd vdd FILL
XFILL_1_OAI21X1_1284 gnd vdd FILL
XFILL_1_OAI21X1_1262 gnd vdd FILL
XFILL_1_OAI21X1_1273 gnd vdd FILL
XOAI21X1_1097 BUFX4_357/Y INVX2_91/Y NAND2X1_463/Y gnd OAI21X1_1097/Y vdd OAI21X1
XDFFPOSX1_643 INVX1_72/A CLKBUF1_71/Y OAI21X1_871/Y gnd vdd DFFPOSX1
XDFFPOSX1_665 BUFX2_302/A CLKBUF1_75/Y OAI21X1_893/Y gnd vdd DFFPOSX1
XOAI21X1_1075 BUFX4_350/Y INVX8_3/Y NAND2X1_441/Y gnd OAI21X1_1075/Y vdd OAI21X1
XFILL_1_DFFPOSX1_830 gnd vdd FILL
XOAI21X1_1086 BUFX4_364/Y INVX4_44/Y NAND2X1_452/Y gnd OAI21X1_1086/Y vdd OAI21X1
XFILL_1_DFFPOSX1_874 gnd vdd FILL
XFILL_1_OAI21X1_224 gnd vdd FILL
XFILL_1_OAI21X1_235 gnd vdd FILL
XDFFPOSX1_698 BUFX2_335/A CLKBUF1_96/Y OAI21X1_945/Y gnd vdd DFFPOSX1
XNAND2X1_702 BUFX2_694/A BUFX4_195/Y gnd NAND2X1_702/Y vdd NAND2X1
XFILL_1_OAI21X1_1295 gnd vdd FILL
XFILL_1_DFFPOSX1_885 gnd vdd FILL
XFILL_1_DFFPOSX1_852 gnd vdd FILL
XDFFPOSX1_687 BUFX2_354/A CLKBUF1_40/Y OAI21X1_923/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_213 gnd vdd FILL
XDFFPOSX1_676 BUFX2_314/A CLKBUF1_53/Y OAI21X1_904/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_863 gnd vdd FILL
XFILL_1_OAI21X1_202 gnd vdd FILL
XFILL_1_OAI21X1_268 gnd vdd FILL
XFILL_1_OAI21X1_246 gnd vdd FILL
XNAND2X1_746 BUFX2_802/A BUFX4_366/Y gnd NAND2X1_746/Y vdd NAND2X1
XNAND2X1_724 BUFX2_840/A BUFX4_378/Y gnd NAND2X1_724/Y vdd NAND2X1
XFILL_1_DFFPOSX1_896 gnd vdd FILL
XNAND2X1_735 BUFX2_790/A BUFX4_383/Y gnd NAND2X1_735/Y vdd NAND2X1
XFILL_1_OAI21X1_257 gnd vdd FILL
XFILL_0_NOR2X1_7 gnd vdd FILL
XNAND2X1_713 BUFX2_706/A BUFX4_217/Y gnd NAND2X1_713/Y vdd NAND2X1
XNAND2X1_768 BUFX2_826/A BUFX4_380/Y gnd NAND2X1_768/Y vdd NAND2X1
XFILL_1_OAI21X1_279 gnd vdd FILL
XNAND2X1_757 BUFX2_814/A BUFX4_384/Y gnd NAND2X1_757/Y vdd NAND2X1
XFILL_2_XNOR2X1_19 gnd vdd FILL
XFILL_1_NAND2X1_252 gnd vdd FILL
XFILL_1_NAND2X1_274 gnd vdd FILL
XFILL_0_DFFPOSX1_431 gnd vdd FILL
XFILL_0_DFFPOSX1_420 gnd vdd FILL
XFILL_0_DFFPOSX1_442 gnd vdd FILL
XFILL_2_DFFPOSX1_6 gnd vdd FILL
XFILL_0_DFFPOSX1_453 gnd vdd FILL
XFILL_0_DFFPOSX1_464 gnd vdd FILL
XFILL_0_DFFPOSX1_475 gnd vdd FILL
XINVX8_5 bundleLen_i[0] gnd INVX8_5/Y vdd INVX8
XFILL_0_DFFPOSX1_486 gnd vdd FILL
XFILL_0_DFFPOSX1_497 gnd vdd FILL
XFILL_3_DFFPOSX1_902 gnd vdd FILL
XFILL_3_DFFPOSX1_913 gnd vdd FILL
XFILL_3_DFFPOSX1_946 gnd vdd FILL
XFILL_3_DFFPOSX1_935 gnd vdd FILL
XFILL_3_DFFPOSX1_924 gnd vdd FILL
XFILL_3_DFFPOSX1_957 gnd vdd FILL
XFILL_3_DFFPOSX1_968 gnd vdd FILL
XFILL_3_DFFPOSX1_979 gnd vdd FILL
XDFFPOSX1_80 BUFX2_749/A CLKBUF1_45/Y DFFPOSX1_80/D gnd vdd DFFPOSX1
XDFFPOSX1_91 BUFX2_761/A CLKBUF1_32/Y DFFPOSX1_91/D gnd vdd DFFPOSX1
XBUFX4_14 INVX8_6/Y gnd BUFX4_14/Y vdd BUFX4
XBUFX4_25 BUFX4_26/A gnd BUFX4_25/Y vdd BUFX4
XFILL_1_OAI21X1_780 gnd vdd FILL
XFILL_1_OAI21X1_791 gnd vdd FILL
XBUFX4_36 BUFX4_67/A gnd BUFX4_36/Y vdd BUFX4
XBUFX4_47 BUFX4_51/A gnd BUFX4_47/Y vdd BUFX4
XBUFX4_69 BUFX4_72/A gnd BUFX4_69/Y vdd BUFX4
XBUFX4_58 BUFX4_73/A gnd BUFX4_58/Y vdd BUFX4
XFILL_2_DFFPOSX1_503 gnd vdd FILL
XFILL_2_DFFPOSX1_514 gnd vdd FILL
XBUFX2_612 BUFX2_612/A gnd majID4_o[30] vdd BUFX2
XBUFX2_601 BUFX2_601/A gnd majID4_o[40] vdd BUFX2
XBUFX2_623 BUFX2_623/A gnd majID4_o[20] vdd BUFX2
XFILL_2_DFFPOSX1_547 gnd vdd FILL
XFILL_2_DFFPOSX1_525 gnd vdd FILL
XFILL_2_DFFPOSX1_536 gnd vdd FILL
XBUFX2_634 BUFX2_634/A gnd majID4_o[10] vdd BUFX2
XBUFX2_645 BUFX2_645/A gnd majID4_o[0] vdd BUFX2
XBUFX2_656 BUFX2_656/A gnd pid1_o[16] vdd BUFX2
XBUFX2_678 BUFX2_678/A gnd pid1_o[24] vdd BUFX2
XFILL_2_DFFPOSX1_569 gnd vdd FILL
XBUFX2_667 BUFX2_667/A gnd pid1_o[6] vdd BUFX2
XFILL_2_DFFPOSX1_558 gnd vdd FILL
XBUFX2_689 BUFX2_689/A gnd pid2_o[15] vdd BUFX2
XFILL_30_2_1 gnd vdd FILL
XFILL_22_18_1 gnd vdd FILL
XINVX2_130 bundlePid_i[18] gnd INVX2_130/Y vdd INVX2
XFILL_1_DFFPOSX1_104 gnd vdd FILL
XOR2X2_17 OR2X2_18/A OR2X2_17/B gnd OR2X2_17/Y vdd OR2X2
XFILL_0_BUFX2_330 gnd vdd FILL
XFILL_0_BUFX2_341 gnd vdd FILL
XINVX2_141 bundlePid_i[7] gnd INVX2_141/Y vdd INVX2
XINVX2_163 bundleTid_i[46] gnd INVX2_163/Y vdd INVX2
XFILL_1_DFFPOSX1_126 gnd vdd FILL
XFILL_1_DFFPOSX1_115 gnd vdd FILL
XINVX2_152 bundleTid_i[57] gnd INVX2_152/Y vdd INVX2
XFILL_1_DFFPOSX1_137 gnd vdd FILL
XFILL_0_BUFX2_374 gnd vdd FILL
XINVX2_174 bundleTid_i[35] gnd INVX2_174/Y vdd INVX2
XFILL_0_BUFX2_363 gnd vdd FILL
XFILL_0_BUFX2_352 gnd vdd FILL
XINVX2_196 bundleTid_i[13] gnd INVX2_196/Y vdd INVX2
XFILL_0_BUFX2_385 gnd vdd FILL
XFILL_1_DFFPOSX1_148 gnd vdd FILL
XINVX2_185 bundleTid_i[24] gnd INVX2_185/Y vdd INVX2
XFILL_0_BUFX2_396 gnd vdd FILL
XFILL_1_DFFPOSX1_159 gnd vdd FILL
XFILL_4_DFFPOSX1_608 gnd vdd FILL
XFILL_4_DFFPOSX1_619 gnd vdd FILL
XFILL_38_3_1 gnd vdd FILL
XFILL_1_BUFX2_509 gnd vdd FILL
XFILL_27_17_1 gnd vdd FILL
XFILL_21_2_1 gnd vdd FILL
XOAI21X1_504 BUFX4_7/Y BUFX4_365/Y BUFX2_533/A gnd OAI21X1_505/C vdd OAI21X1
XFILL_3_DFFPOSX1_209 gnd vdd FILL
XOAI21X1_526 XNOR2X1_25/Y BUFX4_161/Y OAI21X1_526/C gnd OAI21X1_526/Y vdd OAI21X1
XOAI21X1_548 XNOR2X1_28/Y BUFX4_135/Y OAI21X1_548/C gnd OAI21X1_548/Y vdd OAI21X1
XOAI21X1_537 BUFX4_101/Y BUFX4_358/Y BUFX2_526/A gnd OAI21X1_538/C vdd OAI21X1
XOAI21X1_515 INVX4_29/A OAI21X1_515/B OAI21X1_515/C gnd OAI21X1_515/Y vdd OAI21X1
XOAI21X1_559 NOR2X1_64/Y NOR2X1_65/B OAI21X1_559/C gnd OAI21X1_559/Y vdd OAI21X1
XFILL_21_13_0 gnd vdd FILL
XDFFPOSX1_440 BUFX2_470/A CLKBUF1_18/Y OAI21X1_431/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_660 gnd vdd FILL
XFILL_1_OAI21X1_1081 gnd vdd FILL
XFILL_1_OAI21X1_1070 gnd vdd FILL
XDFFPOSX1_462 BUFX2_494/A CLKBUF1_90/Y OAI21X1_463/Y gnd vdd DFFPOSX1
XDFFPOSX1_451 INVX1_14/A CLKBUF1_63/Y OAI21X1_447/Y gnd vdd DFFPOSX1
XDFFPOSX1_473 BUFX2_506/A CLKBUF1_6/Y OAI21X1_481/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1092 gnd vdd FILL
XNAND2X1_521 BUFX2_84/A BUFX4_229/Y gnd NAND2X1_521/Y vdd NAND2X1
XFILL_2_OAI21X1_214 gnd vdd FILL
XDFFPOSX1_484 BUFX2_521/A CLKBUF1_45/Y OAI21X1_501/Y gnd vdd DFFPOSX1
XDFFPOSX1_495 BUFX2_524/A CLKBUF1_90/Y OAI21X1_534/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_693 gnd vdd FILL
XFILL_1_DFFPOSX1_671 gnd vdd FILL
XFILL_1_DFFPOSX1_682 gnd vdd FILL
XNAND2X1_510 BUFX2_80/A BUFX4_186/Y gnd NAND2X1_510/Y vdd NAND2X1
XNAND2X1_532 BUFX2_92/A BUFX4_202/Y gnd NAND2X1_532/Y vdd NAND2X1
XNAND2X1_554 BUFX4_238/Y NAND2X1_554/B gnd NAND2X1_554/Y vdd NAND2X1
XNAND2X1_543 BUFX2_97/A BUFX4_226/Y gnd NAND2X1_543/Y vdd NAND2X1
XNAND2X1_587 BUFX2_124/A BUFX4_187/Y gnd NAND2X1_587/Y vdd NAND2X1
XNAND2X1_565 AND2X2_24/B AND2X2_24/A gnd NOR3X1_14/C vdd NAND2X1
XFILL_1_OAI22X1_1 gnd vdd FILL
XNAND2X1_576 BUFX2_115/A BUFX4_201/Y gnd NAND2X1_576/Y vdd NAND2X1
XFILL_29_3_1 gnd vdd FILL
XNAND2X1_598 INVX1_201/Y AND2X2_26/A gnd NOR3X1_18/C vdd NAND2X1
XFILL_4_3_1 gnd vdd FILL
XFILL_2_18_1 gnd vdd FILL
XFILL_0_AND2X2_33 gnd vdd FILL
XFILL_0_AND2X2_22 gnd vdd FILL
XFILL_0_AND2X2_11 gnd vdd FILL
XFILL_0_DFFPOSX1_250 gnd vdd FILL
XFILL_0_DFFPOSX1_261 gnd vdd FILL
XFILL_0_DFFPOSX1_272 gnd vdd FILL
XFILL_26_12_0 gnd vdd FILL
XFILL_0_DFFPOSX1_283 gnd vdd FILL
XFILL_12_2_1 gnd vdd FILL
XFILL_0_DFFPOSX1_294 gnd vdd FILL
XFILL_3_DFFPOSX1_710 gnd vdd FILL
XFILL_3_DFFPOSX1_721 gnd vdd FILL
XFILL_3_DFFPOSX1_732 gnd vdd FILL
XFILL_3_DFFPOSX1_754 gnd vdd FILL
XFILL_3_CLKBUF1_42 gnd vdd FILL
XFILL_3_CLKBUF1_31 gnd vdd FILL
XFILL_3_DFFPOSX1_743 gnd vdd FILL
XFILL_3_CLKBUF1_20 gnd vdd FILL
XFILL_3_DFFPOSX1_765 gnd vdd FILL
XFILL_3_DFFPOSX1_776 gnd vdd FILL
XFILL_3_CLKBUF1_64 gnd vdd FILL
XFILL_3_DFFPOSX1_787 gnd vdd FILL
XFILL_3_DFFPOSX1_798 gnd vdd FILL
XFILL_3_CLKBUF1_75 gnd vdd FILL
XFILL_3_CLKBUF1_53 gnd vdd FILL
XFILL_3_CLKBUF1_86 gnd vdd FILL
XFILL_3_CLKBUF1_97 gnd vdd FILL
XFILL_1_NOR2X1_182 gnd vdd FILL
XFILL_1_NOR2X1_193 gnd vdd FILL
XFILL_1_NOR2X1_160 gnd vdd FILL
XFILL_2_NAND3X1_2 gnd vdd FILL
XFILL_7_17_1 gnd vdd FILL
XFILL_2_OAI21X1_792 gnd vdd FILL
XFILL_2_DFFPOSX1_322 gnd vdd FILL
XFILL_2_DFFPOSX1_311 gnd vdd FILL
XFILL_2_DFFPOSX1_300 gnd vdd FILL
XBUFX2_420 BUFX2_420/A gnd majID1_o[30] vdd BUFX2
XFILL_2_DFFPOSX1_333 gnd vdd FILL
XBUFX2_431 BUFX2_431/A gnd majID1_o[20] vdd BUFX2
XBUFX2_442 BUFX2_442/A gnd majID1_o[10] vdd BUFX2
XBUFX2_453 BUFX2_453/A gnd majID1_o[0] vdd BUFX2
XFILL_1_13_0 gnd vdd FILL
XFILL_2_DFFPOSX1_355 gnd vdd FILL
XFILL_2_DFFPOSX1_344 gnd vdd FILL
XBUFX2_475 BUFX2_475/A gnd majID2_o[38] vdd BUFX2
XFILL_2_DFFPOSX1_388 gnd vdd FILL
XBUFX2_486 BUFX2_486/A gnd majID2_o[28] vdd BUFX2
XBUFX2_497 BUFX2_497/A gnd majID2_o[18] vdd BUFX2
XBUFX2_464 BUFX2_464/A gnd majID2_o[48] vdd BUFX2
XFILL_2_DFFPOSX1_377 gnd vdd FILL
XFILL_2_DFFPOSX1_366 gnd vdd FILL
XFILL_2_DFFPOSX1_399 gnd vdd FILL
XFILL_5_DFFPOSX1_804 gnd vdd FILL
XFILL_5_DFFPOSX1_815 gnd vdd FILL
XFILL_5_DFFPOSX1_837 gnd vdd FILL
XFILL_5_DFFPOSX1_826 gnd vdd FILL
XFILL_1_BUFX4_380 gnd vdd FILL
XFILL_5_DFFPOSX1_848 gnd vdd FILL
XFILL_5_DFFPOSX1_859 gnd vdd FILL
XFILL_1_XNOR2X1_16 gnd vdd FILL
XFILL_1_XNOR2X1_27 gnd vdd FILL
XFILL_1_XNOR2X1_38 gnd vdd FILL
XFILL_1_XNOR2X1_49 gnd vdd FILL
XFILL_2_OAI21X1_71 gnd vdd FILL
XFILL_0_BUFX2_171 gnd vdd FILL
XFILL_0_BUFX2_182 gnd vdd FILL
XFILL_0_BUFX2_160 gnd vdd FILL
XFILL_0_BUFX2_193 gnd vdd FILL
XFILL_1_DFFPOSX1_3 gnd vdd FILL
XFILL_4_DFFPOSX1_416 gnd vdd FILL
XFILL_4_DFFPOSX1_405 gnd vdd FILL
XFILL_4_DFFPOSX1_427 gnd vdd FILL
XFILL_4_DFFPOSX1_449 gnd vdd FILL
XFILL_6_12_0 gnd vdd FILL
XFILL_4_DFFPOSX1_438 gnd vdd FILL
XFILL_10_10_1 gnd vdd FILL
XFILL_1_BUFX2_317 gnd vdd FILL
XOAI21X1_301 INVX2_196/Y BUFX4_293/Y OAI21X1_301/C gnd OAI21X1_301/Y vdd OAI21X1
XOAI21X1_312 BUFX4_168/Y BUFX4_36/Y BUFX2_1021/A gnd OAI21X1_313/C vdd OAI21X1
XFILL_1_BUFX2_328 gnd vdd FILL
XOAI21X1_323 INVX2_5/Y BUFX4_290/Y OAI21X1_323/C gnd OAI21X1_323/Y vdd OAI21X1
XOAI21X1_345 BUFX4_387/Y INVX4_7/Y NAND2X1_89/Y gnd OAI21X1_345/Y vdd OAI21X1
XOAI21X1_356 OAI21X1_2/A INVX4_13/Y OAI21X1_356/C gnd OAI21X1_356/Y vdd OAI21X1
XOAI21X1_334 BUFX4_355/Y INVX4_2/Y NAND2X1_78/Y gnd OAI21X1_334/Y vdd OAI21X1
XOAI21X1_378 BUFX4_323/Y INVX2_33/Y OAI21X1_378/C gnd OAI21X1_378/Y vdd OAI21X1
XOAI21X1_367 BUFX4_346/Y INVX4_18/Y OAI21X1_367/C gnd OAI21X1_367/Y vdd OAI21X1
XOAI21X1_389 BUFX4_373/Y INVX4_27/Y OAI21X1_389/C gnd OAI21X1_389/Y vdd OAI21X1
XDFFPOSX1_281 BUFX2_954/A CLKBUF1_95/Y OAI21X1_179/Y gnd vdd DFFPOSX1
XDFFPOSX1_270 BUFX2_942/A CLKBUF1_2/Y OAI21X1_157/Y gnd vdd DFFPOSX1
XDFFPOSX1_292 BUFX2_969/A CLKBUF1_23/Y OAI21X1_201/Y gnd vdd DFFPOSX1
XFILL_3_NOR3X1_12 gnd vdd FILL
XFILL_1_DFFPOSX1_490 gnd vdd FILL
XNAND2X1_362 BUFX4_267/Y bundle_i[7] gnd OAI21X1_868/C vdd NAND2X1
XNAND2X1_340 BUFX4_267/Y bundle_i[29] gnd OAI21X1_846/C vdd NAND2X1
XNAND2X1_351 BUFX4_261/Y bundle_i[18] gnd OAI21X1_857/C vdd NAND2X1
XNAND2X1_384 BUFX2_299/A BUFX4_197/Y gnd OAI21X1_890/C vdd NAND2X1
XNAND2X1_373 BUFX2_316/A BUFX4_205/Y gnd OAI21X1_879/C vdd NAND2X1
XFILL_4_DFFPOSX1_950 gnd vdd FILL
XNAND2X1_395 BUFX2_311/A BUFX4_196/Y gnd OAI21X1_901/C vdd NAND2X1
XFILL_4_DFFPOSX1_961 gnd vdd FILL
XFILL_4_DFFPOSX1_983 gnd vdd FILL
XFILL_4_DFFPOSX1_972 gnd vdd FILL
XFILL_0_INVX1_127 gnd vdd FILL
XFILL_4_DFFPOSX1_994 gnd vdd FILL
XFILL_0_INVX1_116 gnd vdd FILL
XFILL_12_18_0 gnd vdd FILL
XFILL_0_INVX1_105 gnd vdd FILL
XFILL_1_AOI21X1_38 gnd vdd FILL
XFILL_1_AOI21X1_27 gnd vdd FILL
XFILL_1_AOI21X1_49 gnd vdd FILL
XFILL_1_AOI21X1_16 gnd vdd FILL
XFILL_0_INVX1_149 gnd vdd FILL
XFILL_0_INVX1_138 gnd vdd FILL
XFILL_1_BUFX2_840 gnd vdd FILL
XFILL_1_BUFX2_873 gnd vdd FILL
XFILL_1_BUFX2_851 gnd vdd FILL
XFILL_1_BUFX2_884 gnd vdd FILL
XOAI21X1_1608 OAI21X1_1/A INVX2_144/Y NAND2X1_677/Y gnd OAI21X1_1608/Y vdd OAI21X1
XFILL_2_NOR3X1_4 gnd vdd FILL
XFILL_3_DFFPOSX1_540 gnd vdd FILL
XFILL_1_BUFX2_895 gnd vdd FILL
XOAI21X1_1619 INVX2_122/Y BUFX4_206/Y NAND2X1_687/Y gnd DFFPOSX1_9/D vdd OAI21X1
XFILL_1_OAI21X1_1806 gnd vdd FILL
XOAI21X1_890 INVX1_91/Y BUFX4_208/Y OAI21X1_890/C gnd OAI21X1_890/Y vdd OAI21X1
XFILL_1_OAI21X1_1828 gnd vdd FILL
XFILL_1_OAI21X1_1817 gnd vdd FILL
XFILL_3_DFFPOSX1_551 gnd vdd FILL
XFILL_3_DFFPOSX1_573 gnd vdd FILL
XFILL_3_DFFPOSX1_562 gnd vdd FILL
XFILL_3_DFFPOSX1_595 gnd vdd FILL
XFILL_0_OAI21X1_608 gnd vdd FILL
XFILL_3_DFFPOSX1_584 gnd vdd FILL
XFILL_0_OAI21X1_619 gnd vdd FILL
XFILL_7_2 gnd vdd FILL
XFILL_17_17_0 gnd vdd FILL
XFILL_33_10_1 gnd vdd FILL
XFILL_2_DFFPOSX1_130 gnd vdd FILL
XFILL_0_NAND2X1_625 gnd vdd FILL
XFILL_0_NAND2X1_636 gnd vdd FILL
XFILL_0_NAND2X1_603 gnd vdd FILL
XFILL_0_NAND2X1_614 gnd vdd FILL
XFILL_35_1_1 gnd vdd FILL
XFILL_0_NAND2X1_658 gnd vdd FILL
XFILL_0_OAI21X1_1418 gnd vdd FILL
XFILL_0_OAI21X1_1407 gnd vdd FILL
XFILL_0_OAI21X1_1429 gnd vdd FILL
XFILL_0_NAND2X1_647 gnd vdd FILL
XFILL_0_NAND2X1_669 gnd vdd FILL
XBUFX2_250 BUFX2_250/A gnd addr4_o[3] vdd BUFX2
XFILL_2_DFFPOSX1_163 gnd vdd FILL
XBUFX2_272 INVX1_64/A gnd instr1_o[12] vdd BUFX2
XBUFX2_261 INVX1_45/A gnd instr1_o[31] vdd BUFX2
XFILL_2_DFFPOSX1_152 gnd vdd FILL
XFILL_2_DFFPOSX1_141 gnd vdd FILL
XBUFX2_283 INVX1_74/A gnd instr1_o[2] vdd BUFX2
XBUFX2_294 BUFX2_294/A gnd instr2_o[30] vdd BUFX2
XFILL_2_DFFPOSX1_185 gnd vdd FILL
XFILL_2_DFFPOSX1_196 gnd vdd FILL
XFILL_2_DFFPOSX1_174 gnd vdd FILL
XFILL_5_DFFPOSX1_601 gnd vdd FILL
XFILL_5_DFFPOSX1_612 gnd vdd FILL
XFILL_5_DFFPOSX1_645 gnd vdd FILL
XFILL_5_DFFPOSX1_634 gnd vdd FILL
XFILL_5_DFFPOSX1_623 gnd vdd FILL
XFILL_5_DFFPOSX1_656 gnd vdd FILL
XFILL_5_DFFPOSX1_678 gnd vdd FILL
XFILL_5_DFFPOSX1_667 gnd vdd FILL
XFILL_5_DFFPOSX1_689 gnd vdd FILL
XFILL_35_18_0 gnd vdd FILL
XFILL_4_DFFPOSX1_202 gnd vdd FILL
XNAND3X1_2 bundleStartMajId_i[37] INVX1_12/A INVX1_11/Y gnd NAND3X1_2/Y vdd NAND3X1
XFILL_4_DFFPOSX1_213 gnd vdd FILL
XFILL_4_DFFPOSX1_235 gnd vdd FILL
XFILL_4_DFFPOSX1_224 gnd vdd FILL
XFILL_4_DFFPOSX1_246 gnd vdd FILL
XFILL_4_DFFPOSX1_279 gnd vdd FILL
XFILL_4_DFFPOSX1_268 gnd vdd FILL
XFILL_4_DFFPOSX1_257 gnd vdd FILL
XFILL_2_CLKBUF1_50 gnd vdd FILL
XFILL_2_BUFX4_356 gnd vdd FILL
XFILL_26_1_1 gnd vdd FILL
XFILL_2_CLKBUF1_61 gnd vdd FILL
XFILL_2_CLKBUF1_72 gnd vdd FILL
XFILL_2_CLKBUF1_83 gnd vdd FILL
XFILL_1_1_1 gnd vdd FILL
XFILL_2_CLKBUF1_94 gnd vdd FILL
XFILL_1_BUFX2_125 gnd vdd FILL
XFILL_1_BUFX2_114 gnd vdd FILL
XFILL_1_BUFX2_136 gnd vdd FILL
XOAI21X1_120 BUFX4_248/Y BUFX4_361/Y BUFX2_922/A gnd OAI21X1_121/C vdd OAI21X1
XFILL_0_NOR2X1_190 gnd vdd FILL
XFILL_1_BUFX2_169 gnd vdd FILL
XFILL_1_BUFX2_158 gnd vdd FILL
XOAI21X1_131 BUFX4_152/Y INVX2_175/Y OAI21X1_131/C gnd OAI21X1_131/Y vdd OAI21X1
XFILL_0_DFFPOSX1_1020 gnd vdd FILL
XFILL_0_BUFX2_907 gnd vdd FILL
XOAI21X1_142 BUFX4_9/Y BUFX4_376/Y BUFX2_934/A gnd OAI21X1_143/C vdd OAI21X1
XOAI21X1_164 BUFX4_107/Y BUFX4_367/Y BUFX2_946/A gnd OAI21X1_165/C vdd OAI21X1
XOAI21X1_153 BUFX4_133/Y INVX2_186/Y OAI21X1_153/C gnd OAI21X1_153/Y vdd OAI21X1
XFILL_0_BUFX2_929 gnd vdd FILL
XOAI21X1_186 BUFX4_248/Y OAI21X1_1/A BUFX2_958/A gnd OAI21X1_187/C vdd OAI21X1
XFILL_0_BUFX2_918 gnd vdd FILL
XFILL_0_DFFPOSX1_1031 gnd vdd FILL
XINVX1_206 OR2X2_19/Y gnd INVX1_206/Y vdd INVX1
XINVX1_217 INVX1_217/A gnd INVX1_217/Y vdd INVX1
XOAI21X1_197 BUFX4_134/Y INVX2_6/Y OAI21X1_197/C gnd OAI21X1_197/Y vdd OAI21X1
XOAI21X1_175 BUFX4_144/Y INVX2_197/Y OAI21X1_175/C gnd OAI21X1_175/Y vdd OAI21X1
XFILL_9_2_1 gnd vdd FILL
XNAND2X1_17 BUFX2_904/A BUFX4_224/Y gnd OAI21X1_17/C vdd NAND2X1
XNAND2X1_39 BUFX2_866/A BUFX4_230/Y gnd OAI21X1_39/C vdd NAND2X1
XNAND2X1_28 BUFX2_854/A BUFX4_233/Y gnd OAI21X1_28/C vdd NAND2X1
XNAND2X1_170 BUFX2_466/A BUFX4_236/Y gnd OAI21X1_425/C vdd NAND2X1
XNAND2X1_192 bundleStartMajId_i[38] bundleStartMajId_i[37] gnd OR2X2_4/A vdd NAND2X1
XFILL_0_XNOR2X1_35 gnd vdd FILL
XFILL_0_XNOR2X1_13 gnd vdd FILL
XFILL_0_XNOR2X1_24 gnd vdd FILL
XNAND2X1_181 AND2X2_2/Y AND2X2_1/Y gnd NOR2X1_23/A vdd NAND2X1
XFILL_0_XNOR2X1_57 gnd vdd FILL
XFILL_4_DFFPOSX1_791 gnd vdd FILL
XFILL_0_XNOR2X1_79 gnd vdd FILL
XFILL_0_XNOR2X1_46 gnd vdd FILL
XFILL_0_XNOR2X1_68 gnd vdd FILL
XFILL_4_DFFPOSX1_780 gnd vdd FILL
XFILL_1_OAI21X1_90 gnd vdd FILL
XFILL_17_1_1 gnd vdd FILL
XFILL_0_BUFX4_200 gnd vdd FILL
XFILL_1_BUFX2_681 gnd vdd FILL
XOAI21X1_1405 OAI21X1_1405/A BUFX4_290/Y OAI21X1_1405/C gnd OAI21X1_1405/Y vdd OAI21X1
XFILL_0_BUFX4_211 gnd vdd FILL
XFILL_0_BUFX4_222 gnd vdd FILL
XFILL_0_BUFX4_233 gnd vdd FILL
XFILL_1_OAI21X1_1614 gnd vdd FILL
XFILL_1_OAI21X1_1603 gnd vdd FILL
XOAI21X1_1427 OAI21X1_1427/A INVX1_221/A OAI21X1_1427/C gnd OAI21X1_1427/Y vdd OAI21X1
XOAI21X1_1416 BUFX4_171/Y BUFX4_64/Y BUFX2_196/A gnd OAI21X1_1417/C vdd OAI21X1
XOAI21X1_1438 NAND2X1_628/Y BUFX4_291/Y OAI21X1_1438/C gnd OAI21X1_1438/Y vdd OAI21X1
XFILL_0_BUFX4_255 gnd vdd FILL
XFILL_0_BUFX4_266 gnd vdd FILL
XFILL_0_BUFX4_244 gnd vdd FILL
XFILL_1_BUFX2_692 gnd vdd FILL
XFILL_1_OAI21X1_1647 gnd vdd FILL
XFILL_1_OAI21X1_1636 gnd vdd FILL
XFILL_1_OAI21X1_1625 gnd vdd FILL
XFILL_3_DFFPOSX1_381 gnd vdd FILL
XFILL_0_BUFX4_288 gnd vdd FILL
XFILL_0_BUFX4_299 gnd vdd FILL
XOAI21X1_1449 OR2X2_17/Y NOR2X1_222/B OAI21X1_1449/C gnd OAI21X1_1451/A vdd OAI21X1
XFILL_0_BUFX4_277 gnd vdd FILL
XNOR3X1_5 bundleStartMajId_i[24] NOR3X1_5/B NOR3X1_5/C gnd NOR3X1_5/Y vdd NOR3X1
XFILL_3_DFFPOSX1_370 gnd vdd FILL
XFILL_1_OAI21X1_1658 gnd vdd FILL
XFILL_1_OAI21X1_1669 gnd vdd FILL
XFILL_3_DFFPOSX1_392 gnd vdd FILL
XFILL_1_OAI21X1_609 gnd vdd FILL
XFILL_0_OAI21X1_438 gnd vdd FILL
XFILL_0_OAI21X1_427 gnd vdd FILL
XFILL_0_OAI21X1_416 gnd vdd FILL
XFILL_0_OAI21X1_405 gnd vdd FILL
XFILL_0_OAI21X1_449 gnd vdd FILL
XFILL_6_DFFPOSX1_830 gnd vdd FILL
XFILL_0_INVX4_30 gnd vdd FILL
XFILL_3_DFFPOSX1_1013 gnd vdd FILL
XFILL_6_DFFPOSX1_841 gnd vdd FILL
XFILL_3_DFFPOSX1_1024 gnd vdd FILL
XFILL_6_DFFPOSX1_852 gnd vdd FILL
XFILL_3_DFFPOSX1_1002 gnd vdd FILL
XFILL_0_INVX4_41 gnd vdd FILL
XFILL_6_DFFPOSX1_863 gnd vdd FILL
XFILL_6_DFFPOSX1_874 gnd vdd FILL
XXNOR2X1_92 INVX1_221/A bundleAddress_i[48] gnd XNOR2X1_92/Y vdd XNOR2X1
XXNOR2X1_81 OR2X2_20/A bundleAddress_i[32] gnd XNOR2X1_81/Y vdd XNOR2X1
XXNOR2X1_70 INVX1_193/A INVX8_3/Y gnd XNOR2X1_70/Y vdd XNOR2X1
XFILL_37_9_0 gnd vdd FILL
XFILL_0_NAND2X1_400 gnd vdd FILL
XFILL_1_XNOR2X1_4 gnd vdd FILL
XFILL_0_OAI21X1_1215 gnd vdd FILL
XFILL_0_NAND2X1_411 gnd vdd FILL
XFILL_0_NAND2X1_433 gnd vdd FILL
XFILL_0_OAI21X1_1204 gnd vdd FILL
XFILL_0_NAND2X1_444 gnd vdd FILL
XFILL_0_NAND2X1_422 gnd vdd FILL
XFILL_0_NAND2X1_466 gnd vdd FILL
XFILL_0_OAI21X1_1237 gnd vdd FILL
XFILL_0_OAI21X1_1226 gnd vdd FILL
XFILL_0_DFFPOSX1_816 gnd vdd FILL
XFILL_0_NAND2X1_477 gnd vdd FILL
XFILL_0_OAI21X1_1248 gnd vdd FILL
XFILL_1_NAND2X1_637 gnd vdd FILL
XFILL_0_NAND2X1_455 gnd vdd FILL
XFILL_0_DFFPOSX1_805 gnd vdd FILL
XBUFX2_80 BUFX2_80/A gnd addr2_o[41] vdd BUFX2
XBUFX2_91 BUFX2_91/A gnd addr2_o[31] vdd BUFX2
XFILL_0_OAI21X1_1259 gnd vdd FILL
XFILL_0_NAND2X1_488 gnd vdd FILL
XFILL_0_NAND2X1_499 gnd vdd FILL
XFILL_0_DFFPOSX1_838 gnd vdd FILL
XFILL_0_DFFPOSX1_849 gnd vdd FILL
XFILL_0_DFFPOSX1_827 gnd vdd FILL
XFILL_5_DFFPOSX1_420 gnd vdd FILL
XFILL_20_8_0 gnd vdd FILL
XFILL_5_DFFPOSX1_431 gnd vdd FILL
XFILL_5_DFFPOSX1_442 gnd vdd FILL
XFILL_5_DFFPOSX1_453 gnd vdd FILL
XFILL_24_15_1 gnd vdd FILL
XFILL_5_DFFPOSX1_486 gnd vdd FILL
XFILL_5_DFFPOSX1_497 gnd vdd FILL
XFILL_5_DFFPOSX1_464 gnd vdd FILL
XFILL_5_DFFPOSX1_475 gnd vdd FILL
XFILL_1_BUFX4_80 gnd vdd FILL
XFILL_1_BUFX4_91 gnd vdd FILL
XFILL_0_AOI21X1_13 gnd vdd FILL
XFILL_0_AOI21X1_24 gnd vdd FILL
XFILL_0_AOI21X1_46 gnd vdd FILL
XFILL_0_AOI21X1_35 gnd vdd FILL
XFILL_0_AOI21X1_57 gnd vdd FILL
XFILL_0_OAI21X1_950 gnd vdd FILL
XFILL_2_CLKBUF1_4 gnd vdd FILL
XFILL_0_OAI21X1_961 gnd vdd FILL
XFILL_0_OAI21X1_983 gnd vdd FILL
XFILL_0_OAI21X1_972 gnd vdd FILL
XFILL_0_OAI21X1_994 gnd vdd FILL
XFILL_28_9_0 gnd vdd FILL
XFILL_3_9_0 gnd vdd FILL
XFILL_2_BUFX4_131 gnd vdd FILL
XFILL_6_DFFPOSX1_1017 gnd vdd FILL
XFILL_6_DFFPOSX1_1006 gnd vdd FILL
XFILL_2_MUX2X1_2 gnd vdd FILL
XFILL_29_14_1 gnd vdd FILL
XFILL_0_OAI21X1_1760 gnd vdd FILL
XFILL_0_OAI21X1_1793 gnd vdd FILL
XFILL_0_OAI21X1_1782 gnd vdd FILL
XFILL_0_OAI21X1_1771 gnd vdd FILL
XFILL_11_8_0 gnd vdd FILL
XFILL_0_BUFX2_715 gnd vdd FILL
XFILL_23_10_0 gnd vdd FILL
XFILL_0_NOR2X1_33 gnd vdd FILL
XFILL_0_NOR2X1_22 gnd vdd FILL
XFILL_0_NOR2X1_11 gnd vdd FILL
XFILL_0_BUFX2_704 gnd vdd FILL
XFILL_0_BUFX2_726 gnd vdd FILL
XFILL_0_BUFX2_748 gnd vdd FILL
XFILL_0_NOR2X1_44 gnd vdd FILL
XFILL_0_NOR2X1_55 gnd vdd FILL
XFILL_0_BUFX2_737 gnd vdd FILL
XFILL_0_NOR2X1_66 gnd vdd FILL
XFILL_0_BUFX2_759 gnd vdd FILL
XFILL_0_NOR2X1_99 gnd vdd FILL
XFILL_0_NOR2X1_77 gnd vdd FILL
XFILL_0_NOR2X1_88 gnd vdd FILL
XFILL_6_DFFPOSX1_104 gnd vdd FILL
XFILL_6_DFFPOSX1_126 gnd vdd FILL
XFILL_6_DFFPOSX1_115 gnd vdd FILL
XFILL_6_DFFPOSX1_137 gnd vdd FILL
XFILL_6_DFFPOSX1_148 gnd vdd FILL
XFILL_6_DFFPOSX1_159 gnd vdd FILL
XBUFX4_312 BUFX4_386/A gnd BUFX4_312/Y vdd BUFX4
XBUFX4_301 BUFX4_303/A gnd BUFX4_301/Y vdd BUFX4
XFILL_0_INVX2_200 gnd vdd FILL
XFILL_2_OAI21X1_1810 gnd vdd FILL
XBUFX4_323 BUFX4_376/A gnd BUFX4_323/Y vdd BUFX4
XBUFX4_334 BUFX4_378/A gnd BUFX4_334/Y vdd BUFX4
XFILL_19_9_0 gnd vdd FILL
XBUFX4_345 BUFX4_388/A gnd BUFX4_345/Y vdd BUFX4
XFILL_4_15_1 gnd vdd FILL
XBUFX4_356 BUFX4_385/A gnd BUFX4_356/Y vdd BUFX4
XBUFX4_378 BUFX4_378/A gnd BUFX4_378/Y vdd BUFX4
XBUFX4_367 BUFX4_376/A gnd BUFX4_367/Y vdd BUFX4
XFILL_19_3 gnd vdd FILL
XOAI21X1_1213 BUFX4_132/Y INVX4_32/Y OAI21X1_1213/C gnd OAI21X1_1213/Y vdd OAI21X1
XOAI21X1_1202 NOR3X1_15/C INVX4_49/Y BUFX4_243/Y gnd OAI21X1_1203/B vdd OAI21X1
XDFFPOSX1_814 BUFX2_121/A CLKBUF1_12/Y OAI21X1_1111/Y gnd vdd DFFPOSX1
XOAI21X1_1224 OAI21X1_1224/A BUFX4_126/Y OAI21X1_1224/C gnd OAI21X1_1224/Y vdd OAI21X1
XFILL_1_OAI21X1_1433 gnd vdd FILL
XOAI21X1_1235 XNOR2X1_75/Y BUFX4_132/Y OAI21X1_1235/C gnd OAI21X1_1235/Y vdd OAI21X1
XOAI21X1_1246 INVX1_201/A NOR2X1_183/A INVX2_66/Y gnd OAI21X1_1247/C vdd OAI21X1
XFILL_1_OAI21X1_1422 gnd vdd FILL
XFILL_1_OAI21X1_1400 gnd vdd FILL
XFILL_1_OAI21X1_1411 gnd vdd FILL
XDFFPOSX1_803 BUFX2_56/A CLKBUF1_97/Y OAI21X1_1095/Y gnd vdd DFFPOSX1
XOAI21X1_1257 BUFX4_94/Y BUFX4_340/Y BUFX2_138/A gnd OAI21X1_1258/C vdd OAI21X1
XDFFPOSX1_825 BUFX2_74/A CLKBUF1_23/Y OAI21X1_1131/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1466 gnd vdd FILL
XFILL_1_CLKBUF1_91 gnd vdd FILL
XDFFPOSX1_836 BUFX2_86/A CLKBUF1_50/Y OAI21X1_1148/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1455 gnd vdd FILL
XFILL_1_CLKBUF1_80 gnd vdd FILL
XOAI21X1_1279 AND2X2_27/A INVX4_37/Y MUX2X1_2/S gnd OAI21X1_1280/B vdd OAI21X1
XOAI21X1_1268 NOR3X1_18/C OR2X2_18/A OR2X2_18/B gnd OAI21X1_1269/C vdd OAI21X1
XFILL_1_OAI21X1_1444 gnd vdd FILL
XDFFPOSX1_847 BUFX2_98/A CLKBUF1_53/Y OAI21X1_1164/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_202 gnd vdd FILL
XFILL_0_OAI21X1_224 gnd vdd FILL
XFILL_0_OAI21X1_235 gnd vdd FILL
XFILL_0_OAI21X1_246 gnd vdd FILL
XFILL_1_OAI21X1_1477 gnd vdd FILL
XDFFPOSX1_869 BUFX2_123/A CLKBUF1_97/Y OAI21X1_1203/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_213 gnd vdd FILL
XDFFPOSX1_858 BUFX2_111/A CLKBUF1_85/Y OAI21X1_1181/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_406 gnd vdd FILL
XFILL_1_OAI21X1_417 gnd vdd FILL
XFILL_1_OAI21X1_1488 gnd vdd FILL
XFILL_1_OAI21X1_1499 gnd vdd FILL
XFILL_0_OAI21X1_268 gnd vdd FILL
XFILL_0_OAI21X1_279 gnd vdd FILL
XFILL_1_OAI21X1_428 gnd vdd FILL
XINVX2_19 bundleStartMajId_i[44] gnd OR2X2_5/B vdd INVX2
XFILL_0_OAI21X1_257 gnd vdd FILL
XFILL_1_OAI21X1_439 gnd vdd FILL
XFILL_9_14_1 gnd vdd FILL
XFILL_3_10_0 gnd vdd FILL
XFILL_1_NAND2X1_412 gnd vdd FILL
XFILL_0_OAI21X1_1023 gnd vdd FILL
XFILL_0_NAND2X1_241 gnd vdd FILL
XFILL_0_NAND2X1_252 gnd vdd FILL
XFILL_0_NAND2X1_230 gnd vdd FILL
XFILL_0_OAI21X1_1001 gnd vdd FILL
XFILL_0_OAI21X1_1012 gnd vdd FILL
XFILL_0_OAI21X1_1045 gnd vdd FILL
XFILL_0_DFFPOSX1_624 gnd vdd FILL
XFILL_0_DFFPOSX1_613 gnd vdd FILL
XFILL_0_NAND2X1_263 gnd vdd FILL
XFILL_1_BUFX4_209 gnd vdd FILL
XFILL_0_NAND2X1_285 gnd vdd FILL
XFILL_0_DFFPOSX1_602 gnd vdd FILL
XFILL_0_NAND2X1_274 gnd vdd FILL
XFILL_0_OAI21X1_1034 gnd vdd FILL
XFILL_0_OAI21X1_1056 gnd vdd FILL
XFILL_1_NAND2X1_478 gnd vdd FILL
XFILL_1_NAND2X1_489 gnd vdd FILL
XFILL_0_OAI21X1_1067 gnd vdd FILL
XFILL_0_NAND2X1_296 gnd vdd FILL
XFILL_0_OAI21X1_1078 gnd vdd FILL
XFILL_0_OAI21X1_1089 gnd vdd FILL
XFILL_0_DFFPOSX1_635 gnd vdd FILL
XFILL_0_DFFPOSX1_657 gnd vdd FILL
XFILL_0_DFFPOSX1_646 gnd vdd FILL
XFILL_0_DFFPOSX1_679 gnd vdd FILL
XFILL_0_DFFPOSX1_668 gnd vdd FILL
XFILL_5_DFFPOSX1_261 gnd vdd FILL
XFILL_5_DFFPOSX1_272 gnd vdd FILL
XFILL_5_DFFPOSX1_250 gnd vdd FILL
XFILL_5_DFFPOSX1_283 gnd vdd FILL
XFILL_5_DFFPOSX1_294 gnd vdd FILL
XOAI21X1_1791 BUFX4_385/Y INVX2_163/Y NAND2X1_732/Y gnd OAI21X1_1791/Y vdd OAI21X1
XOAI21X1_1780 BUFX4_344/Y INVX2_152/Y NAND2X1_721/Y gnd OAI21X1_1780/Y vdd OAI21X1
XFILL_2_BUFX4_14 gnd vdd FILL
XFILL_1_OAI21X1_940 gnd vdd FILL
XFILL_1_OAI21X1_951 gnd vdd FILL
XFILL_0_OAI21X1_780 gnd vdd FILL
XFILL_0_OAI21X1_791 gnd vdd FILL
XFILL_1_OR2X2_3 gnd vdd FILL
XFILL_1_OAI21X1_962 gnd vdd FILL
XFILL_1_OAI21X1_973 gnd vdd FILL
XFILL_1_OAI21X1_984 gnd vdd FILL
XFILL_1_OAI21X1_995 gnd vdd FILL
XFILL_6_0_1 gnd vdd FILL
XBUFX2_805 BUFX2_805/A gnd tid1_o[29] vdd BUFX2
XFILL_2_DFFPOSX1_718 gnd vdd FILL
XBUFX2_816 BUFX2_816/A gnd tid1_o[19] vdd BUFX2
XBUFX2_827 BUFX2_827/A gnd tid1_o[9] vdd BUFX2
XFILL_2_DFFPOSX1_729 gnd vdd FILL
XFILL_2_DFFPOSX1_707 gnd vdd FILL
XBUFX2_849 BUFX2_849/A gnd tid2_o[47] vdd BUFX2
XBUFX2_838 BUFX2_838/A gnd tid1_o[56] vdd BUFX2
XFILL_2_BUFX4_1 gnd vdd FILL
XFILL_0_OAI21X1_1590 gnd vdd FILL
XFILL_0_BUFX2_512 gnd vdd FILL
XFILL_0_BUFX2_501 gnd vdd FILL
XFILL_0_BUFX2_523 gnd vdd FILL
XFILL_1_DFFPOSX1_319 gnd vdd FILL
XFILL_1_DFFPOSX1_308 gnd vdd FILL
XFILL_0_BUFX2_545 gnd vdd FILL
XCLKBUF1_4 BUFX4_83/Y gnd CLKBUF1_4/Y vdd CLKBUF1
XFILL_0_BUFX2_534 gnd vdd FILL
XFILL_0_BUFX2_556 gnd vdd FILL
XFILL_0_BUFX2_578 gnd vdd FILL
XFILL_0_BUFX2_567 gnd vdd FILL
XFILL_0_BUFX2_589 gnd vdd FILL
XFILL_14_15_0 gnd vdd FILL
XBUFX4_120 INVX8_4/Y gnd BUFX4_384/A vdd BUFX4
XBUFX4_164 BUFX4_19/Y gnd BUFX4_164/Y vdd BUFX4
XBUFX4_142 BUFX4_17/Y gnd BUFX4_142/Y vdd BUFX4
XFILL_0_INVX1_42 gnd vdd FILL
XFILL_0_INVX1_31 gnd vdd FILL
XFILL_4_CLKBUF1_24 gnd vdd FILL
XFILL_0_INVX1_20 gnd vdd FILL
XFILL_4_CLKBUF1_13 gnd vdd FILL
XBUFX4_153 BUFX4_13/Y gnd BUFX4_153/Y vdd BUFX4
XBUFX4_131 BUFX4_13/Y gnd BUFX4_131/Y vdd BUFX4
XFILL_1_AND2X2_1 gnd vdd FILL
XBUFX4_197 BUFX4_24/Y gnd BUFX4_197/Y vdd BUFX4
XFILL_0_INVX1_53 gnd vdd FILL
XFILL_4_CLKBUF1_57 gnd vdd FILL
XFILL_4_CLKBUF1_68 gnd vdd FILL
XNOR2X1_224 INVX1_189/A INVX4_51/Y gnd INVX2_109/A vdd NOR2X1
XFILL_4_CLKBUF1_35 gnd vdd FILL
XBUFX4_175 BUFX4_19/Y gnd BUFX4_175/Y vdd BUFX4
XNOR2X1_213 INVX2_91/Y INVX2_92/Y gnd INVX1_218/A vdd NOR2X1
XNOR2X1_202 BUFX4_160/Y NOR3X1_17/Y gnd NOR2X1_202/Y vdd NOR2X1
XFILL_2_OAI21X1_1673 gnd vdd FILL
XFILL_0_INVX1_75 gnd vdd FILL
XFILL_0_INVX1_64 gnd vdd FILL
XFILL_0_INVX1_86 gnd vdd FILL
XBUFX4_186 BUFX4_26/Y gnd BUFX4_186/Y vdd BUFX4
XFILL_4_CLKBUF1_46 gnd vdd FILL
XFILL_34_7_0 gnd vdd FILL
XFILL_0_INVX1_97 gnd vdd FILL
XFILL_31_2 gnd vdd FILL
XFILL_4_CLKBUF1_79 gnd vdd FILL
XFILL_0_BUFX2_17 gnd vdd FILL
XFILL_0_BUFX2_28 gnd vdd FILL
XFILL_0_BUFX2_39 gnd vdd FILL
XFILL_24_1 gnd vdd FILL
XOAI21X1_708 XNOR2X1_43/Y BUFX4_300/Y OAI21X1_708/C gnd OAI21X1_708/Y vdd OAI21X1
XOAI21X1_719 BUFX4_177/Y BUFX4_41/Y BUFX2_599/A gnd OAI21X1_720/C vdd OAI21X1
XOAI21X1_1021 BUFX4_296/Y INVX1_165/Y OAI21X1_1021/C gnd OAI21X1_1021/Y vdd OAI21X1
XOAI21X1_1010 BUFX4_158/Y BUFX4_39/Y BUFX2_368/A gnd OAI21X1_1011/C vdd OAI21X1
XOAI21X1_1032 BUFX4_172/Y BUFX4_55/Y BUFX2_381/A gnd OAI21X1_1033/C vdd OAI21X1
XOAI21X1_1043 BUFX4_353/Y INVX2_60/Y NAND2X1_409/Y gnd OAI21X1_1043/Y vdd OAI21X1
XFILL_1_OAI21X1_1230 gnd vdd FILL
XFILL_1_OAI21X1_1241 gnd vdd FILL
XDFFPOSX1_600 BUFX2_633/A CLKBUF1_72/Y OAI21X1_813/Y gnd vdd DFFPOSX1
XOAI21X1_1054 BUFX4_311/Y INVX2_69/Y NAND2X1_420/Y gnd OAI21X1_1054/Y vdd OAI21X1
XDFFPOSX1_611 BUFX2_645/A CLKBUF1_9/Y OAI21X1_843/Y gnd vdd DFFPOSX1
XDFFPOSX1_622 INVX1_51/A CLKBUF1_6/Y OAI21X1_850/Y gnd vdd DFFPOSX1
XDFFPOSX1_655 BUFX2_322/A CLKBUF1_96/Y OAI21X1_883/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_820 gnd vdd FILL
XFILL_1_OAI21X1_1252 gnd vdd FILL
XDFFPOSX1_633 INVX1_62/A CLKBUF1_61/Y OAI21X1_861/Y gnd vdd DFFPOSX1
XOAI21X1_1065 BUFX4_377/Y INVX4_38/Y NAND2X1_431/Y gnd OAI21X1_1065/Y vdd OAI21X1
XOAI21X1_1098 BUFX4_360/Y INVX2_92/Y NAND2X1_464/Y gnd OAI21X1_1098/Y vdd OAI21X1
XFILL_1_OAI21X1_1263 gnd vdd FILL
XFILL_1_OAI21X1_1274 gnd vdd FILL
XFILL_1_DFFPOSX1_842 gnd vdd FILL
XDFFPOSX1_644 INVX1_73/A CLKBUF1_10/Y OAI21X1_872/Y gnd vdd DFFPOSX1
XDFFPOSX1_666 BUFX2_303/A CLKBUF1_58/Y OAI21X1_894/Y gnd vdd DFFPOSX1
XOAI21X1_1076 BUFX4_350/Y INVX2_79/Y NAND2X1_442/Y gnd OAI21X1_1076/Y vdd OAI21X1
XFILL_1_DFFPOSX1_831 gnd vdd FILL
XOAI21X1_1087 BUFX4_364/Y INVX2_84/Y NAND2X1_453/Y gnd OAI21X1_1087/Y vdd OAI21X1
XFILL_1_OAI21X1_225 gnd vdd FILL
XFILL_1_DFFPOSX1_875 gnd vdd FILL
XDFFPOSX1_688 BUFX2_355/A CLKBUF1_61/Y OAI21X1_925/Y gnd vdd DFFPOSX1
XNAND2X1_703 BUFX2_695/A BUFX4_211/Y gnd NAND2X1_703/Y vdd NAND2X1
XFILL_1_OAI21X1_1285 gnd vdd FILL
XFILL_1_DFFPOSX1_853 gnd vdd FILL
XFILL_1_OAI21X1_1296 gnd vdd FILL
XFILL_1_OAI21X1_214 gnd vdd FILL
XFILL_1_DFFPOSX1_864 gnd vdd FILL
XDFFPOSX1_677 BUFX2_315/A CLKBUF1_81/Y OAI21X1_905/Y gnd vdd DFFPOSX1
XDFFPOSX1_699 BUFX2_336/A CLKBUF1_37/Y OAI21X1_947/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_203 gnd vdd FILL
XFILL_1_OAI21X1_269 gnd vdd FILL
XNAND2X1_736 BUFX2_791/A BUFX4_329/Y gnd NAND2X1_736/Y vdd NAND2X1
XFILL_1_OAI21X1_247 gnd vdd FILL
XNAND2X1_714 bundleLen_i[1] BUFX4_305/Y gnd BUFX4_303/A vdd NAND2X1
XFILL_1_DFFPOSX1_886 gnd vdd FILL
XFILL_1_OAI21X1_258 gnd vdd FILL
XFILL_19_14_0 gnd vdd FILL
XFILL_1_OAI21X1_236 gnd vdd FILL
XFILL_1_DFFPOSX1_897 gnd vdd FILL
XFILL_0_NOR2X1_8 gnd vdd FILL
XNAND2X1_725 BUFX2_779/A BUFX4_326/Y gnd NAND2X1_725/Y vdd NAND2X1
XNAND2X1_769 BUFX2_827/A BUFX4_352/Y gnd NAND2X1_769/Y vdd NAND2X1
XNAND2X1_758 BUFX2_815/A BUFX4_313/Y gnd NAND2X1_758/Y vdd NAND2X1
XNAND2X1_747 BUFX2_803/A BUFX4_320/Y gnd NAND2X1_747/Y vdd NAND2X1
XFILL_6_DFFPOSX1_490 gnd vdd FILL
XFILL_32_16_0 gnd vdd FILL
XFILL_25_7_0 gnd vdd FILL
XFILL_0_7_0 gnd vdd FILL
XFILL_1_NAND2X1_264 gnd vdd FILL
XFILL_0_DFFPOSX1_421 gnd vdd FILL
XFILL_0_DFFPOSX1_410 gnd vdd FILL
XFILL_1_NAND2X1_275 gnd vdd FILL
XFILL_0_DFFPOSX1_432 gnd vdd FILL
XFILL_1_NAND2X1_297 gnd vdd FILL
XFILL_0_DFFPOSX1_443 gnd vdd FILL
XFILL_0_DFFPOSX1_465 gnd vdd FILL
XFILL_2_DFFPOSX1_7 gnd vdd FILL
XFILL_0_DFFPOSX1_454 gnd vdd FILL
XFILL_0_DFFPOSX1_476 gnd vdd FILL
XINVX8_6 INVX8_6/A gnd INVX8_6/Y vdd INVX8
XFILL_0_DFFPOSX1_498 gnd vdd FILL
XFILL_0_DFFPOSX1_487 gnd vdd FILL
XFILL_3_DFFPOSX1_903 gnd vdd FILL
XFILL_3_DFFPOSX1_914 gnd vdd FILL
XFILL_3_DFFPOSX1_936 gnd vdd FILL
XFILL_3_DFFPOSX1_947 gnd vdd FILL
XFILL_3_DFFPOSX1_925 gnd vdd FILL
XFILL_3_DFFPOSX1_969 gnd vdd FILL
XFILL_3_DFFPOSX1_958 gnd vdd FILL
XDFFPOSX1_70 BUFX2_757/A CLKBUF1_8/Y DFFPOSX1_70/D gnd vdd DFFPOSX1
XDFFPOSX1_81 BUFX2_750/A CLKBUF1_55/Y DFFPOSX1_81/D gnd vdd DFFPOSX1
XDFFPOSX1_92 BUFX2_762/A CLKBUF1_3/Y DFFPOSX1_92/D gnd vdd DFFPOSX1
XFILL_37_15_0 gnd vdd FILL
XFILL_8_8_0 gnd vdd FILL
XFILL_1_OAI21X1_781 gnd vdd FILL
XBUFX4_26 BUFX4_26/A gnd BUFX4_26/Y vdd BUFX4
XBUFX4_15 INVX8_6/Y gnd BUFX4_15/Y vdd BUFX4
XFILL_1_OAI21X1_770 gnd vdd FILL
XFILL_2_OAI21X1_985 gnd vdd FILL
XBUFX4_48 BUFX4_64/A gnd BUFX4_48/Y vdd BUFX4
XBUFX4_59 BUFX4_59/A gnd BUFX4_59/Y vdd BUFX4
XBUFX4_37 BUFX4_82/A gnd BUFX4_37/Y vdd BUFX4
XFILL_1_OAI21X1_792 gnd vdd FILL
XFILL_2_DFFPOSX1_504 gnd vdd FILL
XBUFX2_602 BUFX2_602/A gnd majID4_o[39] vdd BUFX2
XFILL_2_DFFPOSX1_515 gnd vdd FILL
XBUFX2_613 BUFX2_613/A gnd majID4_o[29] vdd BUFX2
XFILL_2_DFFPOSX1_537 gnd vdd FILL
XFILL_2_DFFPOSX1_526 gnd vdd FILL
XBUFX2_646 BUFX2_646/A gnd majID4_o[56] vdd BUFX2
XBUFX2_624 BUFX2_624/A gnd majID4_o[19] vdd BUFX2
XBUFX2_635 BUFX2_635/A gnd majID4_o[9] vdd BUFX2
XBUFX2_657 BUFX2_657/A gnd pid1_o[15] vdd BUFX2
XBUFX2_679 BUFX2_679/A gnd pid1_o[23] vdd BUFX2
XFILL_2_DFFPOSX1_548 gnd vdd FILL
XBUFX2_668 BUFX2_668/A gnd pid1_o[5] vdd BUFX2
XFILL_16_7_0 gnd vdd FILL
XFILL_2_DFFPOSX1_559 gnd vdd FILL
XFILL_0_BUFX2_331 gnd vdd FILL
XINVX2_131 bundlePid_i[17] gnd INVX2_131/Y vdd INVX2
XFILL_0_BUFX2_320 gnd vdd FILL
XOR2X2_18 OR2X2_18/A OR2X2_18/B gnd OR2X2_18/Y vdd OR2X2
XINVX2_120 bundlePid_i[28] gnd INVX2_120/Y vdd INVX2
XFILL_1_DFFPOSX1_127 gnd vdd FILL
XFILL_0_BUFX2_342 gnd vdd FILL
XFILL_1_DFFPOSX1_138 gnd vdd FILL
XINVX2_164 bundleTid_i[45] gnd INVX2_164/Y vdd INVX2
XFILL_0_BUFX2_375 gnd vdd FILL
XFILL_1_DFFPOSX1_116 gnd vdd FILL
XINVX2_153 bundleTid_i[56] gnd INVX2_153/Y vdd INVX2
XFILL_0_BUFX2_364 gnd vdd FILL
XINVX2_175 bundleTid_i[34] gnd INVX2_175/Y vdd INVX2
XINVX2_142 bundlePid_i[6] gnd INVX2_142/Y vdd INVX2
XFILL_1_DFFPOSX1_105 gnd vdd FILL
XFILL_0_BUFX2_353 gnd vdd FILL
XFILL_1_DFFPOSX1_149 gnd vdd FILL
XINVX2_197 bundleTid_i[12] gnd INVX2_197/Y vdd INVX2
XFILL_0_BUFX2_386 gnd vdd FILL
XINVX2_186 bundleTid_i[23] gnd INVX2_186/Y vdd INVX2
XFILL_0_BUFX2_397 gnd vdd FILL
XFILL_4_DFFPOSX1_609 gnd vdd FILL
XFILL_2_OAI21X1_1481 gnd vdd FILL
XOAI21X1_505 OAI21X1_505/A BUFX4_135/Y OAI21X1_505/C gnd OAI21X1_505/Y vdd OAI21X1
XOAI21X1_538 OAI22X1_1/Y BUFX4_167/Y OAI21X1_538/C gnd OAI21X1_538/Y vdd OAI21X1
XOAI21X1_527 INVX4_30/Y INVX4_3/Y INVX2_15/Y gnd OAI21X1_528/C vdd OAI21X1
XOAI21X1_516 BUFX4_7/A BUFX4_388/Y BUFX2_577/A gnd OAI21X1_517/C vdd OAI21X1
XOAI21X1_549 OR2X2_10/B INVX4_7/Y INVX2_18/Y gnd OAI21X1_550/C vdd OAI21X1
XFILL_21_13_1 gnd vdd FILL
XFILL_1_NAND3X1_60 gnd vdd FILL
XDFFPOSX1_430 BUFX2_459/A CLKBUF1_13/Y OAI21X1_415/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_650 gnd vdd FILL
XFILL_1_OAI21X1_1082 gnd vdd FILL
XDFFPOSX1_463 BUFX2_495/A CLKBUF1_22/Y OAI21X1_464/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1071 gnd vdd FILL
XDFFPOSX1_452 BUFX2_483/A CLKBUF1_92/Y OAI21X1_449/Y gnd vdd DFFPOSX1
XDFFPOSX1_441 BUFX2_471/A CLKBUF1_18/Y OAI21X1_432/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1060 gnd vdd FILL
XDFFPOSX1_474 BUFX2_507/A CLKBUF1_48/Y OAI21X1_483/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_672 gnd vdd FILL
XFILL_1_DFFPOSX1_683 gnd vdd FILL
XNAND2X1_500 bundleAddress_i[47] bundleAddress_i[46] gnd NOR2X1_133/B vdd NAND2X1
XFILL_1_DFFPOSX1_661 gnd vdd FILL
XDFFPOSX1_485 BUFX2_522/A CLKBUF1_94/Y OAI21X1_503/Y gnd vdd DFFPOSX1
XNAND2X1_511 BUFX2_81/A BUFX4_192/Y gnd NAND2X1_511/Y vdd NAND2X1
XFILL_1_OAI21X1_1093 gnd vdd FILL
XDFFPOSX1_496 BUFX2_525/A CLKBUF1_46/Y OAI21X1_536/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_694 gnd vdd FILL
XNAND2X1_522 BUFX2_85/A BUFX4_229/Y gnd NAND2X1_522/Y vdd NAND2X1
XNAND2X1_533 AND2X2_23/B INVX1_188/A gnd NOR2X1_160/B vdd NAND2X1
XNAND2X1_544 BUFX2_98/A BUFX4_189/Y gnd NAND2X1_544/Y vdd NAND2X1
XNAND2X1_555 BUFX2_105/A BUFX4_203/Y gnd NAND2X1_555/Y vdd NAND2X1
XNAND2X1_588 BUFX4_243/Y NAND2X1_588/B gnd NAND2X1_588/Y vdd NAND2X1
XFILL_2_OAI21X1_259 gnd vdd FILL
XFILL_1_OAI22X1_2 gnd vdd FILL
XNAND2X1_566 BUFX4_242/Y NOR3X1_14/C gnd NAND2X1_566/Y vdd NAND2X1
XNAND2X1_577 BUFX2_116/A BUFX4_201/Y gnd NAND2X1_577/Y vdd NAND2X1
XNAND2X1_599 INVX1_202/Y NOR2X1_187/B gnd MUX2X1_2/A vdd NAND2X1
XFILL_0_AND2X2_23 gnd vdd FILL
XFILL_0_AND2X2_12 gnd vdd FILL
XFILL_0_DFFPOSX1_240 gnd vdd FILL
XFILL_0_DFFPOSX1_273 gnd vdd FILL
XFILL_0_DFFPOSX1_262 gnd vdd FILL
XFILL_0_DFFPOSX1_284 gnd vdd FILL
XFILL_0_DFFPOSX1_251 gnd vdd FILL
XFILL_26_12_1 gnd vdd FILL
XFILL_0_DFFPOSX1_295 gnd vdd FILL
XFILL_3_DFFPOSX1_700 gnd vdd FILL
XFILL_3_DFFPOSX1_711 gnd vdd FILL
XFILL_3_DFFPOSX1_722 gnd vdd FILL
XFILL_3_DFFPOSX1_755 gnd vdd FILL
XFILL_3_DFFPOSX1_744 gnd vdd FILL
XFILL_3_CLKBUF1_32 gnd vdd FILL
XFILL_3_CLKBUF1_21 gnd vdd FILL
XFILL_3_DFFPOSX1_733 gnd vdd FILL
XFILL_3_CLKBUF1_10 gnd vdd FILL
XFILL_3_CLKBUF1_65 gnd vdd FILL
XFILL_3_CLKBUF1_43 gnd vdd FILL
XFILL_3_DFFPOSX1_788 gnd vdd FILL
XFILL_3_DFFPOSX1_777 gnd vdd FILL
XFILL_3_DFFPOSX1_799 gnd vdd FILL
XFILL_3_CLKBUF1_54 gnd vdd FILL
XFILL_3_DFFPOSX1_766 gnd vdd FILL
XFILL_3_CLKBUF1_76 gnd vdd FILL
XFILL_3_CLKBUF1_98 gnd vdd FILL
XFILL_3_CLKBUF1_87 gnd vdd FILL
XFILL_1_NOR2X1_150 gnd vdd FILL
XFILL_1_NOR2X1_161 gnd vdd FILL
XFILL_1_NOR2X1_172 gnd vdd FILL
XFILL_1_NOR2X1_194 gnd vdd FILL
XFILL_2_DFFPOSX1_301 gnd vdd FILL
XFILL_2_DFFPOSX1_312 gnd vdd FILL
XBUFX2_410 BUFX2_410/A gnd majID1_o[39] vdd BUFX2
XFILL_2_DFFPOSX1_345 gnd vdd FILL
XFILL_2_DFFPOSX1_323 gnd vdd FILL
XFILL_2_DFFPOSX1_356 gnd vdd FILL
XBUFX2_432 BUFX2_432/A gnd majID1_o[19] vdd BUFX2
XBUFX2_443 BUFX2_443/A gnd majID1_o[9] vdd BUFX2
XFILL_1_13_1 gnd vdd FILL
XBUFX2_421 BUFX2_421/A gnd majID1_o[29] vdd BUFX2
XBUFX2_454 BUFX2_454/A gnd majID1_o[56] vdd BUFX2
XFILL_2_DFFPOSX1_334 gnd vdd FILL
XBUFX2_487 BUFX2_487/A gnd majID2_o[27] vdd BUFX2
XBUFX2_476 BUFX2_476/A gnd majID2_o[37] vdd BUFX2
XFILL_2_DFFPOSX1_378 gnd vdd FILL
XFILL_2_DFFPOSX1_367 gnd vdd FILL
XBUFX2_465 BUFX2_465/A gnd majID2_o[47] vdd BUFX2
XFILL_2_DFFPOSX1_389 gnd vdd FILL
XBUFX2_498 BUFX2_498/A gnd majID2_o[17] vdd BUFX2
XFILL_5_DFFPOSX1_816 gnd vdd FILL
XFILL_31_5_0 gnd vdd FILL
XFILL_5_DFFPOSX1_805 gnd vdd FILL
XFILL_5_DFFPOSX1_827 gnd vdd FILL
XFILL_5_DFFPOSX1_838 gnd vdd FILL
XFILL_1_BUFX4_381 gnd vdd FILL
XFILL_1_BUFX4_370 gnd vdd FILL
XFILL_5_DFFPOSX1_849 gnd vdd FILL
XFILL_1_XNOR2X1_17 gnd vdd FILL
XFILL_1_XNOR2X1_28 gnd vdd FILL
XFILL_1_XNOR2X1_39 gnd vdd FILL
XFILL_0_BUFX2_150 gnd vdd FILL
XFILL_0_BUFX2_172 gnd vdd FILL
XFILL_0_BUFX2_183 gnd vdd FILL
XFILL_0_BUFX2_161 gnd vdd FILL
XFILL_0_BUFX2_194 gnd vdd FILL
XFILL_1_DFFPOSX1_4 gnd vdd FILL
XFILL_4_DFFPOSX1_406 gnd vdd FILL
XFILL_4_DFFPOSX1_428 gnd vdd FILL
XFILL_4_DFFPOSX1_417 gnd vdd FILL
XFILL_4_DFFPOSX1_439 gnd vdd FILL
XFILL_6_12_1 gnd vdd FILL
XFILL_2_DFFPOSX1_890 gnd vdd FILL
XFILL_1_BUFX2_318 gnd vdd FILL
XFILL_22_5_0 gnd vdd FILL
XFILL_1_BUFX2_307 gnd vdd FILL
XOAI21X1_313 INVX2_202/Y BUFX4_291/Y OAI21X1_313/C gnd OAI21X1_313/Y vdd OAI21X1
XOAI21X1_302 BUFX4_144/Y BUFX4_58/Y BUFX2_1016/A gnd OAI21X1_303/C vdd OAI21X1
XOAI21X1_346 BUFX4_351/Y INVX2_18/Y NAND2X1_90/Y gnd OAI21X1_346/Y vdd OAI21X1
XOAI21X1_324 BUFX4_134/Y BUFX4_72/Y BUFX2_1028/A gnd OAI21X1_325/C vdd OAI21X1
XOAI21X1_335 BUFX4_355/Y INVX2_13/Y NAND2X1_79/Y gnd OAI21X1_335/Y vdd OAI21X1
XOAI21X1_379 BUFX4_323/Y INVX2_34/Y OAI21X1_379/C gnd OAI21X1_379/Y vdd OAI21X1
XOAI21X1_368 BUFX4_358/Y INVX4_19/Y OAI21X1_368/C gnd OAI21X1_368/Y vdd OAI21X1
XOAI21X1_357 BUFX4_314/Y INVX4_14/Y OAI21X1_357/C gnd OAI21X1_357/Y vdd OAI21X1
XDFFPOSX1_282 BUFX2_955/A CLKBUF1_39/Y OAI21X1_181/Y gnd vdd DFFPOSX1
XDFFPOSX1_271 BUFX2_943/A CLKBUF1_57/Y OAI21X1_159/Y gnd vdd DFFPOSX1
XDFFPOSX1_260 BUFX2_931/A CLKBUF1_56/Y OAI21X1_137/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_480 gnd vdd FILL
XFILL_1_DFFPOSX1_491 gnd vdd FILL
XDFFPOSX1_293 BUFX2_970/A CLKBUF1_77/Y OAI21X1_203/Y gnd vdd DFFPOSX1
XNAND2X1_352 BUFX4_263/Y bundle_i[17] gnd OAI21X1_858/C vdd NAND2X1
XNAND2X1_330 INVX1_33/A INVX2_49/A gnd OAI21X1_793/B vdd NAND2X1
XFILL_3_NOR3X1_13 gnd vdd FILL
XNAND2X1_363 BUFX4_264/Y bundle_i[6] gnd OAI21X1_869/C vdd NAND2X1
XNAND2X1_341 INVX8_4/A bundle_i[28] gnd OAI21X1_847/C vdd NAND2X1
XFILL_4_DFFPOSX1_940 gnd vdd FILL
XNAND2X1_374 BUFX2_319/A BUFX4_217/Y gnd OAI21X1_880/C vdd NAND2X1
XNAND2X1_385 BUFX2_300/A BUFX4_206/Y gnd OAI21X1_891/C vdd NAND2X1
XNAND2X1_396 BUFX2_312/A BUFX4_232/Y gnd OAI21X1_902/C vdd NAND2X1
XFILL_5_6_0 gnd vdd FILL
XFILL_4_DFFPOSX1_962 gnd vdd FILL
XFILL_4_DFFPOSX1_951 gnd vdd FILL
XFILL_4_DFFPOSX1_973 gnd vdd FILL
XFILL_0_INVX1_117 gnd vdd FILL
XFILL_4_DFFPOSX1_984 gnd vdd FILL
XFILL_4_DFFPOSX1_995 gnd vdd FILL
XFILL_12_18_1 gnd vdd FILL
XFILL_0_INVX1_128 gnd vdd FILL
XFILL_0_INVX1_106 gnd vdd FILL
XFILL_0_INVX1_139 gnd vdd FILL
XFILL_1_AOI21X1_28 gnd vdd FILL
XFILL_1_AOI21X1_39 gnd vdd FILL
XFILL_1_AOI21X1_17 gnd vdd FILL
XFILL_13_5_0 gnd vdd FILL
XFILL_1_BUFX2_830 gnd vdd FILL
XFILL_1_BUFX2_874 gnd vdd FILL
XFILL_1_BUFX2_863 gnd vdd FILL
XFILL_1_OAI21X1_1807 gnd vdd FILL
XOAI21X1_1609 BUFX4_368/Y INVX2_145/Y NAND2X1_678/Y gnd OAI21X1_1609/Y vdd OAI21X1
XFILL_3_DFFPOSX1_530 gnd vdd FILL
XFILL_2_NOR3X1_5 gnd vdd FILL
XFILL_1_OAI21X1_1818 gnd vdd FILL
XFILL_3_DFFPOSX1_541 gnd vdd FILL
XFILL_3_DFFPOSX1_563 gnd vdd FILL
XFILL_1_OAI21X1_1829 gnd vdd FILL
XFILL_3_DFFPOSX1_574 gnd vdd FILL
XFILL_3_DFFPOSX1_552 gnd vdd FILL
XOAI21X1_880 INVX1_81/Y BUFX4_217/Y OAI21X1_880/C gnd OAI21X1_880/Y vdd OAI21X1
XOAI21X1_891 INVX1_92/Y BUFX4_206/Y OAI21X1_891/C gnd OAI21X1_891/Y vdd OAI21X1
XFILL_3_DFFPOSX1_585 gnd vdd FILL
XFILL_3_DFFPOSX1_596 gnd vdd FILL
XFILL_0_OAI21X1_609 gnd vdd FILL
XFILL_17_17_1 gnd vdd FILL
XFILL_7_3 gnd vdd FILL
XFILL_0_NAND2X1_626 gnd vdd FILL
XFILL_2_DFFPOSX1_131 gnd vdd FILL
XFILL_0_NAND2X1_604 gnd vdd FILL
XFILL_0_NAND2X1_615 gnd vdd FILL
XFILL_11_13_0 gnd vdd FILL
XFILL_2_DFFPOSX1_120 gnd vdd FILL
XFILL_2_DFFPOSX1_153 gnd vdd FILL
XFILL_0_NAND2X1_659 gnd vdd FILL
XFILL_2_DFFPOSX1_164 gnd vdd FILL
XFILL_0_NAND2X1_648 gnd vdd FILL
XFILL_0_OAI21X1_1408 gnd vdd FILL
XFILL_0_OAI21X1_1419 gnd vdd FILL
XBUFX2_251 BUFX2_251/A gnd addr4_o[2] vdd BUFX2
XBUFX2_262 INVX1_46/A gnd instr1_o[30] vdd BUFX2
XFILL_0_NAND2X1_637 gnd vdd FILL
XFILL_2_DFFPOSX1_142 gnd vdd FILL
XBUFX2_240 BUFX2_240/A gnd addr4_o[12] vdd BUFX2
XFILL_2_DFFPOSX1_175 gnd vdd FILL
XFILL_2_DFFPOSX1_197 gnd vdd FILL
XFILL_2_DFFPOSX1_186 gnd vdd FILL
XBUFX2_273 INVX1_47/A gnd instr1_o[29] vdd BUFX2
XBUFX2_295 BUFX2_295/A gnd instr2_o[21] vdd BUFX2
XBUFX2_284 INVX1_48/A gnd instr1_o[28] vdd BUFX2
XFILL_5_DFFPOSX1_602 gnd vdd FILL
XFILL_5_DFFPOSX1_624 gnd vdd FILL
XFILL_5_DFFPOSX1_613 gnd vdd FILL
XFILL_5_DFFPOSX1_635 gnd vdd FILL
XFILL_5_DFFPOSX1_646 gnd vdd FILL
XFILL_5_DFFPOSX1_679 gnd vdd FILL
XFILL_5_DFFPOSX1_668 gnd vdd FILL
XFILL_5_DFFPOSX1_657 gnd vdd FILL
XFILL_35_18_1 gnd vdd FILL
XFILL_4_DFFPOSX1_203 gnd vdd FILL
XNAND3X1_3 bundleStartMajId_i[35] bundleStartMajId_i[32] AND2X2_6/Y gnd NOR2X1_22/B
+ vdd NAND3X1
XFILL_4_DFFPOSX1_214 gnd vdd FILL
XFILL_4_DFFPOSX1_225 gnd vdd FILL
XFILL_16_12_0 gnd vdd FILL
XFILL_4_DFFPOSX1_236 gnd vdd FILL
XFILL_4_DFFPOSX1_258 gnd vdd FILL
XFILL_4_DFFPOSX1_247 gnd vdd FILL
XFILL_4_DFFPOSX1_269 gnd vdd FILL
XFILL_2_BUFX4_324 gnd vdd FILL
XFILL_2_CLKBUF1_40 gnd vdd FILL
XFILL_2_CLKBUF1_73 gnd vdd FILL
XFILL_2_CLKBUF1_84 gnd vdd FILL
XFILL_2_CLKBUF1_51 gnd vdd FILL
XFILL_2_CLKBUF1_62 gnd vdd FILL
XFILL_2_CLKBUF1_95 gnd vdd FILL
XFILL_1_BUFX2_104 gnd vdd FILL
XFILL_1_BUFX2_115 gnd vdd FILL
XOAI21X1_121 BUFX4_168/Y INVX2_170/Y OAI21X1_121/C gnd OAI21X1_121/Y vdd OAI21X1
XFILL_0_NOR2X1_180 gnd vdd FILL
XFILL_1_BUFX2_148 gnd vdd FILL
XOAI21X1_110 BUFX4_95/Y BUFX4_334/Y BUFX2_916/A gnd OAI21X1_111/C vdd OAI21X1
XFILL_0_NOR2X1_191 gnd vdd FILL
XFILL_1_BUFX2_159 gnd vdd FILL
XFILL_0_DFFPOSX1_1021 gnd vdd FILL
XOAI21X1_132 BUFX4_110/Y BUFX4_359/Y BUFX2_929/A gnd OAI21X1_133/C vdd OAI21X1
XOAI21X1_143 BUFX4_125/Y INVX2_181/Y OAI21X1_143/C gnd OAI21X1_143/Y vdd OAI21X1
XOAI21X1_165 BUFX4_134/Y INVX2_192/Y OAI21X1_165/C gnd OAI21X1_165/Y vdd OAI21X1
XOAI21X1_154 BUFX4_1/A BUFX4_374/Y BUFX2_941/A gnd OAI21X1_155/C vdd OAI21X1
XFILL_0_DFFPOSX1_1010 gnd vdd FILL
XFILL_0_BUFX2_908 gnd vdd FILL
XOAI21X1_187 BUFX4_168/Y INVX2_1/Y OAI21X1_187/C gnd OAI21X1_187/Y vdd OAI21X1
XFILL_0_DFFPOSX1_1032 gnd vdd FILL
XFILL_0_BUFX2_919 gnd vdd FILL
XINVX1_207 INVX1_207/A gnd INVX1_207/Y vdd INVX1
XOAI21X1_198 BUFX4_99/Y NAND2X1_7/B BUFX2_965/A gnd OAI21X1_199/C vdd OAI21X1
XOAI21X1_176 BUFX4_4/Y BUFX4_314/Y BUFX2_953/A gnd OAI21X1_177/C vdd OAI21X1
XINVX1_218 INVX1_218/A gnd INVX1_218/Y vdd INVX1
XFILL_6_DFFPOSX1_308 gnd vdd FILL
XFILL_6_DFFPOSX1_319 gnd vdd FILL
XFILL_34_13_0 gnd vdd FILL
XNAND2X1_29 BUFX2_855/A BUFX4_200/Y gnd OAI21X1_29/C vdd NAND2X1
XNAND2X1_171 bundleStartMajId_i[46] bundleStartMajId_i[45] gnd OR2X2_5/A vdd NAND2X1
XNAND2X1_160 BUFX2_461/A BUFX4_181/Y gnd OAI21X1_419/C vdd NAND2X1
XNAND2X1_18 BUFX2_843/A OAI21X1_9/B gnd OAI21X1_18/C vdd NAND2X1
XFILL_0_XNOR2X1_36 gnd vdd FILL
XFILL_0_XNOR2X1_25 gnd vdd FILL
XNAND2X1_182 bundleStartMajId_i[47] bundleStartMajId_i[44] gnd OR2X2_3/B vdd NAND2X1
XNAND2X1_193 BUFX2_477/A BUFX4_214/Y gnd OAI21X1_441/C vdd NAND2X1
XFILL_0_XNOR2X1_14 gnd vdd FILL
XFILL_0_XNOR2X1_58 gnd vdd FILL
XFILL_4_DFFPOSX1_792 gnd vdd FILL
XFILL_4_DFFPOSX1_770 gnd vdd FILL
XFILL_0_XNOR2X1_47 gnd vdd FILL
XFILL_0_XNOR2X1_69 gnd vdd FILL
XFILL_4_DFFPOSX1_781 gnd vdd FILL
XFILL_1_OAI21X1_80 gnd vdd FILL
XFILL_1_OAI21X1_91 gnd vdd FILL
XFILL_0_DFFPOSX1_1 gnd vdd FILL
XFILL_1_BUFX2_682 gnd vdd FILL
XFILL_0_BUFX4_223 gnd vdd FILL
XFILL_1_BUFX2_671 gnd vdd FILL
XFILL_1_BUFX2_660 gnd vdd FILL
XFILL_0_BUFX4_212 gnd vdd FILL
XFILL_0_BUFX4_201 gnd vdd FILL
XFILL_1_OAI21X1_1604 gnd vdd FILL
XFILL_1_OAI21X1_1615 gnd vdd FILL
XFILL_0_BUFX4_234 gnd vdd FILL
XOAI21X1_1406 INVX1_219/A bundleAddress_i[55] BUFX4_285/Y gnd OAI21X1_1408/B vdd OAI21X1
XOAI21X1_1417 XNOR2X1_91/Y BUFX4_289/Y OAI21X1_1417/C gnd OAI21X1_1417/Y vdd OAI21X1
XOAI21X1_1428 BUFX4_171/Y BUFX4_48/Y BUFX2_200/A gnd OAI21X1_1429/C vdd OAI21X1
XFILL_0_BUFX4_256 gnd vdd FILL
XFILL_0_BUFX4_267 gnd vdd FILL
XFILL_0_BUFX4_245 gnd vdd FILL
XFILL_1_OAI21X1_1637 gnd vdd FILL
XFILL_1_OAI21X1_1648 gnd vdd FILL
XFILL_0_BUFX4_289 gnd vdd FILL
XFILL_0_BUFX4_278 gnd vdd FILL
XFILL_3_DFFPOSX1_382 gnd vdd FILL
XFILL_1_OAI21X1_1626 gnd vdd FILL
XOAI21X1_1439 INVX4_51/Y INVX2_69/Y INVX4_35/Y gnd OAI21X1_1440/C vdd OAI21X1
XNOR3X1_6 NOR3X1_6/A NOR3X1_6/B OR2X2_9/Y gnd NOR3X1_6/Y vdd NOR3X1
XFILL_3_DFFPOSX1_360 gnd vdd FILL
XFILL_3_DFFPOSX1_371 gnd vdd FILL
XFILL_0_OAI21X1_428 gnd vdd FILL
XFILL_3_DFFPOSX1_393 gnd vdd FILL
XFILL_0_OAI21X1_406 gnd vdd FILL
XFILL_0_OAI21X1_417 gnd vdd FILL
XFILL_1_OAI21X1_1659 gnd vdd FILL
XFILL_0_INVX4_20 gnd vdd FILL
XFILL_0_OAI21X1_439 gnd vdd FILL
XFILL_3_DFFPOSX1_1014 gnd vdd FILL
XFILL_3_DFFPOSX1_1003 gnd vdd FILL
XFILL_0_INVX4_31 gnd vdd FILL
XFILL_0_INVX4_42 gnd vdd FILL
XFILL_3_DFFPOSX1_1025 gnd vdd FILL
XFILL_6_DFFPOSX1_897 gnd vdd FILL
XXNOR2X1_93 XNOR2X1_93/A INVX2_68/Y gnd XNOR2X1_93/Y vdd XNOR2X1
XXNOR2X1_82 INVX2_106/A bundleAddress_i[28] gnd XNOR2X1_82/Y vdd XNOR2X1
XXNOR2X1_71 XNOR2X1_71/A INVX4_42/Y gnd XNOR2X1_71/Y vdd XNOR2X1
XXNOR2X1_60 INVX1_187/A INVX4_35/Y gnd XNOR2X1_60/Y vdd XNOR2X1
XFILL_0_NAND2X1_401 gnd vdd FILL
XFILL_37_9_1 gnd vdd FILL
XFILL_1_XNOR2X1_5 gnd vdd FILL
XFILL_36_4_0 gnd vdd FILL
XFILL_0_NAND2X1_412 gnd vdd FILL
XFILL_0_NAND2X1_434 gnd vdd FILL
XFILL_1_NAND2X1_605 gnd vdd FILL
XFILL_0_OAI21X1_1205 gnd vdd FILL
XFILL_0_NAND2X1_423 gnd vdd FILL
XBUFX2_70 BUFX2_70/A gnd addr2_o[50] vdd BUFX2
XFILL_0_NAND2X1_478 gnd vdd FILL
XFILL_0_OAI21X1_1227 gnd vdd FILL
XFILL_0_OAI21X1_1216 gnd vdd FILL
XFILL_0_OAI21X1_1238 gnd vdd FILL
XFILL_0_DFFPOSX1_806 gnd vdd FILL
XFILL_0_NAND2X1_445 gnd vdd FILL
XFILL_0_NAND2X1_467 gnd vdd FILL
XFILL_1_NAND2X1_649 gnd vdd FILL
XFILL_1_NAND2X1_627 gnd vdd FILL
XFILL_1_NAND2X1_616 gnd vdd FILL
XBUFX2_81 BUFX2_81/A gnd addr2_o[40] vdd BUFX2
XFILL_0_NAND2X1_456 gnd vdd FILL
XFILL_1_NAND2X1_638 gnd vdd FILL
XBUFX2_92 BUFX2_92/A gnd addr2_o[30] vdd BUFX2
XFILL_0_NAND2X1_489 gnd vdd FILL
XFILL_0_OAI21X1_1249 gnd vdd FILL
XFILL_0_DFFPOSX1_839 gnd vdd FILL
XFILL_0_DFFPOSX1_817 gnd vdd FILL
XFILL_0_DFFPOSX1_828 gnd vdd FILL
XFILL_5_DFFPOSX1_421 gnd vdd FILL
XFILL_5_DFFPOSX1_410 gnd vdd FILL
XFILL_20_8_1 gnd vdd FILL
XFILL_5_DFFPOSX1_443 gnd vdd FILL
XFILL_5_DFFPOSX1_432 gnd vdd FILL
XFILL_5_DFFPOSX1_454 gnd vdd FILL
XFILL_5_DFFPOSX1_476 gnd vdd FILL
XFILL_5_DFFPOSX1_487 gnd vdd FILL
XFILL_5_DFFPOSX1_465 gnd vdd FILL
XFILL_1_BUFX4_70 gnd vdd FILL
XFILL_1_BUFX4_81 gnd vdd FILL
XFILL_5_DFFPOSX1_498 gnd vdd FILL
XFILL_1_BUFX4_92 gnd vdd FILL
XFILL_0_AOI21X1_14 gnd vdd FILL
XFILL_0_AOI21X1_25 gnd vdd FILL
XFILL_0_AOI21X1_36 gnd vdd FILL
XFILL_0_AOI21X1_47 gnd vdd FILL
XFILL_0_OAI21X1_951 gnd vdd FILL
XFILL_2_CLKBUF1_5 gnd vdd FILL
XFILL_0_AOI21X1_58 gnd vdd FILL
XFILL_0_OAI21X1_940 gnd vdd FILL
XFILL_0_OAI21X1_984 gnd vdd FILL
XFILL_0_OAI21X1_962 gnd vdd FILL
XFILL_0_OAI21X1_973 gnd vdd FILL
XFILL_0_OAI21X1_995 gnd vdd FILL
XFILL_28_9_1 gnd vdd FILL
XFILL_3_9_1 gnd vdd FILL
XFILL_27_4_0 gnd vdd FILL
XFILL_2_4_0 gnd vdd FILL
XFILL_2_BUFX4_176 gnd vdd FILL
XFILL_0_OAI21X1_1761 gnd vdd FILL
XFILL_0_OAI21X1_1750 gnd vdd FILL
XFILL_0_OAI21X1_1783 gnd vdd FILL
XFILL_0_OAI21X1_1794 gnd vdd FILL
XFILL_0_OAI21X1_1772 gnd vdd FILL
XFILL_11_8_1 gnd vdd FILL
XFILL_10_3_0 gnd vdd FILL
XFILL_23_10_1 gnd vdd FILL
XFILL_0_NOR2X1_12 gnd vdd FILL
XFILL_0_BUFX2_705 gnd vdd FILL
XFILL_0_NOR2X1_23 gnd vdd FILL
XFILL_0_BUFX2_716 gnd vdd FILL
XFILL_0_BUFX2_727 gnd vdd FILL
XAOI21X1_60 bundleAddress_i[52] INVX2_108/A bundleAddress_i[51] gnd AOI21X1_60/Y vdd
+ AOI21X1
XFILL_0_NOR2X1_56 gnd vdd FILL
XFILL_0_NOR2X1_45 gnd vdd FILL
XFILL_0_BUFX2_749 gnd vdd FILL
XFILL_0_NOR2X1_34 gnd vdd FILL
XFILL_0_BUFX2_738 gnd vdd FILL
XFILL_0_NOR2X1_78 gnd vdd FILL
XFILL_0_NOR2X1_67 gnd vdd FILL
XFILL_0_NOR2X1_89 gnd vdd FILL
XBUFX4_313 BUFX4_380/A gnd BUFX4_313/Y vdd BUFX4
XBUFX4_302 BUFX4_303/A gnd BUFX4_302/Y vdd BUFX4
XFILL_19_9_1 gnd vdd FILL
XBUFX4_346 BUFX4_386/A gnd BUFX4_346/Y vdd BUFX4
XBUFX4_324 BUFX4_378/A gnd BUFX4_324/Y vdd BUFX4
XFILL_0_INVX2_201 gnd vdd FILL
XBUFX4_335 BUFX4_386/A gnd BUFX4_335/Y vdd BUFX4
XBUFX4_368 BUFX4_376/A gnd BUFX4_368/Y vdd BUFX4
XBUFX4_379 BUFX4_385/A gnd OAI21X1_1/A vdd BUFX4
XFILL_18_4_0 gnd vdd FILL
XBUFX4_357 BUFX4_381/A gnd BUFX4_357/Y vdd BUFX4
XFILL_19_4 gnd vdd FILL
XFILL_25_18_0 gnd vdd FILL
XOAI21X1_1203 AOI21X1_45/Y OAI21X1_1203/B NAND2X1_585/Y gnd OAI21X1_1203/Y vdd OAI21X1
XDFFPOSX1_815 BUFX2_126/A CLKBUF1_101/Y OAI21X1_1114/Y gnd vdd DFFPOSX1
XOAI21X1_1214 BUFX4_10/Y BUFX4_353/Y BUFX2_152/A gnd OAI21X1_1215/C vdd OAI21X1
XOAI21X1_1236 BUFX4_251/Y BUFX4_312/Y BUFX2_132/A gnd OAI21X1_1237/C vdd OAI21X1
XOAI21X1_1225 INVX4_47/Y INVX2_60/Y BUFX4_305/Y gnd OAI21X1_1227/A vdd OAI21X1
XOAI21X1_1247 NOR2X1_185/A INVX1_201/A OAI21X1_1247/C gnd OAI21X1_1249/A vdd OAI21X1
XFILL_1_OAI21X1_1401 gnd vdd FILL
XFILL_1_OAI21X1_1423 gnd vdd FILL
XFILL_1_OAI21X1_1412 gnd vdd FILL
XDFFPOSX1_804 BUFX2_58/A CLKBUF1_69/Y OAI21X1_1096/Y gnd vdd DFFPOSX1
XFILL_3_DFFPOSX1_190 gnd vdd FILL
XOAI21X1_1258 NAND2X1_597/Y BUFX4_150/Y OAI21X1_1258/C gnd OAI21X1_1258/Y vdd OAI21X1
XFILL_1_CLKBUF1_70 gnd vdd FILL
XDFFPOSX1_837 BUFX2_87/A CLKBUF1_27/Y OAI21X1_1149/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1434 gnd vdd FILL
XFILL_1_OAI21X1_1456 gnd vdd FILL
XOAI21X1_1269 OR2X2_18/Y NOR3X1_18/C OAI21X1_1269/C gnd OAI21X1_1271/A vdd OAI21X1
XFILL_1_OAI21X1_1445 gnd vdd FILL
XFILL_1_CLKBUF1_81 gnd vdd FILL
XFILL_1_CLKBUF1_92 gnd vdd FILL
XDFFPOSX1_848 BUFX2_100/A CLKBUF1_53/Y OAI21X1_1166/Y gnd vdd DFFPOSX1
XDFFPOSX1_826 BUFX2_75/A CLKBUF1_34/Y OAI21X1_1133/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_203 gnd vdd FILL
XFILL_0_OAI21X1_225 gnd vdd FILL
XFILL_1_OAI21X1_1478 gnd vdd FILL
XFILL_1_OAI21X1_1467 gnd vdd FILL
XFILL_0_OAI21X1_214 gnd vdd FILL
XFILL_0_OAI21X1_236 gnd vdd FILL
XFILL_1_OAI21X1_1489 gnd vdd FILL
XFILL_1_OAI21X1_407 gnd vdd FILL
XFILL_1_OAI21X1_418 gnd vdd FILL
XDFFPOSX1_859 BUFX2_112/A CLKBUF1_76/Y OAI21X1_1183/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_269 gnd vdd FILL
XFILL_0_OAI21X1_247 gnd vdd FILL
XFILL_1_OAI21X1_429 gnd vdd FILL
XFILL_0_OAI21X1_258 gnd vdd FILL
XFILL_6_DFFPOSX1_672 gnd vdd FILL
XFILL_6_DFFPOSX1_650 gnd vdd FILL
XFILL_6_DFFPOSX1_661 gnd vdd FILL
XFILL_6_DFFPOSX1_683 gnd vdd FILL
XFILL_6_DFFPOSX1_694 gnd vdd FILL
XFILL_3_10_1 gnd vdd FILL
XFILL_1_NAND2X1_402 gnd vdd FILL
XFILL_0_NAND2X1_242 gnd vdd FILL
XFILL_0_NAND2X1_220 gnd vdd FILL
XFILL_0_NAND2X1_231 gnd vdd FILL
XFILL_0_OAI21X1_1002 gnd vdd FILL
XFILL_0_OAI21X1_1013 gnd vdd FILL
XFILL_0_NAND2X1_264 gnd vdd FILL
XFILL_0_OAI21X1_1046 gnd vdd FILL
XFILL_1_NAND2X1_435 gnd vdd FILL
XFILL_0_NAND2X1_253 gnd vdd FILL
XFILL_0_NAND2X1_286 gnd vdd FILL
XFILL_0_DFFPOSX1_603 gnd vdd FILL
XFILL_1_NAND2X1_457 gnd vdd FILL
XFILL_0_NAND2X1_275 gnd vdd FILL
XFILL_0_OAI21X1_1024 gnd vdd FILL
XFILL_0_DFFPOSX1_614 gnd vdd FILL
XFILL_0_OAI21X1_1035 gnd vdd FILL
XFILL_0_OAI21X1_1057 gnd vdd FILL
XFILL_0_DFFPOSX1_636 gnd vdd FILL
XFILL_0_OAI21X1_1068 gnd vdd FILL
XFILL_0_OAI21X1_1079 gnd vdd FILL
XFILL_0_NAND2X1_297 gnd vdd FILL
XFILL_0_DFFPOSX1_647 gnd vdd FILL
XFILL_0_DFFPOSX1_625 gnd vdd FILL
XFILL_0_DFFPOSX1_658 gnd vdd FILL
XFILL_0_DFFPOSX1_669 gnd vdd FILL
XFILL_5_DFFPOSX1_262 gnd vdd FILL
XFILL_5_DFFPOSX1_240 gnd vdd FILL
XFILL_5_DFFPOSX1_251 gnd vdd FILL
XFILL_5_DFFPOSX1_273 gnd vdd FILL
XFILL_5_DFFPOSX1_284 gnd vdd FILL
XFILL_5_DFFPOSX1_295 gnd vdd FILL
XOAI21X1_1792 BUFX4_318/Y INVX2_164/Y NAND2X1_733/Y gnd OAI21X1_1792/Y vdd OAI21X1
XOAI21X1_1781 BUFX4_348/Y INVX2_153/Y NAND2X1_722/Y gnd OAI21X1_1781/Y vdd OAI21X1
XOAI21X1_1770 BUFX4_131/Y BUFX4_33/Y BUFX2_769/A gnd OAI21X1_1771/C vdd OAI21X1
XFILL_1_OAI21X1_930 gnd vdd FILL
XFILL_0_OAI21X1_781 gnd vdd FILL
XFILL_2_BUFX4_59 gnd vdd FILL
XFILL_0_OAI21X1_770 gnd vdd FILL
XFILL_1_OAI21X1_952 gnd vdd FILL
XFILL_0_OAI21X1_792 gnd vdd FILL
XFILL_1_OR2X2_4 gnd vdd FILL
XFILL_1_OAI21X1_941 gnd vdd FILL
XFILL_1_OAI21X1_963 gnd vdd FILL
XFILL_1_OAI21X1_985 gnd vdd FILL
XFILL_1_OAI21X1_974 gnd vdd FILL
XFILL_1_OAI21X1_996 gnd vdd FILL
XFILL_5_18_0 gnd vdd FILL
XBUFX2_817 BUFX2_817/A gnd tid1_o[18] vdd BUFX2
XBUFX2_806 BUFX2_806/A gnd tid1_o[28] vdd BUFX2
XBUFX2_828 BUFX2_828/A gnd tid1_o[8] vdd BUFX2
XFILL_2_DFFPOSX1_719 gnd vdd FILL
XFILL_2_DFFPOSX1_708 gnd vdd FILL
XFILL_2_NAND3X1_53 gnd vdd FILL
XBUFX2_839 BUFX2_839/A gnd tid1_o[55] vdd BUFX2
XFILL_0_OAI21X1_1591 gnd vdd FILL
XFILL_0_OAI21X1_1580 gnd vdd FILL
XFILL_1_INVX1_6 gnd vdd FILL
XFILL_0_BUFX2_524 gnd vdd FILL
XFILL_0_BUFX2_513 gnd vdd FILL
XFILL_0_BUFX2_502 gnd vdd FILL
XFILL_1_DFFPOSX1_309 gnd vdd FILL
XFILL_0_BUFX2_546 gnd vdd FILL
XCLKBUF1_5 BUFX4_85/Y gnd CLKBUF1_5/Y vdd CLKBUF1
XFILL_0_BUFX2_557 gnd vdd FILL
XFILL_0_BUFX2_535 gnd vdd FILL
XFILL_0_BUFX2_579 gnd vdd FILL
XFILL_0_BUFX2_568 gnd vdd FILL
XBUFX4_110 BUFX4_10/A gnd BUFX4_110/Y vdd BUFX4
XBUFX4_121 BUFX4_14/Y gnd BUFX4_121/Y vdd BUFX4
XFILL_14_15_1 gnd vdd FILL
XFILL_4_CLKBUF1_25 gnd vdd FILL
XBUFX4_143 BUFX4_18/Y gnd BUFX4_143/Y vdd BUFX4
XBUFX4_132 BUFX4_18/Y gnd BUFX4_132/Y vdd BUFX4
XFILL_4_CLKBUF1_14 gnd vdd FILL
XFILL_0_INVX1_43 gnd vdd FILL
XFILL_0_INVX1_21 gnd vdd FILL
XFILL_0_INVX1_32 gnd vdd FILL
XFILL_0_INVX1_10 gnd vdd FILL
XBUFX4_154 BUFX4_16/Y gnd BUFX4_154/Y vdd BUFX4
XFILL_0_INVX1_65 gnd vdd FILL
XBUFX4_165 BUFX4_14/Y gnd BUFX4_165/Y vdd BUFX4
XFILL_4_CLKBUF1_47 gnd vdd FILL
XNOR2X1_225 INVX2_80/Y NOR2X1_226/B gnd INVX2_110/A vdd NOR2X1
XNOR2X1_203 NOR2X1_204/A NOR2X1_203/B gnd XNOR2X1_85/A vdd NOR2X1
XNOR2X1_214 INVX1_199/Y INVX1_218/Y gnd NOR2X1_214/Y vdd NOR2X1
XBUFX4_187 BUFX4_21/Y gnd BUFX4_187/Y vdd BUFX4
XBUFX4_176 BUFX4_13/Y gnd BUFX4_176/Y vdd BUFX4
XFILL_0_INVX1_76 gnd vdd FILL
XFILL_0_INVX1_54 gnd vdd FILL
XFILL_4_CLKBUF1_58 gnd vdd FILL
XFILL_1_AND2X2_2 gnd vdd FILL
XFILL_34_7_1 gnd vdd FILL
XBUFX4_198 BUFX4_25/Y gnd BUFX4_198/Y vdd BUFX4
XFILL_0_INVX1_98 gnd vdd FILL
XFILL_0_INVX1_87 gnd vdd FILL
XFILL_0_BUFX2_18 gnd vdd FILL
XFILL_33_2_0 gnd vdd FILL
XFILL_24_2 gnd vdd FILL
XFILL_0_BUFX2_29 gnd vdd FILL
XFILL_17_1 gnd vdd FILL
XOAI21X1_709 INVX1_36/A OR2X2_5/A BUFX4_287/Y gnd OAI21X1_711/B vdd OAI21X1
XOAI21X1_1022 BUFX4_136/Y BUFX4_75/Y BUFX2_375/A gnd OAI21X1_1023/C vdd OAI21X1
XOAI21X1_1000 BUFX4_158/Y BUFX4_59/Y BUFX2_363/A gnd OAI21X1_1001/C vdd OAI21X1
XOAI21X1_1011 BUFX4_303/Y INVX1_160/Y OAI21X1_1011/C gnd OAI21X1_1011/Y vdd OAI21X1
XOAI21X1_1033 BUFX4_301/Y INVX1_171/Y OAI21X1_1033/C gnd OAI21X1_1033/Y vdd OAI21X1
XOAI21X1_1044 BUFX4_353/Y INVX2_61/Y NAND2X1_410/Y gnd OAI21X1_1044/Y vdd OAI21X1
XFILL_1_OAI21X1_1231 gnd vdd FILL
XFILL_1_OAI21X1_1220 gnd vdd FILL
XOAI21X1_1055 OAI21X1_5/A INVX4_35/Y NAND2X1_421/Y gnd OAI21X1_1055/Y vdd OAI21X1
XDFFPOSX1_601 BUFX2_634/A CLKBUF1_24/Y OAI21X1_815/Y gnd vdd DFFPOSX1
XDFFPOSX1_612 BUFX2_257/A CLKBUF1_10/Y BUFX4_262/Y gnd vdd DFFPOSX1
XDFFPOSX1_623 INVX1_52/A CLKBUF1_58/Y OAI21X1_851/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_821 gnd vdd FILL
XFILL_1_DFFPOSX1_810 gnd vdd FILL
XDFFPOSX1_645 INVX1_74/A CLKBUF1_96/Y OAI21X1_873/Y gnd vdd DFFPOSX1
XDFFPOSX1_634 INVX1_63/A CLKBUF1_14/Y OAI21X1_862/Y gnd vdd DFFPOSX1
XDFFPOSX1_656 BUFX2_323/A CLKBUF1_39/Y OAI21X1_884/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_832 gnd vdd FILL
XOAI21X1_1066 BUFX4_377/Y INVX2_73/Y NAND2X1_432/Y gnd OAI21X1_1066/Y vdd OAI21X1
XFILL_1_OAI21X1_1253 gnd vdd FILL
XFILL_1_OAI21X1_1242 gnd vdd FILL
XFILL_1_OAI21X1_1264 gnd vdd FILL
XOAI21X1_1088 BUFX4_364/Y INVX2_85/Y NAND2X1_454/Y gnd OAI21X1_1088/Y vdd OAI21X1
XFILL_1_OAI21X1_1275 gnd vdd FILL
XOAI21X1_1077 BUFX4_350/Y INVX4_42/Y NAND2X1_443/Y gnd OAI21X1_1077/Y vdd OAI21X1
XFILL_1_DFFPOSX1_876 gnd vdd FILL
XFILL_1_OAI21X1_1297 gnd vdd FILL
XOAI21X1_1099 BUFX4_360/Y INVX4_46/Y NAND2X1_465/Y gnd OAI21X1_1099/Y vdd OAI21X1
XFILL_1_OAI21X1_1286 gnd vdd FILL
XFILL_1_OAI21X1_215 gnd vdd FILL
XFILL_1_DFFPOSX1_854 gnd vdd FILL
XDFFPOSX1_678 BUFX2_317/A CLKBUF1_51/Y OAI21X1_906/Y gnd vdd DFFPOSX1
XDFFPOSX1_667 BUFX2_304/A CLKBUF1_51/Y OAI21X1_895/Y gnd vdd DFFPOSX1
XDFFPOSX1_689 BUFX2_356/A CLKBUF1_52/Y OAI21X1_927/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_843 gnd vdd FILL
XFILL_1_OAI21X1_226 gnd vdd FILL
XFILL_1_OAI21X1_204 gnd vdd FILL
XFILL_1_DFFPOSX1_865 gnd vdd FILL
XFILL_1_OAI21X1_248 gnd vdd FILL
XNAND2X1_726 BUFX2_780/A BUFX4_363/Y gnd NAND2X1_726/Y vdd NAND2X1
XFILL_1_DFFPOSX1_887 gnd vdd FILL
XNAND2X1_704 BUFX2_696/A BUFX4_223/Y gnd NAND2X1_704/Y vdd NAND2X1
XNAND2X1_715 BUFX2_777/A OAI21X1_1/A gnd NAND2X1_715/Y vdd NAND2X1
XNAND2X1_737 BUFX2_792/A BUFX4_375/Y gnd NAND2X1_737/Y vdd NAND2X1
XFILL_1_DFFPOSX1_898 gnd vdd FILL
XFILL_19_14_1 gnd vdd FILL
XFILL_1_OAI21X1_259 gnd vdd FILL
XFILL_1_OAI21X1_237 gnd vdd FILL
XFILL_0_NOR2X1_9 gnd vdd FILL
XNAND2X1_748 BUFX2_804/A BUFX4_329/Y gnd NAND2X1_748/Y vdd NAND2X1
XNAND2X1_759 BUFX2_816/A BUFX4_336/Y gnd NAND2X1_759/Y vdd NAND2X1
XFILL_32_16_1 gnd vdd FILL
XFILL_13_10_0 gnd vdd FILL
XFILL_25_7_1 gnd vdd FILL
XFILL_1_NAND2X1_210 gnd vdd FILL
XFILL_1_NAND2X1_221 gnd vdd FILL
XFILL_0_7_1 gnd vdd FILL
XFILL_1_NAND2X1_265 gnd vdd FILL
XFILL_24_2_0 gnd vdd FILL
XFILL_1_NAND2X1_243 gnd vdd FILL
XFILL_0_DFFPOSX1_422 gnd vdd FILL
XFILL_0_DFFPOSX1_400 gnd vdd FILL
XFILL_0_DFFPOSX1_433 gnd vdd FILL
XFILL_0_DFFPOSX1_411 gnd vdd FILL
XFILL_2_DFFPOSX1_8 gnd vdd FILL
XFILL_1_NAND2X1_298 gnd vdd FILL
XFILL_0_DFFPOSX1_466 gnd vdd FILL
XFILL_0_DFFPOSX1_455 gnd vdd FILL
XFILL_0_DFFPOSX1_444 gnd vdd FILL
XINVX8_7 bundleLen_i[1] gnd INVX8_7/Y vdd INVX8
XFILL_0_DFFPOSX1_477 gnd vdd FILL
XFILL_0_DFFPOSX1_499 gnd vdd FILL
XFILL_0_DFFPOSX1_488 gnd vdd FILL
XFILL_3_DFFPOSX1_904 gnd vdd FILL
XFILL_3_DFFPOSX1_948 gnd vdd FILL
XFILL_3_DFFPOSX1_937 gnd vdd FILL
XFILL_3_DFFPOSX1_915 gnd vdd FILL
XFILL_3_DFFPOSX1_926 gnd vdd FILL
XFILL_3_DFFPOSX1_959 gnd vdd FILL
XDFFPOSX1_60 BUFX2_730/A CLKBUF1_47/Y DFFPOSX1_60/D gnd vdd DFFPOSX1
XDFFPOSX1_71 BUFX2_768/A CLKBUF1_35/Y DFFPOSX1_71/D gnd vdd DFFPOSX1
XDFFPOSX1_82 BUFX2_751/A CLKBUF1_86/Y DFFPOSX1_82/D gnd vdd DFFPOSX1
XDFFPOSX1_93 BUFX2_763/A CLKBUF1_50/Y DFFPOSX1_93/D gnd vdd DFFPOSX1
XFILL_37_15_1 gnd vdd FILL
XFILL_8_8_1 gnd vdd FILL
XFILL_1_OAI21X1_782 gnd vdd FILL
XFILL_1_OAI21X1_771 gnd vdd FILL
XFILL_1_OAI21X1_760 gnd vdd FILL
XBUFX4_16 INVX8_6/Y gnd BUFX4_16/Y vdd BUFX4
XFILL_7_3_0 gnd vdd FILL
XFILL_2_OAI21X1_975 gnd vdd FILL
XBUFX4_38 BUFX4_51/A gnd BUFX4_38/Y vdd BUFX4
XBUFX4_49 BUFX4_81/A gnd BUFX4_49/Y vdd BUFX4
XFILL_1_OAI21X1_793 gnd vdd FILL
XBUFX4_27 BUFX4_79/A gnd BUFX4_27/Y vdd BUFX4
XFILL_2_OAI21X1_964 gnd vdd FILL
XFILL_31_11_0 gnd vdd FILL
XBUFX2_603 BUFX2_603/A gnd majID4_o[38] vdd BUFX2
XFILL_2_DFFPOSX1_505 gnd vdd FILL
XBUFX2_614 BUFX2_614/A gnd majID4_o[28] vdd BUFX2
XFILL_2_DFFPOSX1_516 gnd vdd FILL
XFILL_2_DFFPOSX1_527 gnd vdd FILL
XFILL_2_DFFPOSX1_538 gnd vdd FILL
XBUFX2_636 BUFX2_636/A gnd majID4_o[8] vdd BUFX2
XBUFX2_625 BUFX2_625/A gnd majID4_o[18] vdd BUFX2
XBUFX2_658 BUFX2_658/A gnd pid1_o[14] vdd BUFX2
XBUFX2_669 BUFX2_669/A gnd pid1_o[4] vdd BUFX2
XFILL_16_7_1 gnd vdd FILL
XBUFX2_647 BUFX2_647/A gnd majID4_o[55] vdd BUFX2
XFILL_2_DFFPOSX1_549 gnd vdd FILL
XFILL_15_2_0 gnd vdd FILL
XFILL_0_BUFX2_310 gnd vdd FILL
XINVX2_132 bundlePid_i[16] gnd INVX2_132/Y vdd INVX2
XFILL_0_BUFX2_321 gnd vdd FILL
XOR2X2_19 OR2X2_19/A OR2X2_19/B gnd OR2X2_19/Y vdd OR2X2
XINVX2_110 INVX2_110/A gnd INVX2_110/Y vdd INVX2
XFILL_0_BUFX2_332 gnd vdd FILL
XINVX2_121 bundlePid_i[27] gnd INVX2_121/Y vdd INVX2
XINVX2_165 bundleTid_i[44] gnd INVX2_165/Y vdd INVX2
XFILL_1_DFFPOSX1_117 gnd vdd FILL
XINVX2_143 bundlePid_i[5] gnd INVX2_143/Y vdd INVX2
XFILL_1_DFFPOSX1_106 gnd vdd FILL
XFILL_0_BUFX2_354 gnd vdd FILL
XINVX2_154 bundleTid_i[55] gnd INVX2_154/Y vdd INVX2
XFILL_1_DFFPOSX1_128 gnd vdd FILL
XFILL_0_BUFX2_365 gnd vdd FILL
XFILL_0_BUFX2_343 gnd vdd FILL
XINVX2_176 bundleTid_i[33] gnd INVX2_176/Y vdd INVX2
XFILL_1_DFFPOSX1_139 gnd vdd FILL
XINVX2_187 bundleTid_i[22] gnd INVX2_187/Y vdd INVX2
XFILL_0_BUFX2_376 gnd vdd FILL
XINVX2_198 bundleTid_i[11] gnd INVX2_198/Y vdd INVX2
XFILL_0_BUFX2_387 gnd vdd FILL
XFILL_0_BUFX2_398 gnd vdd FILL
XFILL_36_10_0 gnd vdd FILL
XOAI21X1_506 INVX1_24/Y bundleStartMajId_i[60] NOR2X1_89/B gnd OAI21X1_508/B vdd OAI21X1
XOAI21X1_539 OAI22X1_1/B INVX1_26/Y NOR2X1_9/A gnd OAI21X1_539/Y vdd OAI21X1
XOAI21X1_528 OR2X2_1/A INVX4_30/Y OAI21X1_528/C gnd OAI21X1_530/A vdd OAI21X1
XOAI21X1_517 XNOR2X1_24/Y BUFX4_163/Y OAI21X1_517/C gnd OAI21X1_517/Y vdd OAI21X1
XFILL_1_OAI21X1_1050 gnd vdd FILL
XFILL_1_NAND3X1_50 gnd vdd FILL
XFILL_1_NAND3X1_61 gnd vdd FILL
XDFFPOSX1_431 BUFX2_460/A CLKBUF1_75/Y OAI21X1_416/Y gnd vdd DFFPOSX1
XDFFPOSX1_420 BUFX2_457/A CLKBUF1_10/Y OAI21X1_392/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_640 gnd vdd FILL
XFILL_1_OAI21X1_1083 gnd vdd FILL
XFILL_1_DFFPOSX1_651 gnd vdd FILL
XFILL_1_OAI21X1_1061 gnd vdd FILL
XDFFPOSX1_442 BUFX2_472/A CLKBUF1_18/Y OAI21X1_433/Y gnd vdd DFFPOSX1
XDFFPOSX1_453 BUFX2_484/A CLKBUF1_44/Y OAI21X1_450/Y gnd vdd DFFPOSX1
XDFFPOSX1_464 BUFX2_496/A CLKBUF1_48/Y OAI21X1_466/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1072 gnd vdd FILL
XFILL_1_DFFPOSX1_662 gnd vdd FILL
XNAND2X1_501 NOR2X1_130/Y NOR2X1_133/Y gnd NOR2X1_220/A vdd NAND2X1
XFILL_1_OAI21X1_1094 gnd vdd FILL
XDFFPOSX1_486 BUFX2_533/A CLKBUF1_45/Y OAI21X1_505/Y gnd vdd DFFPOSX1
XNAND2X1_512 bundleAddress_i[45] bundleAddress_i[42] gnd NOR2X1_140/B vdd NAND2X1
XDFFPOSX1_497 BUFX2_526/A CLKBUF1_46/Y OAI21X1_538/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_673 gnd vdd FILL
XFILL_1_DFFPOSX1_684 gnd vdd FILL
XDFFPOSX1_475 BUFX2_508/A CLKBUF1_48/Y OAI21X1_485/Y gnd vdd DFFPOSX1
XNAND2X1_523 bundleAddress_i[37] bundleAddress_i[36] gnd NOR2X1_144/A vdd NAND2X1
XFILL_1_DFFPOSX1_695 gnd vdd FILL
XNAND2X1_534 BUFX2_93/A INVX8_1/A gnd NAND2X1_534/Y vdd NAND2X1
XFILL_2_OAI21X1_227 gnd vdd FILL
XNAND2X1_545 BUFX2_100/A BUFX4_226/Y gnd NAND2X1_545/Y vdd NAND2X1
XNAND2X1_556 bundleAddress_i[21] bundleAddress_i[18] gnd NOR2X1_163/B vdd NAND2X1
XNAND2X1_567 BUFX2_111/A INVX8_1/A gnd NAND2X1_567/Y vdd NAND2X1
XNAND2X1_578 BUFX2_117/A BUFX4_188/Y gnd NAND2X1_578/Y vdd NAND2X1
XNAND2X1_589 BUFX2_125/A BUFX4_187/Y gnd NAND2X1_589/Y vdd NAND2X1
XFILL_0_AND2X2_24 gnd vdd FILL
XFILL_0_AND2X2_13 gnd vdd FILL
XFILL_0_DFFPOSX1_230 gnd vdd FILL
XFILL_0_DFFPOSX1_241 gnd vdd FILL
XFILL_0_DFFPOSX1_252 gnd vdd FILL
XFILL_0_DFFPOSX1_263 gnd vdd FILL
XFILL_0_DFFPOSX1_274 gnd vdd FILL
XFILL_0_DFFPOSX1_296 gnd vdd FILL
XFILL_0_DFFPOSX1_285 gnd vdd FILL
XFILL_3_DFFPOSX1_701 gnd vdd FILL
XFILL_3_DFFPOSX1_712 gnd vdd FILL
XFILL_3_DFFPOSX1_723 gnd vdd FILL
XFILL_3_DFFPOSX1_756 gnd vdd FILL
XFILL_3_CLKBUF1_11 gnd vdd FILL
XFILL_3_CLKBUF1_22 gnd vdd FILL
XFILL_3_DFFPOSX1_745 gnd vdd FILL
XFILL_3_DFFPOSX1_734 gnd vdd FILL
XFILL_3_CLKBUF1_33 gnd vdd FILL
XFILL_3_DFFPOSX1_789 gnd vdd FILL
XFILL_3_CLKBUF1_55 gnd vdd FILL
XFILL_3_DFFPOSX1_778 gnd vdd FILL
XFILL_3_CLKBUF1_44 gnd vdd FILL
XFILL_3_DFFPOSX1_767 gnd vdd FILL
XFILL_3_CLKBUF1_66 gnd vdd FILL
XFILL_3_CLKBUF1_99 gnd vdd FILL
XFILL_3_CLKBUF1_88 gnd vdd FILL
XFILL_3_CLKBUF1_77 gnd vdd FILL
XFILL_1_NOR2X1_140 gnd vdd FILL
XFILL_1_NOR2X1_151 gnd vdd FILL
XFILL_1_NOR2X1_162 gnd vdd FILL
XFILL_1_OAI21X1_590 gnd vdd FILL
XFILL_1_NOR2X1_195 gnd vdd FILL
XFILL_2_OAI21X1_783 gnd vdd FILL
XFILL_2_DFFPOSX1_313 gnd vdd FILL
XBUFX2_411 BUFX2_411/A gnd majID1_o[38] vdd BUFX2
XFILL_2_DFFPOSX1_302 gnd vdd FILL
XBUFX2_400 BUFX2_400/A gnd majID1_o[48] vdd BUFX2
XFILL_2_DFFPOSX1_346 gnd vdd FILL
XFILL_2_DFFPOSX1_335 gnd vdd FILL
XBUFX2_433 BUFX2_433/A gnd majID1_o[18] vdd BUFX2
XBUFX2_422 BUFX2_422/A gnd majID1_o[28] vdd BUFX2
XBUFX2_444 BUFX2_444/A gnd majID1_o[8] vdd BUFX2
XFILL_2_DFFPOSX1_324 gnd vdd FILL
XBUFX2_488 BUFX2_488/A gnd majID2_o[26] vdd BUFX2
XFILL_2_DFFPOSX1_357 gnd vdd FILL
XFILL_2_DFFPOSX1_368 gnd vdd FILL
XBUFX2_466 BUFX2_466/A gnd majID2_o[46] vdd BUFX2
XBUFX2_455 BUFX2_455/A gnd majID1_o[55] vdd BUFX2
XFILL_2_DFFPOSX1_379 gnd vdd FILL
XBUFX2_477 BUFX2_477/A gnd majID2_o[36] vdd BUFX2
XBUFX2_499 BUFX2_499/A gnd majID2_o[16] vdd BUFX2
XFILL_31_5_1 gnd vdd FILL
XFILL_5_DFFPOSX1_806 gnd vdd FILL
XFILL_5_DFFPOSX1_817 gnd vdd FILL
XFILL_5_DFFPOSX1_828 gnd vdd FILL
XFILL_1_BUFX4_382 gnd vdd FILL
XFILL_30_0_0 gnd vdd FILL
XFILL_5_DFFPOSX1_839 gnd vdd FILL
XFILL_1_BUFX4_360 gnd vdd FILL
XFILL_1_BUFX4_371 gnd vdd FILL
XFILL_1_XNOR2X1_18 gnd vdd FILL
XFILL_22_16_0 gnd vdd FILL
XFILL_1_XNOR2X1_29 gnd vdd FILL
XFILL_2_OAI21X1_84 gnd vdd FILL
XFILL_0_BUFX2_140 gnd vdd FILL
XFILL_0_BUFX2_151 gnd vdd FILL
XFILL_0_BUFX2_173 gnd vdd FILL
XFILL_0_BUFX2_162 gnd vdd FILL
XFILL_0_BUFX2_195 gnd vdd FILL
XFILL_0_BUFX2_184 gnd vdd FILL
XFILL_1_DFFPOSX1_5 gnd vdd FILL
XFILL_4_DFFPOSX1_418 gnd vdd FILL
XFILL_4_DFFPOSX1_407 gnd vdd FILL
XFILL_4_DFFPOSX1_429 gnd vdd FILL
XFILL_38_1_0 gnd vdd FILL
XFILL_2_DFFPOSX1_880 gnd vdd FILL
XFILL_2_DFFPOSX1_891 gnd vdd FILL
XFILL_22_5_1 gnd vdd FILL
XFILL_27_15_0 gnd vdd FILL
XOAI21X1_314 BUFX4_147/Y BUFX4_31/Y BUFX2_1022/A gnd OAI21X1_315/C vdd OAI21X1
XFILL_21_0_0 gnd vdd FILL
XOAI21X1_303 INVX2_197/Y BUFX4_303/Y OAI21X1_303/C gnd OAI21X1_303/Y vdd OAI21X1
XOAI21X1_347 BUFX4_319/Y OR2X2_5/B NAND2X1_91/Y gnd OAI21X1_347/Y vdd OAI21X1
XOAI21X1_325 INVX2_6/Y BUFX4_302/Y OAI21X1_325/C gnd OAI21X1_325/Y vdd OAI21X1
XOAI21X1_336 BUFX4_387/Y NOR2X1_5/A NAND2X1_80/Y gnd OAI21X1_336/Y vdd OAI21X1
XOAI21X1_369 BUFX4_362/Y INVX4_20/Y OAI21X1_369/C gnd OAI21X1_369/Y vdd OAI21X1
XOAI21X1_358 BUFX4_314/Y NOR3X1_7/A OAI21X1_358/C gnd OAI21X1_358/Y vdd OAI21X1
XBUFX4_1 BUFX4_1/A gnd BUFX4_1/Y vdd BUFX4
XDFFPOSX1_261 BUFX2_932/A CLKBUF1_39/Y OAI21X1_139/Y gnd vdd DFFPOSX1
XDFFPOSX1_272 BUFX2_944/A CLKBUF1_3/Y OAI21X1_161/Y gnd vdd DFFPOSX1
XDFFPOSX1_250 BUFX2_920/A CLKBUF1_97/Y OAI21X1_117/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_470 gnd vdd FILL
XFILL_1_DFFPOSX1_481 gnd vdd FILL
XDFFPOSX1_283 BUFX2_956/A CLKBUF1_87/Y OAI21X1_183/Y gnd vdd DFFPOSX1
XNAND2X1_320 OAI21X1_727/Y INVX1_38/Y gnd OAI21X1_729/A vdd NAND2X1
XDFFPOSX1_294 BUFX2_981/A CLKBUF1_92/Y OAI21X1_205/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_492 gnd vdd FILL
XNAND2X1_331 OAI21X1_797/Y INVX2_53/Y gnd OAI21X1_799/A vdd NAND2X1
XFILL_3_NOR3X1_14 gnd vdd FILL
XNAND2X1_342 BUFX4_268/Y bundle_i[27] gnd OAI21X1_848/C vdd NAND2X1
XNAND2X1_353 BUFX4_262/Y bundle_i[16] gnd OAI21X1_859/C vdd NAND2X1
XNAND2X1_386 BUFX2_301/A BUFX4_184/Y gnd OAI21X1_892/C vdd NAND2X1
XNAND2X1_375 BUFX2_320/A BUFX4_206/Y gnd OAI21X1_881/C vdd NAND2X1
XFILL_4_DFFPOSX1_941 gnd vdd FILL
XNAND2X1_364 BUFX4_261/Y bundle_i[5] gnd OAI21X1_870/C vdd NAND2X1
XFILL_4_DFFPOSX1_930 gnd vdd FILL
XFILL_5_6_1 gnd vdd FILL
XFILL_4_DFFPOSX1_952 gnd vdd FILL
XFILL_29_1_0 gnd vdd FILL
XFILL_4_DFFPOSX1_963 gnd vdd FILL
XNAND2X1_397 BUFX2_313/A BUFX4_181/Y gnd OAI21X1_903/C vdd NAND2X1
XFILL_4_1_0 gnd vdd FILL
XFILL_4_DFFPOSX1_974 gnd vdd FILL
XFILL_4_DFFPOSX1_985 gnd vdd FILL
XFILL_4_DFFPOSX1_996 gnd vdd FILL
XFILL_0_INVX1_107 gnd vdd FILL
XFILL_0_INVX1_118 gnd vdd FILL
XFILL_2_16_0 gnd vdd FILL
XFILL_0_INVX1_129 gnd vdd FILL
XFILL_1_AOI21X1_18 gnd vdd FILL
XFILL_1_AOI21X1_29 gnd vdd FILL
XFILL_13_5_1 gnd vdd FILL
XINVX4_1 bundleStartMajId_i[63] gnd INVX4_1/Y vdd INVX4
XFILL_12_0_0 gnd vdd FILL
XFILL_1_BUFX2_842 gnd vdd FILL
XFILL_1_BUFX2_853 gnd vdd FILL
XFILL_1_BUFX2_864 gnd vdd FILL
XFILL_1_BUFX2_897 gnd vdd FILL
XFILL_2_NOR3X1_6 gnd vdd FILL
XFILL_3_DFFPOSX1_520 gnd vdd FILL
XFILL_3_DFFPOSX1_531 gnd vdd FILL
XFILL_1_BUFX2_886 gnd vdd FILL
XFILL_1_OAI21X1_1808 gnd vdd FILL
XFILL_1_OAI21X1_1819 gnd vdd FILL
XOAI21X1_892 INVX1_93/Y BUFX4_184/Y OAI21X1_892/C gnd OAI21X1_892/Y vdd OAI21X1
XFILL_3_DFFPOSX1_542 gnd vdd FILL
XOAI21X1_881 INVX1_82/Y BUFX4_206/Y OAI21X1_881/C gnd OAI21X1_881/Y vdd OAI21X1
XOAI21X1_870 INVX1_71/Y BUFX4_261/Y OAI21X1_870/C gnd OAI21X1_870/Y vdd OAI21X1
XFILL_3_DFFPOSX1_564 gnd vdd FILL
XFILL_3_DFFPOSX1_553 gnd vdd FILL
XFILL_3_DFFPOSX1_575 gnd vdd FILL
XFILL_3_DFFPOSX1_586 gnd vdd FILL
XFILL_3_DFFPOSX1_597 gnd vdd FILL
XFILL_7_15_0 gnd vdd FILL
XFILL_2_DFFPOSX1_121 gnd vdd FILL
XFILL_0_NAND2X1_605 gnd vdd FILL
XFILL_0_NAND2X1_627 gnd vdd FILL
XFILL_0_NAND2X1_616 gnd vdd FILL
XFILL_2_DFFPOSX1_110 gnd vdd FILL
XFILL_2_DFFPOSX1_154 gnd vdd FILL
XFILL_2_DFFPOSX1_143 gnd vdd FILL
XFILL_0_OAI21X1_1409 gnd vdd FILL
XBUFX2_252 BUFX2_252/A gnd addr4_o[1] vdd BUFX2
XFILL_0_NAND2X1_649 gnd vdd FILL
XBUFX2_230 BUFX2_230/A gnd addr4_o[21] vdd BUFX2
XFILL_11_13_1 gnd vdd FILL
XBUFX2_241 BUFX2_241/A gnd addr4_o[11] vdd BUFX2
XFILL_2_DFFPOSX1_132 gnd vdd FILL
XFILL_0_NAND2X1_638 gnd vdd FILL
XFILL_2_DFFPOSX1_198 gnd vdd FILL
XBUFX2_274 INVX1_65/A gnd instr1_o[11] vdd BUFX2
XFILL_2_DFFPOSX1_176 gnd vdd FILL
XFILL_2_DFFPOSX1_187 gnd vdd FILL
XBUFX2_285 INVX1_75/A gnd instr1_o[1] vdd BUFX2
XBUFX2_296 BUFX2_296/A gnd instr2_o[20] vdd BUFX2
XBUFX2_263 INVX1_55/A gnd instr1_o[21] vdd BUFX2
XFILL_2_DFFPOSX1_165 gnd vdd FILL
XFILL_5_DFFPOSX1_603 gnd vdd FILL
XFILL_5_DFFPOSX1_636 gnd vdd FILL
XFILL_5_DFFPOSX1_625 gnd vdd FILL
XFILL_5_DFFPOSX1_614 gnd vdd FILL
XFILL_5_DFFPOSX1_647 gnd vdd FILL
XFILL_1_BUFX4_190 gnd vdd FILL
XFILL_5_DFFPOSX1_658 gnd vdd FILL
XFILL_5_DFFPOSX1_669 gnd vdd FILL
XNAND3X1_4 AND2X2_4/Y AND2X2_5/Y NOR2X1_27/Y gnd NOR2X1_30/A vdd NAND3X1
XFILL_4_DFFPOSX1_215 gnd vdd FILL
XFILL_16_12_1 gnd vdd FILL
XFILL_4_DFFPOSX1_226 gnd vdd FILL
XFILL_4_DFFPOSX1_204 gnd vdd FILL
XFILL_4_DFFPOSX1_237 gnd vdd FILL
XFILL_4_DFFPOSX1_248 gnd vdd FILL
XFILL_4_DFFPOSX1_259 gnd vdd FILL
XFILL_2_CLKBUF1_30 gnd vdd FILL
XFILL_2_CLKBUF1_41 gnd vdd FILL
XFILL_2_CLKBUF1_74 gnd vdd FILL
XFILL_2_CLKBUF1_63 gnd vdd FILL
XFILL_2_CLKBUF1_52 gnd vdd FILL
XFILL_2_CLKBUF1_96 gnd vdd FILL
XFILL_2_CLKBUF1_85 gnd vdd FILL
XFILL_2_BUFX4_369 gnd vdd FILL
XOAI21X1_100 BUFX4_11/A BUFX4_341/Y BUFX2_911/A gnd OAI21X1_101/C vdd OAI21X1
XFILL_1_BUFX2_138 gnd vdd FILL
XFILL_1_BUFX2_127 gnd vdd FILL
XFILL_0_NOR2X1_181 gnd vdd FILL
XOAI21X1_111 BUFX4_127/Y INVX2_165/Y OAI21X1_111/C gnd OAI21X1_111/Y vdd OAI21X1
XFILL_1_BUFX2_149 gnd vdd FILL
XOAI21X1_122 BUFX4_4/A BUFX4_317/Y BUFX2_923/A gnd OAI21X1_123/C vdd OAI21X1
XFILL_0_NOR2X1_170 gnd vdd FILL
XFILL_0_DFFPOSX1_1011 gnd vdd FILL
XOAI21X1_133 BUFX4_149/Y INVX2_176/Y OAI21X1_133/C gnd OAI21X1_133/Y vdd OAI21X1
XFILL_0_DFFPOSX1_1000 gnd vdd FILL
XFILL_0_NOR2X1_192 gnd vdd FILL
XOAI21X1_144 BUFX4_5/Y BUFX4_317/Y BUFX2_935/A gnd OAI21X1_145/C vdd OAI21X1
XOAI21X1_155 BUFX4_139/Y INVX2_187/Y OAI21X1_155/C gnd OAI21X1_155/Y vdd OAI21X1
XFILL_0_BUFX2_909 gnd vdd FILL
XOAI21X1_166 BUFX4_104/Y BUFX4_361/Y BUFX2_947/A gnd OAI21X1_167/C vdd OAI21X1
XFILL_0_DFFPOSX1_1022 gnd vdd FILL
XINVX1_208 INVX1_208/A gnd INVX1_208/Y vdd INVX1
XOAI21X1_188 BUFX4_4/A BUFX4_354/Y BUFX2_959/A gnd OAI21X1_189/C vdd OAI21X1
XOAI21X1_177 BUFX4_130/Y INVX2_198/Y OAI21X1_177/C gnd OAI21X1_177/Y vdd OAI21X1
XINVX1_219 INVX1_219/A gnd INVX1_219/Y vdd INVX1
XOAI21X1_199 BUFX4_144/Y INVX2_7/Y OAI21X1_199/C gnd OAI21X1_199/Y vdd OAI21X1
XNAND2X1_19 BUFX2_844/A BUFX4_220/Y gnd OAI21X1_19/C vdd NAND2X1
XFILL_34_13_1 gnd vdd FILL
XNAND2X1_150 NOR2X1_3/Y NOR2X1_4/Y gnd NOR2X1_5/B vdd NAND2X1
XNAND2X1_161 BUFX2_462/A BUFX4_225/Y gnd OAI21X1_420/C vdd NAND2X1
XFILL_0_XNOR2X1_15 gnd vdd FILL
XNAND2X1_172 BUFX4_245/Y OAI21X1_426/Y gnd OAI21X1_427/A vdd NAND2X1
XFILL_0_XNOR2X1_26 gnd vdd FILL
XNAND2X1_194 bundleStartMajId_i[36] bundleStartMajId_i[35] gnd NOR2X1_19/B vdd NAND2X1
XNAND2X1_183 BUFX2_472/A BUFX4_194/Y gnd OAI21X1_433/C vdd NAND2X1
XFILL_0_XNOR2X1_59 gnd vdd FILL
XFILL_4_DFFPOSX1_771 gnd vdd FILL
XFILL_4_DFFPOSX1_760 gnd vdd FILL
XFILL_0_XNOR2X1_37 gnd vdd FILL
XFILL_0_XNOR2X1_48 gnd vdd FILL
XFILL_1_OAI21X1_70 gnd vdd FILL
XFILL_4_DFFPOSX1_782 gnd vdd FILL
XFILL_1_OAI21X1_81 gnd vdd FILL
XFILL_4_DFFPOSX1_793 gnd vdd FILL
XFILL_1_OAI21X1_92 gnd vdd FILL
XFILL_0_DFFPOSX1_2 gnd vdd FILL
XFILL_1_BUFX2_650 gnd vdd FILL
XFILL_1_BUFX2_661 gnd vdd FILL
XFILL_0_BUFX4_202 gnd vdd FILL
XFILL_0_BUFX4_224 gnd vdd FILL
XFILL_0_BUFX4_213 gnd vdd FILL
XFILL_0_BUFX4_235 gnd vdd FILL
XFILL_0_BUFX4_246 gnd vdd FILL
XOAI21X1_1418 INVX2_108/Y INVX2_96/A BUFX4_288/Y gnd OAI21X1_1420/A vdd OAI21X1
XFILL_0_BUFX4_257 gnd vdd FILL
XOAI21X1_1407 BUFX4_179/Y BUFX4_75/Y BUFX2_255/A gnd OAI21X1_1408/C vdd OAI21X1
XOAI21X1_1429 XNOR2X1_92/Y BUFX4_291/Y OAI21X1_1429/C gnd OAI21X1_1429/Y vdd OAI21X1
XFILL_1_BUFX2_694 gnd vdd FILL
XFILL_1_OAI21X1_1605 gnd vdd FILL
XFILL_1_OAI21X1_1649 gnd vdd FILL
XFILL_1_OAI21X1_1616 gnd vdd FILL
XFILL_0_BUFX4_279 gnd vdd FILL
XFILL_1_OAI21X1_1627 gnd vdd FILL
XNOR3X1_7 NOR3X1_7/A bundleStartMajId_i[32] NOR3X1_7/C gnd NOR3X1_7/Y vdd NOR3X1
XFILL_0_BUFX4_268 gnd vdd FILL
XFILL_3_DFFPOSX1_350 gnd vdd FILL
XFILL_1_OAI21X1_1638 gnd vdd FILL
XFILL_3_DFFPOSX1_361 gnd vdd FILL
XFILL_3_DFFPOSX1_372 gnd vdd FILL
XFILL_3_DFFPOSX1_394 gnd vdd FILL
XFILL_0_OAI21X1_429 gnd vdd FILL
XFILL_0_OAI21X1_407 gnd vdd FILL
XFILL_0_OAI21X1_418 gnd vdd FILL
XFILL_3_DFFPOSX1_383 gnd vdd FILL
XFILL_0_INVX4_21 gnd vdd FILL
XFILL_0_INVX4_10 gnd vdd FILL
XFILL_3_DFFPOSX1_1004 gnd vdd FILL
XFILL_6_DFFPOSX1_832 gnd vdd FILL
XFILL_0_INVX4_32 gnd vdd FILL
XFILL_3_DFFPOSX1_1015 gnd vdd FILL
XFILL_6_DFFPOSX1_854 gnd vdd FILL
XFILL_0_INVX4_43 gnd vdd FILL
XFILL_6_DFFPOSX1_843 gnd vdd FILL
XFILL_5_1 gnd vdd FILL
XFILL_6_DFFPOSX1_887 gnd vdd FILL
XFILL_6_DFFPOSX1_876 gnd vdd FILL
XFILL_3_DFFPOSX1_1026 gnd vdd FILL
XXNOR2X1_50 XNOR2X1_50/A bundleStartMajId_i[26] gnd XNOR2X1_50/Y vdd XNOR2X1
XFILL_6_DFFPOSX1_865 gnd vdd FILL
XXNOR2X1_72 INVX1_194/A INVX4_43/Y gnd XNOR2X1_72/Y vdd XNOR2X1
XXNOR2X1_83 XNOR2X1_83/A INVX4_41/Y gnd XNOR2X1_83/Y vdd XNOR2X1
XXNOR2X1_61 XNOR2X1_61/A bundleAddress_i[40] gnd XNOR2X1_61/Y vdd XNOR2X1
XXNOR2X1_94 INVX1_222/A OR2X2_18/B gnd XNOR2X1_94/Y vdd XNOR2X1
XFILL_36_4_1 gnd vdd FILL
XFILL_0_NAND2X1_402 gnd vdd FILL
XFILL_0_NAND2X1_413 gnd vdd FILL
XFILL_0_NAND2X1_435 gnd vdd FILL
XFILL_0_OAI21X1_1206 gnd vdd FILL
XFILL_0_NAND2X1_424 gnd vdd FILL
XFILL_1_XNOR2X1_6 gnd vdd FILL
XFILL_0_NAND2X1_468 gnd vdd FILL
XBUFX2_71 BUFX2_71/A gnd addr2_o[49] vdd BUFX2
XFILL_0_OAI21X1_1228 gnd vdd FILL
XFILL_0_OAI21X1_1217 gnd vdd FILL
XFILL_0_OAI21X1_1239 gnd vdd FILL
XFILL_0_NAND2X1_446 gnd vdd FILL
XBUFX2_60 BUFX2_60/A gnd addr1_o[1] vdd BUFX2
XFILL_0_DFFPOSX1_807 gnd vdd FILL
XFILL_1_NAND2X1_617 gnd vdd FILL
XFILL_0_NAND2X1_457 gnd vdd FILL
XBUFX2_82 BUFX2_82/A gnd addr2_o[39] vdd BUFX2
XFILL_0_NAND2X1_479 gnd vdd FILL
XFILL_0_DFFPOSX1_818 gnd vdd FILL
XBUFX2_93 BUFX2_93/A gnd addr2_o[29] vdd BUFX2
XFILL_0_DFFPOSX1_829 gnd vdd FILL
XFILL_5_DFFPOSX1_400 gnd vdd FILL
XFILL_5_DFFPOSX1_411 gnd vdd FILL
XFILL_5_DFFPOSX1_422 gnd vdd FILL
XFILL_5_DFFPOSX1_433 gnd vdd FILL
XFILL_5_DFFPOSX1_444 gnd vdd FILL
XFILL_5_DFFPOSX1_477 gnd vdd FILL
XFILL_5_DFFPOSX1_466 gnd vdd FILL
XFILL_5_DFFPOSX1_488 gnd vdd FILL
XFILL_5_DFFPOSX1_455 gnd vdd FILL
XFILL_1_BUFX4_60 gnd vdd FILL
XFILL_1_BUFX4_71 gnd vdd FILL
XFILL_5_DFFPOSX1_499 gnd vdd FILL
XFILL_1_BUFX4_82 gnd vdd FILL
XFILL_1_BUFX4_93 gnd vdd FILL
XFILL_0_AOI21X1_26 gnd vdd FILL
XFILL_0_AOI21X1_37 gnd vdd FILL
XFILL_0_AOI21X1_48 gnd vdd FILL
XFILL_0_AOI21X1_15 gnd vdd FILL
XFILL_0_OAI21X1_930 gnd vdd FILL
XFILL_0_AOI21X1_59 gnd vdd FILL
XFILL_0_OAI21X1_941 gnd vdd FILL
XFILL_2_CLKBUF1_6 gnd vdd FILL
XFILL_0_OAI21X1_974 gnd vdd FILL
XFILL_0_OAI21X1_952 gnd vdd FILL
XFILL_0_OAI21X1_963 gnd vdd FILL
XFILL_0_OAI21X1_985 gnd vdd FILL
XFILL_0_OAI21X1_996 gnd vdd FILL
XFILL_27_4_1 gnd vdd FILL
XFILL_2_BUFX4_111 gnd vdd FILL
XFILL_2_4_1 gnd vdd FILL
XFILL_6_DFFPOSX1_1008 gnd vdd FILL
XFILL_2_BUFX4_144 gnd vdd FILL
XFILL_6_DFFPOSX1_1019 gnd vdd FILL
XFILL_0_OAI21X1_1740 gnd vdd FILL
XFILL_0_OAI21X1_1751 gnd vdd FILL
XFILL_0_OAI21X1_1762 gnd vdd FILL
XFILL_0_OAI21X1_1795 gnd vdd FILL
XFILL_0_OAI21X1_1784 gnd vdd FILL
XFILL_0_OAI21X1_1773 gnd vdd FILL
XFILL_10_3_1 gnd vdd FILL
XFILL_0_BUFX2_706 gnd vdd FILL
XFILL_0_NOR2X1_24 gnd vdd FILL
XFILL_0_NOR2X1_13 gnd vdd FILL
XFILL_0_BUFX2_728 gnd vdd FILL
XFILL_0_NOR2X1_57 gnd vdd FILL
XFILL_0_NOR2X1_46 gnd vdd FILL
XAOI21X1_61 bundleAddress_i[20] INVX2_110/A bundleAddress_i[19] gnd AOI21X1_61/Y vdd
+ AOI21X1
XFILL_0_BUFX2_717 gnd vdd FILL
XFILL_0_NOR2X1_35 gnd vdd FILL
XFILL_0_BUFX2_739 gnd vdd FILL
XAOI21X1_50 INVX2_101/Y AND2X2_31/Y bundleAddress_i[22] gnd AOI21X1_50/Y vdd AOI21X1
XFILL_0_NOR2X1_79 gnd vdd FILL
XFILL_0_NOR2X1_68 gnd vdd FILL
XOAI21X1_1 OAI21X1_1/A INVX2_1/Y OAI21X1_1/C gnd OAI21X1_1/Y vdd OAI21X1
XFILL_6_DFFPOSX1_117 gnd vdd FILL
XFILL_6_DFFPOSX1_139 gnd vdd FILL
XFILL_6_DFFPOSX1_128 gnd vdd FILL
XFILL_9_0_0 gnd vdd FILL
XBUFX4_303 BUFX4_303/A gnd BUFX4_303/Y vdd BUFX4
XBUFX4_336 BUFX4_380/A gnd BUFX4_336/Y vdd BUFX4
XFILL_2_OAI21X1_1823 gnd vdd FILL
XBUFX4_325 BUFX4_386/A gnd BUFX4_325/Y vdd BUFX4
XBUFX4_314 BUFX4_378/A gnd BUFX4_314/Y vdd BUFX4
XFILL_0_INVX2_202 gnd vdd FILL
XBUFX4_347 BUFX4_376/A gnd BUFX4_347/Y vdd BUFX4
XFILL_18_4_1 gnd vdd FILL
XFILL_4_DFFPOSX1_590 gnd vdd FILL
XBUFX4_358 BUFX4_388/A gnd BUFX4_358/Y vdd BUFX4
XBUFX4_369 BUFX4_384/A gnd OAI21X1_4/A vdd BUFX4
XFILL_25_18_1 gnd vdd FILL
XOAI21X1_1204 NOR3X1_15/C INVX4_49/Y INVX2_92/Y gnd NAND2X1_588/B vdd OAI21X1
XOAI21X1_1215 BUFX4_126/Y bundleAddress_i[60] OAI21X1_1215/C gnd OAI21X1_1215/Y vdd
+ OAI21X1
XOAI21X1_1237 XNOR2X1_76/Y BUFX4_146/Y OAI21X1_1237/C gnd OAI21X1_1237/Y vdd OAI21X1
XOAI21X1_1226 BUFX4_8/A BUFX4_382/Y BUFX2_190/A gnd OAI21X1_1227/C vdd OAI21X1
XFILL_1_OAI21X1_1413 gnd vdd FILL
XFILL_1_OAI21X1_1402 gnd vdd FILL
XFILL_1_OAI21X1_1424 gnd vdd FILL
XDFFPOSX1_805 BUFX2_59/A CLKBUF1_20/Y OAI21X1_1097/Y gnd vdd DFFPOSX1
XFILL_1_BUFX2_491 gnd vdd FILL
XFILL_3_DFFPOSX1_191 gnd vdd FILL
XDFFPOSX1_816 BUFX2_127/A CLKBUF1_74/Y OAI21X1_1116/Y gnd vdd DFFPOSX1
XFILL_3_DFFPOSX1_180 gnd vdd FILL
XOAI21X1_1259 BUFX4_10/Y BUFX4_356/Y BUFX2_139/A gnd OAI21X1_1261/C vdd OAI21X1
XDFFPOSX1_838 BUFX2_89/A CLKBUF1_27/Y OAI21X1_1150/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1435 gnd vdd FILL
XOAI21X1_1248 BUFX4_108/Y BUFX4_328/Y BUFX2_135/A gnd OAI21X1_1249/C vdd OAI21X1
XFILL_1_OAI21X1_1457 gnd vdd FILL
XFILL_1_CLKBUF1_60 gnd vdd FILL
XFILL_1_OAI21X1_1446 gnd vdd FILL
XFILL_1_CLKBUF1_82 gnd vdd FILL
XFILL_1_CLKBUF1_71 gnd vdd FILL
XDFFPOSX1_827 BUFX2_76/A CLKBUF1_52/Y OAI21X1_1134/Y gnd vdd DFFPOSX1
XFILL_1_CLKBUF1_93 gnd vdd FILL
XFILL_1_OAI21X1_1479 gnd vdd FILL
XFILL_1_OAI21X1_1468 gnd vdd FILL
XFILL_0_OAI21X1_215 gnd vdd FILL
XFILL_0_OAI21X1_237 gnd vdd FILL
XFILL_0_OAI21X1_226 gnd vdd FILL
XFILL_0_OAI21X1_204 gnd vdd FILL
XDFFPOSX1_849 BUFX2_101/A CLKBUF1_62/Y OAI21X1_1167/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_408 gnd vdd FILL
XFILL_0_OAI21X1_248 gnd vdd FILL
XFILL_0_OAI21X1_259 gnd vdd FILL
XFILL_1_OAI21X1_419 gnd vdd FILL
XFILL_6_DFFPOSX1_640 gnd vdd FILL
XFILL_0_NAND2X1_210 gnd vdd FILL
XFILL_1_NAND2X1_414 gnd vdd FILL
XFILL_0_NAND2X1_243 gnd vdd FILL
XFILL_1_NAND2X1_403 gnd vdd FILL
XFILL_0_NAND2X1_232 gnd vdd FILL
XFILL_0_NAND2X1_221 gnd vdd FILL
XFILL_0_OAI21X1_1014 gnd vdd FILL
XFILL_0_OAI21X1_1003 gnd vdd FILL
XFILL_0_OAI21X1_1036 gnd vdd FILL
XFILL_0_NAND2X1_265 gnd vdd FILL
XFILL_0_OAI21X1_1047 gnd vdd FILL
XFILL_1_NAND2X1_447 gnd vdd FILL
XFILL_0_DFFPOSX1_615 gnd vdd FILL
XFILL_0_DFFPOSX1_604 gnd vdd FILL
XFILL_0_NAND2X1_254 gnd vdd FILL
XFILL_0_NAND2X1_276 gnd vdd FILL
XFILL_1_NAND2X1_425 gnd vdd FILL
XFILL_0_OAI21X1_1025 gnd vdd FILL
XFILL_1_NAND2X1_469 gnd vdd FILL
XFILL_0_OAI21X1_1069 gnd vdd FILL
XFILL_0_NAND2X1_287 gnd vdd FILL
XFILL_0_NAND2X1_298 gnd vdd FILL
XFILL_0_DFFPOSX1_648 gnd vdd FILL
XFILL_0_DFFPOSX1_626 gnd vdd FILL
XFILL_0_DFFPOSX1_637 gnd vdd FILL
XFILL_0_OAI21X1_1058 gnd vdd FILL
XFILL_0_DFFPOSX1_659 gnd vdd FILL
XFILL_5_DFFPOSX1_252 gnd vdd FILL
XFILL_5_DFFPOSX1_263 gnd vdd FILL
XFILL_5_DFFPOSX1_230 gnd vdd FILL
XFILL_5_DFFPOSX1_241 gnd vdd FILL
XFILL_5_DFFPOSX1_296 gnd vdd FILL
XFILL_5_DFFPOSX1_285 gnd vdd FILL
XFILL_24_13_0 gnd vdd FILL
XFILL_5_DFFPOSX1_274 gnd vdd FILL
XOAI21X1_1760 BUFX4_147/Y BUFX4_54/Y BUFX2_763/A gnd OAI21X1_1761/C vdd OAI21X1
XOAI21X1_1793 BUFX4_353/Y INVX2_165/Y NAND2X1_734/Y gnd OAI21X1_1793/Y vdd OAI21X1
XOAI21X1_1782 BUFX4_315/Y INVX2_154/Y NAND2X1_723/Y gnd OAI21X1_1782/Y vdd OAI21X1
XOAI21X1_1771 INVX2_115/Y BUFX4_299/Y OAI21X1_1771/C gnd DFFPOSX1_98/D vdd OAI21X1
XFILL_1_OAI21X1_931 gnd vdd FILL
XFILL_2_BUFX4_27 gnd vdd FILL
XFILL_1_OAI21X1_920 gnd vdd FILL
XFILL_0_OAI21X1_782 gnd vdd FILL
XFILL_0_OAI21X1_771 gnd vdd FILL
XFILL_0_OAI21X1_760 gnd vdd FILL
XFILL_0_OAI21X1_793 gnd vdd FILL
XFILL_1_OR2X2_5 gnd vdd FILL
XFILL_1_OAI21X1_953 gnd vdd FILL
XFILL_1_OAI21X1_964 gnd vdd FILL
XFILL_1_OAI21X1_942 gnd vdd FILL
XFILL_1_OAI21X1_975 gnd vdd FILL
XFILL_1_OAI21X1_986 gnd vdd FILL
XFILL_1_OAI21X1_997 gnd vdd FILL
XFILL_2_OAI21X1_1108 gnd vdd FILL
XFILL_5_18_1 gnd vdd FILL
XBUFX2_807 BUFX2_807/A gnd tid1_o[27] vdd BUFX2
XBUFX2_818 BUFX2_818/A gnd tid1_o[17] vdd BUFX2
XFILL_2_DFFPOSX1_709 gnd vdd FILL
XBUFX2_829 BUFX2_829/A gnd tid1_o[7] vdd BUFX2
XFILL_2_NAND3X1_54 gnd vdd FILL
XFILL_29_12_0 gnd vdd FILL
XFILL_0_OAI21X1_1570 gnd vdd FILL
XFILL_0_OAI21X1_1581 gnd vdd FILL
XFILL_0_OAI21X1_1592 gnd vdd FILL
XFILL_0_BUFX2_503 gnd vdd FILL
XFILL_0_BUFX2_514 gnd vdd FILL
XFILL_0_BUFX2_547 gnd vdd FILL
XFILL_0_BUFX2_536 gnd vdd FILL
XFILL_0_BUFX2_525 gnd vdd FILL
XFILL_0_BUFX2_558 gnd vdd FILL
XFILL_0_BUFX2_569 gnd vdd FILL
XCLKBUF1_6 BUFX4_84/Y gnd CLKBUF1_6/Y vdd CLKBUF1
XBUFX4_100 BUFX4_2/A gnd BUFX4_100/Y vdd BUFX4
XBUFX4_111 BUFX4_1/A gnd BUFX4_111/Y vdd BUFX4
XFILL_0_INVX1_22 gnd vdd FILL
XBUFX4_155 BUFX4_17/Y gnd BUFX4_155/Y vdd BUFX4
XBUFX4_133 BUFX4_19/Y gnd BUFX4_133/Y vdd BUFX4
XBUFX4_122 BUFX4_13/Y gnd BUFX4_122/Y vdd BUFX4
XFILL_0_INVX1_11 gnd vdd FILL
XFILL_0_INVX1_33 gnd vdd FILL
XBUFX4_144 BUFX4_16/Y gnd BUFX4_144/Y vdd BUFX4
XFILL_4_13_0 gnd vdd FILL
XFILL_4_CLKBUF1_15 gnd vdd FILL
XFILL_2_OAI21X1_1653 gnd vdd FILL
XNOR2X1_215 INVX1_185/A NOR2X1_215/B gnd INVX4_50/A vdd NOR2X1
XFILL_4_CLKBUF1_59 gnd vdd FILL
XFILL_4_CLKBUF1_26 gnd vdd FILL
XNOR2X1_204 NOR2X1_204/A NOR2X1_204/B gnd INVX1_211/A vdd NOR2X1
XFILL_0_INVX1_44 gnd vdd FILL
XBUFX4_166 BUFX4_15/Y gnd OR2X2_20/B vdd BUFX4
XBUFX4_177 BUFX4_17/Y gnd BUFX4_177/Y vdd BUFX4
XBUFX4_188 BUFX4_21/Y gnd BUFX4_188/Y vdd BUFX4
XFILL_0_INVX1_77 gnd vdd FILL
XFILL_0_INVX1_55 gnd vdd FILL
XFILL_0_INVX1_66 gnd vdd FILL
XFILL_4_CLKBUF1_48 gnd vdd FILL
XFILL_4_CLKBUF1_37 gnd vdd FILL
XFILL_1_AND2X2_3 gnd vdd FILL
XFILL_0_INVX1_99 gnd vdd FILL
XFILL_2_OAI21X1_1686 gnd vdd FILL
XNOR2X1_226 INVX2_111/Y NOR2X1_226/B gnd NOR2X1_226/Y vdd NOR2X1
XFILL_0_INVX1_88 gnd vdd FILL
XBUFX4_199 BUFX4_20/Y gnd BUFX4_199/Y vdd BUFX4
XFILL_33_2_1 gnd vdd FILL
XFILL_24_3 gnd vdd FILL
XFILL_0_BUFX2_19 gnd vdd FILL
XFILL_17_2 gnd vdd FILL
XOAI21X1_1001 BUFX4_303/Y INVX1_155/Y OAI21X1_1001/C gnd OAI21X1_1001/Y vdd OAI21X1
XOAI21X1_1012 BUFX4_158/Y BUFX4_35/Y BUFX2_370/A gnd OAI21X1_1013/C vdd OAI21X1
XFILL_1_OAI21X1_1232 gnd vdd FILL
XOAI21X1_1045 BUFX4_382/Y INVX2_62/Y NAND2X1_411/Y gnd OAI21X1_1045/Y vdd OAI21X1
XFILL_1_OAI21X1_1221 gnd vdd FILL
XOAI21X1_1023 BUFX4_296/Y INVX1_166/Y OAI21X1_1023/C gnd OAI21X1_1023/Y vdd OAI21X1
XDFFPOSX1_613 BUFX2_258/A CLKBUF1_67/Y BUFX4_243/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1210 gnd vdd FILL
XDFFPOSX1_602 BUFX2_635/A CLKBUF1_79/Y OAI21X1_818/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_800 gnd vdd FILL
XOAI21X1_1034 BUFX4_154/Y BUFX4_51/Y BUFX2_382/A gnd OAI21X1_1035/C vdd OAI21X1
XFILL_1_DFFPOSX1_822 gnd vdd FILL
XFILL_1_OAI21X1_1254 gnd vdd FILL
XFILL_1_OAI21X1_1243 gnd vdd FILL
XDFFPOSX1_624 INVX1_53/A CLKBUF1_61/Y OAI21X1_852/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_811 gnd vdd FILL
XOAI21X1_1067 BUFX4_341/Y INVX4_39/Y NAND2X1_433/Y gnd OAI21X1_1067/Y vdd OAI21X1
XFILL_1_DFFPOSX1_833 gnd vdd FILL
XOAI21X1_1078 BUFX4_342/Y INVX2_80/Y NAND2X1_444/Y gnd OAI21X1_1078/Y vdd OAI21X1
XFILL_1_OAI21X1_1265 gnd vdd FILL
XOAI21X1_1089 NAND2X1_7/B INVX2_86/Y NAND2X1_455/Y gnd OAI21X1_1089/Y vdd OAI21X1
XDFFPOSX1_635 INVX1_64/A CLKBUF1_82/Y OAI21X1_863/Y gnd vdd DFFPOSX1
XDFFPOSX1_657 BUFX2_324/A CLKBUF1_54/Y OAI21X1_885/Y gnd vdd DFFPOSX1
XDFFPOSX1_646 INVX1_75/A CLKBUF1_54/Y OAI21X1_874/Y gnd vdd DFFPOSX1
XOAI21X1_1056 BUFX4_354/Y INVX1_173/Y NAND2X1_422/Y gnd OAI21X1_1056/Y vdd OAI21X1
XDFFPOSX1_679 BUFX2_318/A CLKBUF1_96/Y OAI21X1_907/Y gnd vdd DFFPOSX1
XDFFPOSX1_668 BUFX2_306/A CLKBUF1_96/Y OAI21X1_896/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_855 gnd vdd FILL
XFILL_1_OAI21X1_1287 gnd vdd FILL
XFILL_1_OAI21X1_1298 gnd vdd FILL
XFILL_1_DFFPOSX1_866 gnd vdd FILL
XFILL_1_OAI21X1_1276 gnd vdd FILL
XFILL_1_OAI21X1_216 gnd vdd FILL
XFILL_1_DFFPOSX1_844 gnd vdd FILL
XFILL_1_OAI21X1_205 gnd vdd FILL
XNAND2X1_705 BUFX2_697/A BUFX4_205/Y gnd NAND2X1_705/Y vdd NAND2X1
XFILL_1_OAI21X1_249 gnd vdd FILL
XNAND2X1_727 BUFX2_781/A BUFX4_322/Y gnd NAND2X1_727/Y vdd NAND2X1
XFILL_1_DFFPOSX1_888 gnd vdd FILL
XFILL_1_DFFPOSX1_877 gnd vdd FILL
XFILL_1_OAI21X1_238 gnd vdd FILL
XFILL_1_DFFPOSX1_899 gnd vdd FILL
XNAND2X1_716 BUFX2_778/A BUFX4_343/Y gnd NAND2X1_716/Y vdd NAND2X1
XFILL_1_OAI21X1_227 gnd vdd FILL
XFILL_9_12_0 gnd vdd FILL
XNAND2X1_749 BUFX2_805/A BUFX4_316/Y gnd NAND2X1_749/Y vdd NAND2X1
XNAND2X1_738 BUFX2_793/A BUFX4_375/Y gnd NAND2X1_738/Y vdd NAND2X1
XFILL_6_DFFPOSX1_481 gnd vdd FILL
XFILL_6_DFFPOSX1_492 gnd vdd FILL
XFILL_13_10_1 gnd vdd FILL
XFILL_1_NAND2X1_200 gnd vdd FILL
XFILL_1_NAND2X1_211 gnd vdd FILL
XFILL_1_NAND2X1_222 gnd vdd FILL
XFILL_24_2_1 gnd vdd FILL
XFILL_0_DFFPOSX1_412 gnd vdd FILL
XFILL_1_NAND2X1_255 gnd vdd FILL
XFILL_1_NAND2X1_233 gnd vdd FILL
XFILL_1_NAND2X1_266 gnd vdd FILL
XFILL_0_DFFPOSX1_423 gnd vdd FILL
XFILL_0_DFFPOSX1_401 gnd vdd FILL
XFILL_0_DFFPOSX1_456 gnd vdd FILL
XFILL_0_DFFPOSX1_445 gnd vdd FILL
XFILL_1_NAND2X1_288 gnd vdd FILL
XFILL_0_DFFPOSX1_434 gnd vdd FILL
XFILL_2_DFFPOSX1_9 gnd vdd FILL
XFILL_1_NAND2X1_277 gnd vdd FILL
XFILL_0_DFFPOSX1_478 gnd vdd FILL
XFILL_0_DFFPOSX1_489 gnd vdd FILL
XFILL_0_DFFPOSX1_467 gnd vdd FILL
XFILL_3_DFFPOSX1_905 gnd vdd FILL
XFILL_3_DFFPOSX1_938 gnd vdd FILL
XFILL_3_DFFPOSX1_916 gnd vdd FILL
XFILL_3_DFFPOSX1_927 gnd vdd FILL
XFILL_3_DFFPOSX1_949 gnd vdd FILL
XDFFPOSX1_50 BUFX2_719/A CLKBUF1_25/Y DFFPOSX1_50/D gnd vdd DFFPOSX1
XDFFPOSX1_61 BUFX2_731/A CLKBUF1_47/Y DFFPOSX1_61/D gnd vdd DFFPOSX1
XDFFPOSX1_72 BUFX2_771/A CLKBUF1_87/Y DFFPOSX1_72/D gnd vdd DFFPOSX1
XOAI21X1_1590 BUFX4_380/Y INVX2_126/Y NAND2X1_659/Y gnd OAI21X1_1590/Y vdd OAI21X1
XDFFPOSX1_94 BUFX2_764/A CLKBUF1_99/Y DFFPOSX1_94/D gnd vdd DFFPOSX1
XDFFPOSX1_83 BUFX2_752/A CLKBUF1_86/Y DFFPOSX1_83/D gnd vdd DFFPOSX1
XBUFX4_17 INVX8_6/Y gnd BUFX4_17/Y vdd BUFX4
XFILL_1_OAI21X1_772 gnd vdd FILL
XFILL_1_OAI21X1_761 gnd vdd FILL
XFILL_1_OAI21X1_750 gnd vdd FILL
XFILL_7_3_1 gnd vdd FILL
XFILL_0_OAI21X1_590 gnd vdd FILL
XFILL_1_INVX1_211 gnd vdd FILL
XFILL_1_OAI21X1_794 gnd vdd FILL
XFILL_15_18_0 gnd vdd FILL
XFILL_1_OAI21X1_783 gnd vdd FILL
XBUFX4_39 BUFX4_66/A gnd BUFX4_39/Y vdd BUFX4
XFILL_2_OAI21X1_954 gnd vdd FILL
XBUFX4_28 BUFX4_73/A gnd BUFX4_28/Y vdd BUFX4
XFILL_31_11_1 gnd vdd FILL
XBUFX2_637 BUFX2_637/A gnd majID4_o[7] vdd BUFX2
XBUFX2_615 BUFX2_615/A gnd majID4_o[27] vdd BUFX2
XFILL_2_DFFPOSX1_528 gnd vdd FILL
XBUFX2_604 BUFX2_604/A gnd majID4_o[37] vdd BUFX2
XFILL_2_DFFPOSX1_506 gnd vdd FILL
XFILL_2_DFFPOSX1_517 gnd vdd FILL
XBUFX2_626 BUFX2_626/A gnd majID4_o[17] vdd BUFX2
XBUFX2_659 BUFX2_659/A gnd pid1_o[13] vdd BUFX2
XFILL_2_DFFPOSX1_539 gnd vdd FILL
XFILL_0_CLKBUF1_90 gnd vdd FILL
XBUFX2_648 BUFX2_648/A gnd majID4_o[54] vdd BUFX2
XFILL_15_2_1 gnd vdd FILL
XFILL_0_DFFPOSX1_990 gnd vdd FILL
XFILL_0_BUFX2_322 gnd vdd FILL
XINVX2_111 INVX2_111/A gnd INVX2_111/Y vdd INVX2
XINVX2_100 INVX2_100/A gnd INVX2_100/Y vdd INVX2
XFILL_0_BUFX2_300 gnd vdd FILL
XFILL_0_BUFX2_311 gnd vdd FILL
XINVX2_122 bundlePid_i[26] gnd INVX2_122/Y vdd INVX2
XINVX2_133 bundlePid_i[15] gnd INVX2_133/Y vdd INVX2
XINVX2_155 bundleTid_i[54] gnd INVX2_155/Y vdd INVX2
XFILL_0_BUFX2_355 gnd vdd FILL
XFILL_1_DFFPOSX1_118 gnd vdd FILL
XFILL_0_BUFX2_366 gnd vdd FILL
XFILL_1_DFFPOSX1_107 gnd vdd FILL
XFILL_0_BUFX2_333 gnd vdd FILL
XFILL_0_BUFX2_344 gnd vdd FILL
XFILL_1_DFFPOSX1_129 gnd vdd FILL
XINVX2_144 bundlePid_i[4] gnd INVX2_144/Y vdd INVX2
XINVX2_166 bundleTid_i[43] gnd INVX2_166/Y vdd INVX2
XINVX2_199 bundleTid_i[10] gnd INVX2_199/Y vdd INVX2
XFILL_0_BUFX2_388 gnd vdd FILL
XINVX2_177 bundleTid_i[32] gnd INVX2_177/Y vdd INVX2
XFILL_0_BUFX2_399 gnd vdd FILL
XINVX2_188 bundleTid_i[21] gnd INVX2_188/Y vdd INVX2
XFILL_0_BUFX2_377 gnd vdd FILL
XFILL_36_10_1 gnd vdd FILL
XFILL_2_OAI21X1_1494 gnd vdd FILL
XOAI21X1_507 BUFX4_2/Y BUFX4_320/Y BUFX2_544/A gnd OAI21X1_508/C vdd OAI21X1
XOAI21X1_529 BUFX4_7/A BUFX4_388/Y BUFX2_523/A gnd OAI21X1_530/C vdd OAI21X1
XOAI21X1_518 INVX4_29/Y INVX4_2/Y INVX2_13/Y gnd OAI21X1_519/C vdd OAI21X1
XFILL_1_OAI21X1_1040 gnd vdd FILL
XFILL_1_NAND3X1_40 gnd vdd FILL
XFILL_1_NAND3X1_62 gnd vdd FILL
XFILL_1_NAND3X1_51 gnd vdd FILL
XDFFPOSX1_421 INVX1_6/A CLKBUF1_94/Y OAI21X1_393/Y gnd vdd DFFPOSX1
XDFFPOSX1_410 BUFX2_443/A CLKBUF1_79/Y OAI21X1_382/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1051 gnd vdd FILL
XFILL_1_DFFPOSX1_630 gnd vdd FILL
XFILL_1_OAI21X1_1062 gnd vdd FILL
XFILL_1_OAI21X1_1073 gnd vdd FILL
XFILL_1_DFFPOSX1_641 gnd vdd FILL
XDFFPOSX1_443 BUFX2_473/A CLKBUF1_18/Y OAI21X1_434/Y gnd vdd DFFPOSX1
XDFFPOSX1_432 BUFX2_461/A CLKBUF1_13/Y OAI21X1_419/Y gnd vdd DFFPOSX1
XDFFPOSX1_465 BUFX2_497/A CLKBUF1_75/Y OAI21X1_467/Y gnd vdd DFFPOSX1
XDFFPOSX1_454 BUFX2_485/A CLKBUF1_44/Y OAI21X1_452/Y gnd vdd DFFPOSX1
XFILL_38_18_0 gnd vdd FILL
XFILL_1_OAI21X1_1084 gnd vdd FILL
XFILL_1_OAI21X1_1095 gnd vdd FILL
XDFFPOSX1_476 BUFX2_509/A CLKBUF1_9/Y OAI21X1_487/Y gnd vdd DFFPOSX1
XDFFPOSX1_498 BUFX2_527/A CLKBUF1_80/Y OAI21X1_541/Y gnd vdd DFFPOSX1
XNAND2X1_502 bundleAddress_i[45] INVX1_188/A gnd INVX1_187/A vdd NAND2X1
XFILL_1_DFFPOSX1_652 gnd vdd FILL
XDFFPOSX1_487 BUFX2_544/A CLKBUF1_94/Y OAI21X1_508/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_663 gnd vdd FILL
XFILL_1_DFFPOSX1_674 gnd vdd FILL
XNAND2X1_524 BUFX2_86/A BUFX4_209/Y gnd NAND2X1_524/Y vdd NAND2X1
XNAND2X1_513 NOR2X1_140/Y INVX1_188/A gnd NOR2X1_141/B vdd NAND2X1
XFILL_1_DFFPOSX1_696 gnd vdd FILL
XNAND2X1_535 BUFX2_94/A BUFX4_226/Y gnd NAND2X1_535/Y vdd NAND2X1
XFILL_1_DFFPOSX1_685 gnd vdd FILL
XNAND2X1_557 BUFX4_243/Y INVX2_102/A gnd NAND2X1_557/Y vdd NAND2X1
XNAND2X1_568 NAND2X1_568/A NOR3X1_13/C gnd NAND2X1_568/Y vdd NAND2X1
XNAND2X1_546 bundleAddress_i[24] bundleAddress_i[23] gnd NOR3X1_16/B vdd NAND2X1
XNAND2X1_579 BUFX2_118/A BUFX4_201/Y gnd NAND2X1_579/Y vdd NAND2X1
XFILL_0_AND2X2_25 gnd vdd FILL
XFILL_0_AND2X2_14 gnd vdd FILL
XFILL_0_DFFPOSX1_220 gnd vdd FILL
XFILL_0_DFFPOSX1_231 gnd vdd FILL
XFILL_0_DFFPOSX1_242 gnd vdd FILL
XFILL_0_DFFPOSX1_275 gnd vdd FILL
XFILL_0_DFFPOSX1_253 gnd vdd FILL
XFILL_0_DFFPOSX1_264 gnd vdd FILL
XFILL_0_DFFPOSX1_297 gnd vdd FILL
XFILL_0_DFFPOSX1_286 gnd vdd FILL
XFILL_3_DFFPOSX1_713 gnd vdd FILL
XFILL_3_DFFPOSX1_702 gnd vdd FILL
XFILL_3_DFFPOSX1_746 gnd vdd FILL
XFILL_3_CLKBUF1_12 gnd vdd FILL
XFILL_3_CLKBUF1_23 gnd vdd FILL
XFILL_3_DFFPOSX1_735 gnd vdd FILL
XFILL_3_DFFPOSX1_724 gnd vdd FILL
XFILL_3_DFFPOSX1_757 gnd vdd FILL
XFILL_3_CLKBUF1_67 gnd vdd FILL
XFILL_3_CLKBUF1_45 gnd vdd FILL
XFILL_3_CLKBUF1_34 gnd vdd FILL
XFILL_3_DFFPOSX1_779 gnd vdd FILL
XFILL_3_CLKBUF1_56 gnd vdd FILL
XFILL_3_DFFPOSX1_768 gnd vdd FILL
XFILL_3_CLKBUF1_89 gnd vdd FILL
XFILL_3_CLKBUF1_78 gnd vdd FILL
XFILL_1_NOR2X1_130 gnd vdd FILL
XFILL_1_NOR2X1_141 gnd vdd FILL
XFILL_1_NOR2X1_152 gnd vdd FILL
XFILL_1_NOR2X1_174 gnd vdd FILL
XFILL_1_OAI21X1_580 gnd vdd FILL
XFILL_2_NAND3X1_5 gnd vdd FILL
XFILL_1_OAI21X1_591 gnd vdd FILL
XFILL_2_DFFPOSX1_303 gnd vdd FILL
XBUFX2_401 BUFX2_401/A gnd majID1_o[47] vdd BUFX2
XBUFX2_412 BUFX2_412/A gnd majID1_o[37] vdd BUFX2
XFILL_2_DFFPOSX1_336 gnd vdd FILL
XFILL_2_DFFPOSX1_325 gnd vdd FILL
XBUFX2_423 BUFX2_423/A gnd majID1_o[27] vdd BUFX2
XFILL_2_DFFPOSX1_314 gnd vdd FILL
XBUFX2_445 BUFX2_445/A gnd majID1_o[7] vdd BUFX2
XFILL_2_DFFPOSX1_347 gnd vdd FILL
XBUFX2_434 BUFX2_434/A gnd majID1_o[17] vdd BUFX2
XFILL_2_DFFPOSX1_358 gnd vdd FILL
XBUFX2_478 BUFX2_478/A gnd majID2_o[35] vdd BUFX2
XBUFX2_456 BUFX2_456/A gnd majID1_o[54] vdd BUFX2
XBUFX2_467 BUFX2_467/A gnd majID2_o[45] vdd BUFX2
XFILL_2_DFFPOSX1_369 gnd vdd FILL
XBUFX2_489 BUFX2_489/A gnd majID2_o[25] vdd BUFX2
XFILL_5_DFFPOSX1_818 gnd vdd FILL
XFILL_5_DFFPOSX1_807 gnd vdd FILL
XFILL_1_BUFX4_361 gnd vdd FILL
XFILL_30_0_1 gnd vdd FILL
XFILL_1_BUFX4_372 gnd vdd FILL
XFILL_1_BUFX4_383 gnd vdd FILL
XFILL_5_DFFPOSX1_829 gnd vdd FILL
XFILL_1_BUFX4_350 gnd vdd FILL
XFILL_1_XNOR2X1_19 gnd vdd FILL
XFILL_2_OAI21X1_41 gnd vdd FILL
XFILL_22_16_1 gnd vdd FILL
XFILL_0_BUFX2_130 gnd vdd FILL
XFILL_0_BUFX2_141 gnd vdd FILL
XFILL_0_BUFX2_163 gnd vdd FILL
XFILL_0_BUFX2_152 gnd vdd FILL
XFILL_0_BUFX2_174 gnd vdd FILL
XFILL_0_BUFX2_196 gnd vdd FILL
XFILL_0_BUFX2_185 gnd vdd FILL
XFILL_1_DFFPOSX1_6 gnd vdd FILL
XFILL_4_DFFPOSX1_408 gnd vdd FILL
XFILL_4_DFFPOSX1_419 gnd vdd FILL
XFILL_38_1_1 gnd vdd FILL
XFILL_2_DFFPOSX1_881 gnd vdd FILL
XFILL_2_DFFPOSX1_870 gnd vdd FILL
XFILL_2_DFFPOSX1_892 gnd vdd FILL
XBUFX2_990 BUFX2_990/A gnd tid4_o[35] vdd BUFX2
XFILL_1_BUFX2_309 gnd vdd FILL
XFILL_27_15_1 gnd vdd FILL
XFILL_21_0_1 gnd vdd FILL
XOAI21X1_304 BUFX4_130/Y BUFX4_54/Y BUFX2_1017/A gnd OAI21X1_305/C vdd OAI21X1
XOAI21X1_315 INVX2_1/Y BUFX4_295/Y OAI21X1_315/C gnd OAI21X1_315/Y vdd OAI21X1
XOAI21X1_337 BUFX4_387/Y INVX4_3/Y NAND2X1_81/Y gnd OAI21X1_337/Y vdd OAI21X1
XOAI21X1_326 BUFX4_139/Y BUFX4_68/Y BUFX2_1029/A gnd OAI21X1_327/C vdd OAI21X1
XOAI21X1_348 BUFX4_383/Y INVX2_20/Y NAND2X1_92/Y gnd OAI21X1_348/Y vdd OAI21X1
XOAI21X1_359 BUFX4_314/Y INVX2_24/Y OAI21X1_359/C gnd OAI21X1_359/Y vdd OAI21X1
XFILL_21_11_0 gnd vdd FILL
XDFFPOSX1_240 BUFX2_909/A CLKBUF1_25/Y OAI21X1_97/Y gnd vdd DFFPOSX1
XBUFX4_2 BUFX4_2/A gnd BUFX4_2/Y vdd BUFX4
XDFFPOSX1_273 BUFX2_945/A CLKBUF1_102/Y OAI21X1_163/Y gnd vdd DFFPOSX1
XDFFPOSX1_262 BUFX2_933/A CLKBUF1_11/Y OAI21X1_141/Y gnd vdd DFFPOSX1
XDFFPOSX1_251 BUFX2_921/A CLKBUF1_86/Y OAI21X1_119/Y gnd vdd DFFPOSX1
XDFFPOSX1_284 BUFX2_957/A CLKBUF1_43/Y OAI21X1_185/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_493 gnd vdd FILL
XFILL_1_DFFPOSX1_471 gnd vdd FILL
XFILL_1_DFFPOSX1_482 gnd vdd FILL
XFILL_1_DFFPOSX1_460 gnd vdd FILL
XDFFPOSX1_295 BUFX2_992/A CLKBUF1_88/Y OAI21X1_207/Y gnd vdd DFFPOSX1
XNAND2X1_310 bundleStartMajId_i[55] AND2X2_18/Y gnd INVX1_35/A vdd NAND2X1
XNAND2X1_354 BUFX4_265/Y bundle_i[15] gnd OAI21X1_860/C vdd NAND2X1
XNAND2X1_343 BUFX4_265/Y bundle_i[26] gnd OAI21X1_849/C vdd NAND2X1
XFILL_3_NOR3X1_15 gnd vdd FILL
XNAND2X1_332 NAND3X1_34/Y OAI21X1_820/Y gnd OAI21X1_821/A vdd NAND2X1
XNAND2X1_321 INVX2_42/Y INVX1_38/A gnd XNOR2X1_46/A vdd NAND2X1
XFILL_4_DFFPOSX1_920 gnd vdd FILL
XNAND2X1_376 BUFX2_321/A BUFX4_205/Y gnd OAI21X1_882/C vdd NAND2X1
XFILL_4_DFFPOSX1_931 gnd vdd FILL
XNAND2X1_365 BUFX4_264/Y bundle_i[4] gnd OAI21X1_871/C vdd NAND2X1
XNAND2X1_387 BUFX2_302/A BUFX4_199/Y gnd OAI21X1_893/C vdd NAND2X1
XFILL_4_DFFPOSX1_942 gnd vdd FILL
XFILL_29_1_1 gnd vdd FILL
XFILL_4_DFFPOSX1_953 gnd vdd FILL
XFILL_4_DFFPOSX1_964 gnd vdd FILL
XNAND2X1_398 BUFX2_314/A BUFX4_189/Y gnd OAI21X1_904/C vdd NAND2X1
XFILL_4_1_1 gnd vdd FILL
XFILL_0_INVX1_119 gnd vdd FILL
XFILL_0_INVX1_108 gnd vdd FILL
XFILL_4_DFFPOSX1_997 gnd vdd FILL
XFILL_2_16_1 gnd vdd FILL
XFILL_4_DFFPOSX1_986 gnd vdd FILL
XFILL_4_DFFPOSX1_975 gnd vdd FILL
XFILL_1_AOI21X1_19 gnd vdd FILL
XFILL_1_BUFX2_821 gnd vdd FILL
XFILL_12_0_1 gnd vdd FILL
XFILL_26_10_0 gnd vdd FILL
XFILL_1_INVX2_87 gnd vdd FILL
XFILL_1_BUFX2_832 gnd vdd FILL
XFILL_1_BUFX2_843 gnd vdd FILL
XINVX4_2 bundleStartMajId_i[57] gnd INVX4_2/Y vdd INVX4
XFILL_1_BUFX2_887 gnd vdd FILL
XOAI21X1_860 INVX1_61/Y BUFX4_265/Y OAI21X1_860/C gnd OAI21X1_860/Y vdd OAI21X1
XFILL_3_DFFPOSX1_510 gnd vdd FILL
XFILL_2_NOR3X1_7 gnd vdd FILL
XFILL_3_DFFPOSX1_521 gnd vdd FILL
XFILL_1_BUFX2_876 gnd vdd FILL
XOAI21X1_882 INVX1_83/Y BUFX4_205/Y OAI21X1_882/C gnd OAI21X1_882/Y vdd OAI21X1
XFILL_3_DFFPOSX1_543 gnd vdd FILL
XFILL_1_OAI21X1_1809 gnd vdd FILL
XFILL_3_DFFPOSX1_565 gnd vdd FILL
XFILL_3_DFFPOSX1_532 gnd vdd FILL
XOAI21X1_871 INVX1_72/Y BUFX4_264/Y OAI21X1_871/C gnd OAI21X1_871/Y vdd OAI21X1
XOAI21X1_893 INVX1_94/Y BUFX4_199/Y OAI21X1_893/C gnd OAI21X1_893/Y vdd OAI21X1
XFILL_3_DFFPOSX1_554 gnd vdd FILL
XFILL_3_DFFPOSX1_598 gnd vdd FILL
XFILL_3_DFFPOSX1_587 gnd vdd FILL
XFILL_3_DFFPOSX1_576 gnd vdd FILL
XFILL_7_15_1 gnd vdd FILL
XFILL_2_DFFPOSX1_111 gnd vdd FILL
XFILL_2_DFFPOSX1_100 gnd vdd FILL
XFILL_2_DFFPOSX1_122 gnd vdd FILL
XBUFX2_220 BUFX2_220/A gnd addr4_o[30] vdd BUFX2
XFILL_0_NAND2X1_617 gnd vdd FILL
XFILL_0_NAND2X1_606 gnd vdd FILL
XFILL_2_DFFPOSX1_133 gnd vdd FILL
XFILL_2_DFFPOSX1_144 gnd vdd FILL
XFILL_0_NAND2X1_628 gnd vdd FILL
XBUFX2_253 BUFX2_253/A gnd addr4_o[0] vdd BUFX2
XFILL_2_DFFPOSX1_155 gnd vdd FILL
XFILL_0_NAND2X1_639 gnd vdd FILL
XBUFX2_231 BUFX2_231/A gnd addr4_o[20] vdd BUFX2
XFILL_1_11_0 gnd vdd FILL
XBUFX2_242 BUFX2_242/A gnd addr4_o[10] vdd BUFX2
XFILL_2_DFFPOSX1_188 gnd vdd FILL
XBUFX2_264 INVX1_56/A gnd instr1_o[20] vdd BUFX2
XFILL_2_DFFPOSX1_166 gnd vdd FILL
XBUFX2_286 INVX1_76/A gnd instr1_o[0] vdd BUFX2
XBUFX2_275 INVX1_66/A gnd instr1_o[10] vdd BUFX2
XFILL_2_DFFPOSX1_177 gnd vdd FILL
XFILL_32_8_0 gnd vdd FILL
XFILL_2_DFFPOSX1_199 gnd vdd FILL
XBUFX2_297 BUFX2_297/A gnd instr2_o[19] vdd BUFX2
XFILL_5_DFFPOSX1_615 gnd vdd FILL
XFILL_5_DFFPOSX1_604 gnd vdd FILL
XFILL_5_DFFPOSX1_626 gnd vdd FILL
XFILL_5_DFFPOSX1_637 gnd vdd FILL
XFILL_1_BUFX4_191 gnd vdd FILL
XFILL_1_BUFX4_180 gnd vdd FILL
XFILL_5_DFFPOSX1_648 gnd vdd FILL
XFILL_5_DFFPOSX1_659 gnd vdd FILL
XNAND3X1_5 NOR2X1_29/Y AND2X2_6/Y NOR2X1_28/Y gnd NOR2X1_30/B vdd NAND3X1
XFILL_4_DFFPOSX1_205 gnd vdd FILL
XFILL_4_DFFPOSX1_216 gnd vdd FILL
XFILL_4_DFFPOSX1_227 gnd vdd FILL
XFILL_4_DFFPOSX1_249 gnd vdd FILL
XFILL_4_DFFPOSX1_238 gnd vdd FILL
XFILL_6_10_0 gnd vdd FILL
XFILL_2_CLKBUF1_31 gnd vdd FILL
XFILL_2_BUFX4_304 gnd vdd FILL
XFILL_2_CLKBUF1_20 gnd vdd FILL
XFILL_2_CLKBUF1_42 gnd vdd FILL
XFILL_2_CLKBUF1_64 gnd vdd FILL
XFILL_2_BUFX4_337 gnd vdd FILL
XFILL_2_CLKBUF1_75 gnd vdd FILL
XFILL_2_CLKBUF1_53 gnd vdd FILL
XFILL_2_CLKBUF1_86 gnd vdd FILL
XFILL_2_CLKBUF1_97 gnd vdd FILL
XFILL_23_8_0 gnd vdd FILL
XFILL_1_BUFX2_106 gnd vdd FILL
XFILL_1_BUFX2_117 gnd vdd FILL
XOAI21X1_101 BUFX4_165/Y INVX2_160/Y OAI21X1_101/C gnd OAI21X1_101/Y vdd OAI21X1
XOAI21X1_112 BUFX4_10/Y BUFX4_340/Y BUFX2_918/A gnd OAI21X1_113/C vdd OAI21X1
XFILL_0_NOR2X1_182 gnd vdd FILL
XFILL_0_NOR2X1_160 gnd vdd FILL
XFILL_1_BUFX2_128 gnd vdd FILL
XFILL_0_NOR2X1_171 gnd vdd FILL
XFILL_0_DFFPOSX1_1012 gnd vdd FILL
XOAI21X1_123 BUFX4_138/Y INVX2_171/Y OAI21X1_123/C gnd OAI21X1_123/Y vdd OAI21X1
XFILL_0_DFFPOSX1_1001 gnd vdd FILL
XOAI21X1_134 BUFX4_107/Y BUFX4_366/Y BUFX2_930/A gnd OAI21X1_135/C vdd OAI21X1
XFILL_0_NOR2X1_193 gnd vdd FILL
XOAI21X1_145 BUFX4_157/Y INVX2_182/Y OAI21X1_145/C gnd OAI21X1_145/Y vdd OAI21X1
XOAI21X1_156 BUFX4_4/A BUFX4_326/Y BUFX2_942/A gnd OAI21X1_157/C vdd OAI21X1
XOAI21X1_178 BUFX4_11/A BUFX4_318/Y BUFX2_954/A gnd OAI21X1_179/C vdd OAI21X1
XOAI21X1_167 BUFX4_159/Y INVX2_193/Y OAI21X1_167/C gnd OAI21X1_167/Y vdd OAI21X1
XFILL_0_DFFPOSX1_1023 gnd vdd FILL
XOAI21X1_189 BUFX4_133/Y INVX2_2/Y OAI21X1_189/C gnd OAI21X1_189/Y vdd OAI21X1
XINVX1_209 INVX1_209/A gnd INVX1_209/Y vdd INVX1
XFILL_1_DFFPOSX1_290 gnd vdd FILL
XNAND2X1_140 BUFX2_469/A BUFX4_180/Y gnd OAI21X1_396/C vdd NAND2X1
XNAND2X1_151 NOR2X1_5/B OAI21X1_408/Y gnd OAI21X1_409/A vdd NAND2X1
XFILL_6_9_0 gnd vdd FILL
XNAND2X1_162 bundleStartMajId_i[55] bundleStartMajId_i[52] gnd NOR2X1_7/B vdd NAND2X1
XFILL_0_XNOR2X1_16 gnd vdd FILL
XNAND2X1_195 NOR2X1_19/Y NOR2X1_17/Y gnd XNOR2X1_11/A vdd NAND2X1
XFILL_0_XNOR2X1_27 gnd vdd FILL
XNAND2X1_184 BUFX2_473/A BUFX4_233/Y gnd OAI21X1_434/C vdd NAND2X1
XNAND2X1_173 BUFX2_467/A BUFX4_236/Y gnd OAI21X1_427/C vdd NAND2X1
XFILL_4_DFFPOSX1_761 gnd vdd FILL
XFILL_4_DFFPOSX1_750 gnd vdd FILL
XFILL_4_DFFPOSX1_772 gnd vdd FILL
XFILL_0_XNOR2X1_38 gnd vdd FILL
XFILL_0_XNOR2X1_49 gnd vdd FILL
XFILL_1_OAI21X1_60 gnd vdd FILL
XFILL_4_DFFPOSX1_783 gnd vdd FILL
XFILL_1_OAI21X1_93 gnd vdd FILL
XFILL_12_16_0 gnd vdd FILL
XFILL_1_OAI21X1_71 gnd vdd FILL
XFILL_1_OAI21X1_82 gnd vdd FILL
XFILL_4_DFFPOSX1_794 gnd vdd FILL
XFILL_14_8_0 gnd vdd FILL
XFILL_0_DFFPOSX1_3 gnd vdd FILL
XFILL_0_BUFX4_203 gnd vdd FILL
XFILL_1_BUFX2_640 gnd vdd FILL
XFILL_1_BUFX2_673 gnd vdd FILL
XFILL_0_BUFX4_214 gnd vdd FILL
XFILL_0_BUFX4_247 gnd vdd FILL
XFILL_3_DFFPOSX1_340 gnd vdd FILL
XFILL_1_BUFX2_695 gnd vdd FILL
XOAI21X1_1408 NOR2X1_217/Y OAI21X1_1408/B OAI21X1_1408/C gnd OAI21X1_1408/Y vdd OAI21X1
XOAI21X1_1419 BUFX4_156/Y BUFX4_62/Y BUFX2_197/A gnd OAI21X1_1420/C vdd OAI21X1
XFILL_1_BUFX2_684 gnd vdd FILL
XFILL_0_BUFX4_258 gnd vdd FILL
XFILL_0_BUFX4_225 gnd vdd FILL
XFILL_1_OAI21X1_1606 gnd vdd FILL
XFILL_0_BUFX4_236 gnd vdd FILL
XFILL_1_OAI21X1_1628 gnd vdd FILL
XFILL_0_BUFX4_269 gnd vdd FILL
XFILL_1_OAI21X1_1639 gnd vdd FILL
XNOR3X1_8 NOR3X1_8/A NOR3X1_8/B NOR3X1_8/C gnd NOR3X1_8/Y vdd NOR3X1
XFILL_3_DFFPOSX1_373 gnd vdd FILL
XFILL_1_OAI21X1_1617 gnd vdd FILL
XFILL_3_DFFPOSX1_362 gnd vdd FILL
XOAI21X1_690 NOR2X1_104/A INVX1_35/A OAI21X1_690/C gnd OAI21X1_692/A vdd OAI21X1
XFILL_3_DFFPOSX1_351 gnd vdd FILL
XFILL_3_DFFPOSX1_395 gnd vdd FILL
XFILL_0_OAI21X1_419 gnd vdd FILL
XFILL_3_DFFPOSX1_384 gnd vdd FILL
XFILL_0_OAI21X1_408 gnd vdd FILL
XFILL_6_DFFPOSX1_811 gnd vdd FILL
XFILL_0_INVX4_11 gnd vdd FILL
XFILL_6_DFFPOSX1_800 gnd vdd FILL
XFILL_3_DFFPOSX1_1005 gnd vdd FILL
XFILL_6_DFFPOSX1_822 gnd vdd FILL
XFILL_0_INVX4_33 gnd vdd FILL
XFILL_0_INVX4_22 gnd vdd FILL
XFILL_0_INVX4_44 gnd vdd FILL
XFILL_3_DFFPOSX1_1027 gnd vdd FILL
XFILL_3_DFFPOSX1_1016 gnd vdd FILL
XFILL_17_15_0 gnd vdd FILL
XXNOR2X1_40 INVX2_52/A bundleStartMajId_i[59] gnd XNOR2X1_40/Y vdd XNOR2X1
XFILL_5_2 gnd vdd FILL
XXNOR2X1_73 XNOR2X1_73/A INVX2_81/Y gnd XNOR2X1_73/Y vdd XNOR2X1
XXNOR2X1_62 XNOR2X1_62/A bundleAddress_i[39] gnd XNOR2X1_62/Y vdd XNOR2X1
XXNOR2X1_51 XNOR2X1_51/A INVX4_18/Y gnd XNOR2X1_51/Y vdd XNOR2X1
XXNOR2X1_84 NOR3X1_16/C INVX8_3/Y gnd XNOR2X1_84/Y vdd XNOR2X1
XXNOR2X1_95 XNOR2X1_95/A bundleAddress_i[40] gnd XNOR2X1_95/Y vdd XNOR2X1
XFILL_0_NAND2X1_414 gnd vdd FILL
XFILL_30_17_0 gnd vdd FILL
XFILL_0_NAND2X1_403 gnd vdd FILL
XFILL_0_NAND2X1_425 gnd vdd FILL
XFILL_1_XNOR2X1_7 gnd vdd FILL
XBUFX2_72 BUFX2_72/A gnd addr2_o[48] vdd BUFX2
XFILL_0_OAI21X1_1229 gnd vdd FILL
XFILL_0_OAI21X1_1218 gnd vdd FILL
XFILL_0_NAND2X1_469 gnd vdd FILL
XFILL_0_NAND2X1_447 gnd vdd FILL
XFILL_1_NAND2X1_607 gnd vdd FILL
XBUFX2_61 BUFX2_61/A gnd addr1_o[0] vdd BUFX2
XFILL_1_NAND2X1_618 gnd vdd FILL
XFILL_0_OAI21X1_1207 gnd vdd FILL
XFILL_0_NAND2X1_436 gnd vdd FILL
XFILL_0_NAND2X1_458 gnd vdd FILL
XBUFX2_50 BUFX2_50/A gnd addr1_o[10] vdd BUFX2
XFILL_0_DFFPOSX1_808 gnd vdd FILL
XBUFX2_83 BUFX2_83/A gnd addr2_o[38] vdd BUFX2
XFILL_0_DFFPOSX1_819 gnd vdd FILL
XBUFX2_94 BUFX2_94/A gnd addr2_o[28] vdd BUFX2
XFILL_5_DFFPOSX1_412 gnd vdd FILL
XFILL_5_DFFPOSX1_401 gnd vdd FILL
XFILL_5_DFFPOSX1_445 gnd vdd FILL
XFILL_5_DFFPOSX1_423 gnd vdd FILL
XFILL_5_DFFPOSX1_434 gnd vdd FILL
XFILL_5_DFFPOSX1_478 gnd vdd FILL
XFILL_5_DFFPOSX1_456 gnd vdd FILL
XFILL_5_DFFPOSX1_467 gnd vdd FILL
XFILL_1_BUFX4_50 gnd vdd FILL
XFILL_1_BUFX4_72 gnd vdd FILL
XFILL_1_BUFX4_61 gnd vdd FILL
XFILL_5_DFFPOSX1_489 gnd vdd FILL
XFILL_1_BUFX4_94 gnd vdd FILL
XFILL_1_BUFX4_83 gnd vdd FILL
XFILL_0_AOI21X1_38 gnd vdd FILL
XFILL_0_AOI21X1_27 gnd vdd FILL
XFILL_0_AOI21X1_16 gnd vdd FILL
XFILL_0_OAI21X1_931 gnd vdd FILL
XFILL_2_CLKBUF1_7 gnd vdd FILL
XFILL_0_AOI21X1_49 gnd vdd FILL
XFILL_0_OAI21X1_942 gnd vdd FILL
XFILL_0_OAI21X1_920 gnd vdd FILL
XFILL_0_OAI21X1_975 gnd vdd FILL
XFILL_0_OAI21X1_953 gnd vdd FILL
XFILL_0_OAI21X1_964 gnd vdd FILL
XFILL_35_16_0 gnd vdd FILL
XFILL_0_OAI21X1_986 gnd vdd FILL
XFILL_0_OAI21X1_997 gnd vdd FILL
XFILL_1_OR2X2_20 gnd vdd FILL
XFILL_0_OAI21X1_1730 gnd vdd FILL
XFILL_0_OAI21X1_1741 gnd vdd FILL
XFILL_0_OAI21X1_1752 gnd vdd FILL
XFILL_2_BUFX4_189 gnd vdd FILL
XFILL_0_OAI21X1_1785 gnd vdd FILL
XFILL_0_OAI21X1_1763 gnd vdd FILL
XFILL_0_OAI21X1_1774 gnd vdd FILL
XFILL_0_OAI21X1_1796 gnd vdd FILL
XFILL_5_DFFPOSX1_990 gnd vdd FILL
XFILL_0_NOR2X1_14 gnd vdd FILL
XFILL_0_BUFX2_729 gnd vdd FILL
XAOI21X1_40 bundleAddress_i[16] INVX2_102/Y bundleAddress_i[15] gnd AOI21X1_40/Y vdd
+ AOI21X1
XAOI21X1_62 bundleAddress_i[16] INVX1_225/Y bundleAddress_i[15] gnd AOI21X1_62/Y vdd
+ AOI21X1
XAOI21X1_51 bundleAddress_i[20] NOR3X1_17/Y bundleAddress_i[19] gnd AOI21X1_51/Y vdd
+ AOI21X1
XFILL_0_NOR2X1_47 gnd vdd FILL
XFILL_0_NOR2X1_36 gnd vdd FILL
XFILL_0_BUFX2_707 gnd vdd FILL
XFILL_0_NOR2X1_25 gnd vdd FILL
XFILL_0_BUFX2_718 gnd vdd FILL
XFILL_0_NOR2X1_69 gnd vdd FILL
XFILL_0_NOR2X1_58 gnd vdd FILL
XFILL_6_DFFPOSX1_107 gnd vdd FILL
XOAI21X1_2 OAI21X1_2/A INVX2_2/Y OAI21X1_2/C gnd OAI21X1_2/Y vdd OAI21X1
XFILL_9_0_1 gnd vdd FILL
XBUFX4_304 BUFX4_310/A gnd NOR2X1_89/B vdd BUFX4
XBUFX4_326 BUFX4_378/A gnd BUFX4_326/Y vdd BUFX4
XBUFX4_315 BUFX4_388/A gnd BUFX4_315/Y vdd BUFX4
XBUFX4_337 BUFX4_385/A gnd BUFX4_337/Y vdd BUFX4
XBUFX4_359 BUFX4_385/A gnd BUFX4_359/Y vdd BUFX4
XFILL_4_DFFPOSX1_591 gnd vdd FILL
XBUFX4_348 BUFX4_381/A gnd BUFX4_348/Y vdd BUFX4
XFILL_4_DFFPOSX1_580 gnd vdd FILL
XFILL_1_BUFX2_481 gnd vdd FILL
XFILL_1_BUFX2_470 gnd vdd FILL
XOAI21X1_1227 OAI21X1_1227/A NOR2X1_178/Y OAI21X1_1227/C gnd OAI21X1_1227/Y vdd OAI21X1
XOAI21X1_1216 BUFX4_8/Y BUFX4_368/Y BUFX2_163/A gnd OAI21X1_1217/C vdd OAI21X1
XOAI21X1_1238 INVX1_201/A INVX4_33/Y INVX2_64/Y gnd OAI21X1_1239/C vdd OAI21X1
XFILL_1_OAI21X1_1414 gnd vdd FILL
XFILL_1_OAI21X1_1403 gnd vdd FILL
XDFFPOSX1_806 BUFX2_60/A CLKBUF1_30/Y OAI21X1_1098/Y gnd vdd DFFPOSX1
XOAI21X1_1205 NAND2X1_588/Y NOR3X1_15/Y NAND2X1_587/Y gnd OAI21X1_1205/Y vdd OAI21X1
XFILL_1_INVX8_1 gnd vdd FILL
XFILL_1_BUFX2_492 gnd vdd FILL
XFILL_3_DFFPOSX1_181 gnd vdd FILL
XFILL_1_OAI21X1_1425 gnd vdd FILL
XOAI21X1_1249 OAI21X1_1249/A BUFX4_146/Y OAI21X1_1249/C gnd OAI21X1_1249/Y vdd OAI21X1
XDFFPOSX1_839 BUFX2_90/A CLKBUF1_89/Y OAI21X1_1152/Y gnd vdd DFFPOSX1
XFILL_1_CLKBUF1_61 gnd vdd FILL
XFILL_1_OAI21X1_1436 gnd vdd FILL
XFILL_1_CLKBUF1_72 gnd vdd FILL
XFILL_3_DFFPOSX1_170 gnd vdd FILL
XFILL_1_CLKBUF1_50 gnd vdd FILL
XDFFPOSX1_817 BUFX2_128/A CLKBUF1_84/Y OAI21X1_1119/Y gnd vdd DFFPOSX1
XFILL_1_CLKBUF1_83 gnd vdd FILL
XFILL_1_OAI21X1_1447 gnd vdd FILL
XDFFPOSX1_828 BUFX2_78/A CLKBUF1_34/Y OAI21X1_1136/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1458 gnd vdd FILL
XFILL_1_OAI21X1_1469 gnd vdd FILL
XFILL_1_CLKBUF1_94 gnd vdd FILL
XFILL_0_OAI21X1_216 gnd vdd FILL
XFILL_3_DFFPOSX1_192 gnd vdd FILL
XFILL_0_OAI21X1_205 gnd vdd FILL
XFILL_0_OAI21X1_227 gnd vdd FILL
XFILL_0_OAI21X1_249 gnd vdd FILL
XFILL_0_OAI21X1_238 gnd vdd FILL
XFILL_1_OAI21X1_409 gnd vdd FILL
XFILL_6_DFFPOSX1_663 gnd vdd FILL
XFILL_6_DFFPOSX1_696 gnd vdd FILL
XFILL_6_DFFPOSX1_674 gnd vdd FILL
XFILL_6_DFFPOSX1_685 gnd vdd FILL
XFILL_37_7_0 gnd vdd FILL
XFILL_0_NAND2X1_200 gnd vdd FILL
XFILL_1_NAND2X1_404 gnd vdd FILL
XFILL_1_NAND2X1_415 gnd vdd FILL
XFILL_0_NAND2X1_211 gnd vdd FILL
XFILL_0_NAND2X1_222 gnd vdd FILL
XFILL_0_NAND2X1_233 gnd vdd FILL
XFILL_0_OAI21X1_1004 gnd vdd FILL
XFILL_0_OAI21X1_1048 gnd vdd FILL
XFILL_0_DFFPOSX1_605 gnd vdd FILL
XFILL_1_NAND2X1_448 gnd vdd FILL
XFILL_0_OAI21X1_1037 gnd vdd FILL
XFILL_0_NAND2X1_255 gnd vdd FILL
XFILL_0_NAND2X1_266 gnd vdd FILL
XFILL_0_NAND2X1_244 gnd vdd FILL
XFILL_0_OAI21X1_1015 gnd vdd FILL
XFILL_0_OAI21X1_1026 gnd vdd FILL
XFILL_1_NAND2X1_426 gnd vdd FILL
XFILL_0_NAND2X1_277 gnd vdd FILL
XFILL_0_DFFPOSX1_649 gnd vdd FILL
XFILL_0_DFFPOSX1_627 gnd vdd FILL
XFILL_0_NAND2X1_299 gnd vdd FILL
XFILL_0_NAND2X1_288 gnd vdd FILL
XFILL_0_DFFPOSX1_616 gnd vdd FILL
XFILL_0_DFFPOSX1_638 gnd vdd FILL
XFILL_0_OAI21X1_1059 gnd vdd FILL
XFILL_5_DFFPOSX1_220 gnd vdd FILL
XFILL_5_DFFPOSX1_242 gnd vdd FILL
XFILL_5_DFFPOSX1_253 gnd vdd FILL
XFILL_20_6_0 gnd vdd FILL
XFILL_5_DFFPOSX1_231 gnd vdd FILL
XFILL_5_DFFPOSX1_275 gnd vdd FILL
XFILL_24_13_1 gnd vdd FILL
XFILL_5_DFFPOSX1_264 gnd vdd FILL
XFILL_5_DFFPOSX1_286 gnd vdd FILL
XFILL_5_DFFPOSX1_297 gnd vdd FILL
XFILL_0_OAI21X1_90 gnd vdd FILL
XOAI21X1_1750 BUFX4_144/Y BUFX4_73/Y BUFX2_758/A gnd OAI21X1_1751/C vdd OAI21X1
XOAI21X1_1783 BUFX4_378/Y INVX2_155/Y NAND2X1_724/Y gnd OAI21X1_1783/Y vdd OAI21X1
XOAI21X1_1761 INVX2_142/Y BUFX4_295/Y OAI21X1_1761/C gnd DFFPOSX1_93/D vdd OAI21X1
XOAI21X1_1794 BUFX4_383/Y INVX2_166/Y NAND2X1_735/Y gnd OAI21X1_1794/Y vdd OAI21X1
XOAI21X1_1772 BUFX4_163/Y BUFX4_30/Y BUFX2_770/A gnd OAI21X1_1773/C vdd OAI21X1
XFILL_1_OAI21X1_910 gnd vdd FILL
XFILL_0_OAI21X1_750 gnd vdd FILL
XFILL_1_OAI21X1_921 gnd vdd FILL
XFILL_1_OAI21X1_932 gnd vdd FILL
XFILL_0_OAI21X1_772 gnd vdd FILL
XFILL_0_OAI21X1_761 gnd vdd FILL
XFILL_0_OAI21X1_783 gnd vdd FILL
XFILL_1_OAI21X1_954 gnd vdd FILL
XFILL_1_OAI21X1_943 gnd vdd FILL
XFILL_1_OAI21X1_998 gnd vdd FILL
XFILL_1_OAI21X1_976 gnd vdd FILL
XFILL_0_OAI21X1_794 gnd vdd FILL
XFILL_1_OR2X2_6 gnd vdd FILL
XFILL_1_OAI21X1_987 gnd vdd FILL
XFILL_1_OAI21X1_965 gnd vdd FILL
XFILL_2_OAI21X1_1109 gnd vdd FILL
XBUFX2_808 BUFX2_808/A gnd tid1_o[26] vdd BUFX2
XBUFX2_819 BUFX2_819/A gnd tid1_o[16] vdd BUFX2
XFILL_28_7_0 gnd vdd FILL
XFILL_3_7_0 gnd vdd FILL
XFILL_29_12_1 gnd vdd FILL
XFILL_0_OAI21X1_1560 gnd vdd FILL
XFILL_0_OAI21X1_1582 gnd vdd FILL
XFILL_0_OAI21X1_1571 gnd vdd FILL
XFILL_0_OAI21X1_1593 gnd vdd FILL
XFILL_11_6_0 gnd vdd FILL
XFILL_0_BUFX2_504 gnd vdd FILL
XFILL_0_BUFX2_515 gnd vdd FILL
XFILL_0_BUFX2_537 gnd vdd FILL
XFILL_0_BUFX2_548 gnd vdd FILL
XFILL_0_BUFX2_526 gnd vdd FILL
XCLKBUF1_7 BUFX4_86/Y gnd CLKBUF1_7/Y vdd CLKBUF1
XFILL_0_BUFX2_559 gnd vdd FILL
XBUFX4_101 BUFX4_94/A gnd BUFX4_101/Y vdd BUFX4
XBUFX4_112 BUFX4_9/A gnd BUFX4_112/Y vdd BUFX4
XBUFX4_123 BUFX4_14/Y gnd BUFX4_123/Y vdd BUFX4
XFILL_4_CLKBUF1_16 gnd vdd FILL
XFILL_0_INVX1_23 gnd vdd FILL
XBUFX4_145 BUFX4_18/Y gnd BUFX4_145/Y vdd BUFX4
XFILL_2_OAI21X1_1632 gnd vdd FILL
XFILL_19_7_0 gnd vdd FILL
XFILL_0_INVX1_12 gnd vdd FILL
XBUFX4_134 BUFX4_13/Y gnd BUFX4_134/Y vdd BUFX4
XFILL_2_OAI21X1_1610 gnd vdd FILL
XFILL_4_13_1 gnd vdd FILL
XFILL_0_INVX1_34 gnd vdd FILL
XBUFX4_178 BUFX4_15/Y gnd BUFX4_178/Y vdd BUFX4
XNOR2X1_216 NOR2X1_216/A INVX4_50/Y gnd INVX1_219/A vdd NOR2X1
XFILL_4_CLKBUF1_27 gnd vdd FILL
XBUFX4_156 BUFX4_17/Y gnd BUFX4_156/Y vdd BUFX4
XNOR2X1_205 bundleAddress_i[16] INVX1_212/Y gnd NOR2X1_205/Y vdd NOR2X1
XFILL_0_INVX1_56 gnd vdd FILL
XBUFX4_167 BUFX4_13/Y gnd BUFX4_167/Y vdd BUFX4
XFILL_1_AND2X2_4 gnd vdd FILL
XFILL_0_INVX1_67 gnd vdd FILL
XFILL_0_INVX1_45 gnd vdd FILL
XFILL_4_CLKBUF1_38 gnd vdd FILL
XFILL_0_INVX1_78 gnd vdd FILL
XNOR2X1_227 bundleAddress_i[16] INVX1_225/Y gnd NOR2X1_227/Y vdd NOR2X1
XFILL_0_INVX1_89 gnd vdd FILL
XBUFX4_189 BUFX4_21/Y gnd BUFX4_189/Y vdd BUFX4
XFILL_24_4 gnd vdd FILL
XOAI21X1_1002 BUFX4_144/Y BUFX4_58/Y BUFX2_364/A gnd OAI21X1_1003/C vdd OAI21X1
XOAI21X1_1013 BUFX4_303/Y INVX1_161/Y OAI21X1_1013/C gnd OAI21X1_1013/Y vdd OAI21X1
XFILL_1_OAI21X1_1222 gnd vdd FILL
XOAI21X1_1046 BUFX4_328/Y INVX2_63/Y NAND2X1_412/Y gnd OAI21X1_1046/Y vdd OAI21X1
XFILL_1_OAI21X1_1211 gnd vdd FILL
XFILL_1_OAI21X1_1200 gnd vdd FILL
XDFFPOSX1_603 BUFX2_636/A CLKBUF1_60/Y OAI21X1_821/Y gnd vdd DFFPOSX1
XOAI21X1_1024 BUFX4_154/Y BUFX4_73/Y BUFX2_376/A gnd OAI21X1_1025/C vdd OAI21X1
XDFFPOSX1_614 BUFX2_259/A CLKBUF1_76/Y BUFX4_308/Y gnd vdd DFFPOSX1
XOAI21X1_1035 BUFX4_303/Y INVX1_172/Y OAI21X1_1035/C gnd OAI21X1_1035/Y vdd OAI21X1
XFILL_1_DFFPOSX1_812 gnd vdd FILL
XFILL_1_OAI21X1_1233 gnd vdd FILL
XDFFPOSX1_636 INVX1_65/A CLKBUF1_96/Y OAI21X1_864/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1255 gnd vdd FILL
XOAI21X1_1068 BUFX4_381/Y INVX2_74/Y NAND2X1_434/Y gnd OAI21X1_1068/Y vdd OAI21X1
XFILL_1_DFFPOSX1_823 gnd vdd FILL
XFILL_1_OAI21X1_1244 gnd vdd FILL
XOAI21X1_1079 BUFX4_344/Y INVX4_43/Y NAND2X1_445/Y gnd OAI21X1_1079/Y vdd OAI21X1
XFILL_1_OAI21X1_1266 gnd vdd FILL
XDFFPOSX1_647 INVX1_76/A CLKBUF1_54/Y OAI21X1_875/Y gnd vdd DFFPOSX1
XDFFPOSX1_625 INVX1_54/A CLKBUF1_10/Y OAI21X1_853/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_801 gnd vdd FILL
XOAI21X1_1057 BUFX4_354/Y OR2X2_18/B NAND2X1_423/Y gnd OAI21X1_1057/Y vdd OAI21X1
XFILL_1_DFFPOSX1_856 gnd vdd FILL
XFILL_1_DFFPOSX1_834 gnd vdd FILL
XFILL_1_OAI21X1_1299 gnd vdd FILL
XFILL_1_OAI21X1_1288 gnd vdd FILL
XFILL_1_DFFPOSX1_867 gnd vdd FILL
XFILL_1_OAI21X1_206 gnd vdd FILL
XFILL_1_OAI21X1_1277 gnd vdd FILL
XFILL_1_DFFPOSX1_845 gnd vdd FILL
XFILL_1_OAI21X1_217 gnd vdd FILL
XDFFPOSX1_658 BUFX2_295/A CLKBUF1_52/Y OAI21X1_886/Y gnd vdd DFFPOSX1
XDFFPOSX1_669 BUFX2_307/A CLKBUF1_81/Y OAI21X1_897/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_228 gnd vdd FILL
XFILL_1_DFFPOSX1_889 gnd vdd FILL
XFILL_1_DFFPOSX1_878 gnd vdd FILL
XFILL_1_OAI21X1_239 gnd vdd FILL
XNAND2X1_717 BUFX2_789/A BUFX4_373/Y gnd NAND2X1_717/Y vdd NAND2X1
XNAND2X1_728 BUFX2_782/A BUFX4_320/Y gnd NAND2X1_728/Y vdd NAND2X1
XNAND2X1_706 BUFX2_698/A BUFX4_192/Y gnd NAND2X1_706/Y vdd NAND2X1
XNAND2X1_739 BUFX2_794/A BUFX4_361/Y gnd NAND2X1_739/Y vdd NAND2X1
XFILL_6_DFFPOSX1_471 gnd vdd FILL
XFILL_6_DFFPOSX1_460 gnd vdd FILL
XFILL_9_12_1 gnd vdd FILL
XFILL_1_NAND2X1_223 gnd vdd FILL
XFILL_1_NAND2X1_201 gnd vdd FILL
XFILL_1_NAND2X1_212 gnd vdd FILL
XFILL_0_DFFPOSX1_413 gnd vdd FILL
XFILL_1_NAND2X1_234 gnd vdd FILL
XFILL_0_DFFPOSX1_402 gnd vdd FILL
XFILL_0_DFFPOSX1_424 gnd vdd FILL
XFILL_1_NAND2X1_245 gnd vdd FILL
XFILL_0_DFFPOSX1_457 gnd vdd FILL
XFILL_1_NAND2X1_289 gnd vdd FILL
XFILL_1_NAND2X1_267 gnd vdd FILL
XFILL_1_NAND2X1_278 gnd vdd FILL
XFILL_0_DFFPOSX1_435 gnd vdd FILL
XFILL_0_DFFPOSX1_446 gnd vdd FILL
XFILL_0_DFFPOSX1_479 gnd vdd FILL
XFILL_0_DFFPOSX1_468 gnd vdd FILL
XFILL_3_DFFPOSX1_939 gnd vdd FILL
XFILL_3_DFFPOSX1_906 gnd vdd FILL
XFILL_3_DFFPOSX1_917 gnd vdd FILL
XFILL_3_DFFPOSX1_928 gnd vdd FILL
XDFFPOSX1_51 BUFX2_720/A CLKBUF1_89/Y DFFPOSX1_51/D gnd vdd DFFPOSX1
XDFFPOSX1_62 BUFX2_732/A CLKBUF1_8/Y DFFPOSX1_62/D gnd vdd DFFPOSX1
XDFFPOSX1_40 BUFX2_739/A CLKBUF1_87/Y DFFPOSX1_40/D gnd vdd DFFPOSX1
XDFFPOSX1_84 BUFX2_753/A CLKBUF1_101/Y DFFPOSX1_84/D gnd vdd DFFPOSX1
XOAI21X1_1591 BUFX4_349/Y INVX2_127/Y NAND2X1_660/Y gnd OAI21X1_1591/Y vdd OAI21X1
XDFFPOSX1_95 BUFX2_765/A CLKBUF1_102/Y DFFPOSX1_95/D gnd vdd DFFPOSX1
XOAI21X1_1580 INVX2_113/Y INVX8_2/A OAI21X1_1580/C gnd OAI21X1_1580/Y vdd OAI21X1
XDFFPOSX1_73 BUFX2_772/A CLKBUF1_58/Y DFFPOSX1_73/D gnd vdd DFFPOSX1
XFILL_2_OAI21X1_900 gnd vdd FILL
XFILL_2_OAI21X1_933 gnd vdd FILL
XFILL_1_OAI21X1_762 gnd vdd FILL
XFILL_0_OAI21X1_580 gnd vdd FILL
XFILL_1_OAI21X1_773 gnd vdd FILL
XFILL_1_OAI21X1_740 gnd vdd FILL
XFILL_0_OAI21X1_591 gnd vdd FILL
XFILL_1_OAI21X1_751 gnd vdd FILL
XBUFX4_29 BUFX4_82/A gnd BUFX4_29/Y vdd BUFX4
XFILL_1_OAI21X1_795 gnd vdd FILL
XBUFX4_18 INVX8_6/Y gnd BUFX4_18/Y vdd BUFX4
XFILL_1_OAI21X1_784 gnd vdd FILL
XFILL_15_18_1 gnd vdd FILL
XBUFX2_616 BUFX2_616/A gnd majID4_o[26] vdd BUFX2
XBUFX2_605 BUFX2_605/A gnd majID4_o[36] vdd BUFX2
XBUFX2_627 BUFX2_627/A gnd majID4_o[16] vdd BUFX2
XFILL_2_DFFPOSX1_529 gnd vdd FILL
XFILL_2_DFFPOSX1_507 gnd vdd FILL
XFILL_2_DFFPOSX1_518 gnd vdd FILL
XBUFX2_649 BUFX2_649/A gnd pid1_o[31] vdd BUFX2
XBUFX2_638 BUFX2_638/A gnd majID4_o[6] vdd BUFX2
XFILL_0_CLKBUF1_91 gnd vdd FILL
XFILL_0_CLKBUF1_80 gnd vdd FILL
XFILL_0_OAI21X1_1390 gnd vdd FILL
XFILL_0_DFFPOSX1_980 gnd vdd FILL
XFILL_0_DFFPOSX1_991 gnd vdd FILL
XFILL_0_BUFX2_301 gnd vdd FILL
XFILL_0_BUFX2_323 gnd vdd FILL
XINVX2_112 INVX2_112/A gnd INVX2_112/Y vdd INVX2
XINVX2_101 NOR3X1_16/B gnd INVX2_101/Y vdd INVX2
XFILL_0_BUFX2_312 gnd vdd FILL
XINVX2_123 bundlePid_i[25] gnd INVX2_123/Y vdd INVX2
XINVX2_134 bundlePid_i[14] gnd INVX2_134/Y vdd INVX2
XINVX2_145 bundlePid_i[3] gnd INVX2_145/Y vdd INVX2
XFILL_1_DFFPOSX1_119 gnd vdd FILL
XFILL_0_BUFX2_345 gnd vdd FILL
XFILL_0_BUFX2_334 gnd vdd FILL
XFILL_0_BUFX2_356 gnd vdd FILL
XINVX2_156 bundleTid_i[53] gnd INVX2_156/Y vdd INVX2
XFILL_1_DFFPOSX1_108 gnd vdd FILL
XINVX2_189 bundleTid_i[20] gnd INVX2_189/Y vdd INVX2
XFILL_0_BUFX2_378 gnd vdd FILL
XINVX2_167 bundleTid_i[42] gnd INVX2_167/Y vdd INVX2
XFILL_0_BUFX2_389 gnd vdd FILL
XINVX2_178 bundleTid_i[31] gnd INVX2_178/Y vdd INVX2
XFILL_0_BUFX2_367 gnd vdd FILL
XFILL_14_13_0 gnd vdd FILL
XFILL_2_OAI21X1_1440 gnd vdd FILL
XFILL_34_5_0 gnd vdd FILL
XFILL_22_1 gnd vdd FILL
XOAI21X1_508 INVX1_25/Y OAI21X1_508/B OAI21X1_508/C gnd OAI21X1_508/Y vdd OAI21X1
XOAI21X1_519 NOR2X1_4/B INVX4_29/Y OAI21X1_519/C gnd OAI21X1_521/A vdd OAI21X1
XFILL_1_NAND3X1_30 gnd vdd FILL
XFILL_1_OAI21X1_1030 gnd vdd FILL
XFILL_1_NAND3X1_63 gnd vdd FILL
XFILL_1_OAI21X1_1041 gnd vdd FILL
XFILL_1_NAND3X1_52 gnd vdd FILL
XFILL_1_NAND3X1_41 gnd vdd FILL
XDFFPOSX1_422 BUFX2_469/A CLKBUF1_45/Y OAI21X1_396/Y gnd vdd DFFPOSX1
XDFFPOSX1_400 BUFX2_432/A CLKBUF1_90/Y OAI21X1_372/Y gnd vdd DFFPOSX1
XDFFPOSX1_411 BUFX2_444/A CLKBUF1_6/Y OAI21X1_383/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1052 gnd vdd FILL
XFILL_1_OAI21X1_1063 gnd vdd FILL
XFILL_1_DFFPOSX1_642 gnd vdd FILL
XFILL_1_DFFPOSX1_620 gnd vdd FILL
XFILL_1_DFFPOSX1_631 gnd vdd FILL
XDFFPOSX1_433 BUFX2_462/A CLKBUF1_13/Y OAI21X1_420/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1074 gnd vdd FILL
XDFFPOSX1_455 BUFX2_486/A CLKBUF1_44/Y OAI21X1_453/Y gnd vdd DFFPOSX1
XDFFPOSX1_444 BUFX2_474/A CLKBUF1_15/Y OAI21X1_436/Y gnd vdd DFFPOSX1
XFILL_38_18_1 gnd vdd FILL
XFILL_0_BUFX2_890 gnd vdd FILL
XFILL_1_DFFPOSX1_664 gnd vdd FILL
XFILL_1_OAI21X1_1085 gnd vdd FILL
XDFFPOSX1_477 BUFX2_510/A CLKBUF1_9/Y OAI21X1_489/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1096 gnd vdd FILL
XDFFPOSX1_499 BUFX2_528/A CLKBUF1_90/Y OAI21X1_543/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_675 gnd vdd FILL
XFILL_1_DFFPOSX1_653 gnd vdd FILL
XDFFPOSX1_466 BUFX2_498/A CLKBUF1_48/Y OAI21X1_469/Y gnd vdd DFFPOSX1
XNAND2X1_503 BUFX2_75/A BUFX4_228/Y gnd NAND2X1_503/Y vdd NAND2X1
XDFFPOSX1_488 BUFX2_555/A CLKBUF1_66/Y OAI21X1_512/Y gnd vdd DFFPOSX1
XNAND2X1_525 BUFX2_87/A BUFX4_202/Y gnd NAND2X1_525/Y vdd NAND2X1
XFILL_19_12_0 gnd vdd FILL
XFILL_2_OAI21X1_207 gnd vdd FILL
XNAND2X1_514 bundleAddress_i[41] bundleAddress_i[40] gnd INVX1_202/A vdd NAND2X1
XNAND2X1_536 bundleAddress_i[29] bundleAddress_i[28] gnd NOR2X1_154/A vdd NAND2X1
XFILL_1_DFFPOSX1_697 gnd vdd FILL
XFILL_1_DFFPOSX1_686 gnd vdd FILL
XNAND2X1_558 BUFX2_106/A BUFX4_187/Y gnd NAND2X1_558/Y vdd NAND2X1
XNAND2X1_547 BUFX4_239/Y NAND2X1_547/B gnd NAND2X1_547/Y vdd NAND2X1
XNAND2X1_569 BUFX2_112/A BUFX4_201/Y gnd NAND2X1_569/Y vdd NAND2X1
XFILL_32_14_0 gnd vdd FILL
XFILL_0_AND2X2_15 gnd vdd FILL
XFILL_0_AND2X2_26 gnd vdd FILL
XFILL_25_5_0 gnd vdd FILL
XFILL_0_5_0 gnd vdd FILL
XFILL_0_DFFPOSX1_232 gnd vdd FILL
XFILL_0_DFFPOSX1_221 gnd vdd FILL
XFILL_0_DFFPOSX1_210 gnd vdd FILL
XFILL_0_DFFPOSX1_254 gnd vdd FILL
XFILL_0_DFFPOSX1_243 gnd vdd FILL
XFILL_0_DFFPOSX1_265 gnd vdd FILL
XFILL_0_DFFPOSX1_276 gnd vdd FILL
XFILL_0_DFFPOSX1_298 gnd vdd FILL
XFILL_0_DFFPOSX1_287 gnd vdd FILL
XFILL_3_DFFPOSX1_714 gnd vdd FILL
XFILL_3_DFFPOSX1_703 gnd vdd FILL
XFILL_3_DFFPOSX1_747 gnd vdd FILL
XFILL_3_DFFPOSX1_725 gnd vdd FILL
XFILL_3_DFFPOSX1_736 gnd vdd FILL
XFILL_3_CLKBUF1_24 gnd vdd FILL
XFILL_3_CLKBUF1_13 gnd vdd FILL
XFILL_3_DFFPOSX1_758 gnd vdd FILL
XFILL_3_CLKBUF1_57 gnd vdd FILL
XFILL_3_CLKBUF1_35 gnd vdd FILL
XFILL_3_DFFPOSX1_769 gnd vdd FILL
XFILL_3_CLKBUF1_46 gnd vdd FILL
XFILL_3_CLKBUF1_68 gnd vdd FILL
XFILL_3_CLKBUF1_79 gnd vdd FILL
XFILL_37_13_0 gnd vdd FILL
XFILL_1_NOR2X1_120 gnd vdd FILL
XFILL_8_6_0 gnd vdd FILL
XFILL_1_NOR2X1_142 gnd vdd FILL
XFILL_1_OAI21X1_570 gnd vdd FILL
XFILL_1_OAI21X1_581 gnd vdd FILL
XFILL_1_NOR2X1_153 gnd vdd FILL
XFILL_2_OAI21X1_752 gnd vdd FILL
XFILL_2_NAND3X1_6 gnd vdd FILL
XFILL_1_NOR2X1_175 gnd vdd FILL
XFILL_1_NOR2X1_197 gnd vdd FILL
XFILL_1_OAI21X1_592 gnd vdd FILL
XFILL_2_DFFPOSX1_304 gnd vdd FILL
XBUFX2_402 BUFX2_402/A gnd majID1_o[46] vdd BUFX2
XFILL_2_DFFPOSX1_337 gnd vdd FILL
XFILL_2_DFFPOSX1_326 gnd vdd FILL
XFILL_2_DFFPOSX1_315 gnd vdd FILL
XBUFX2_435 BUFX2_435/A gnd majID1_o[16] vdd BUFX2
XBUFX2_413 BUFX2_413/A gnd majID1_o[36] vdd BUFX2
XBUFX2_424 BUFX2_424/A gnd majID1_o[26] vdd BUFX2
XFILL_2_DFFPOSX1_348 gnd vdd FILL
XBUFX2_446 BUFX2_446/A gnd majID1_o[6] vdd BUFX2
XBUFX2_468 BUFX2_468/A gnd majID2_o[44] vdd BUFX2
XFILL_16_5_0 gnd vdd FILL
XFILL_2_DFFPOSX1_359 gnd vdd FILL
XBUFX2_457 BUFX2_457/A gnd majID2_o[63] vdd BUFX2
XBUFX2_479 BUFX2_479/A gnd majID2_o[34] vdd BUFX2
XFILL_5_DFFPOSX1_808 gnd vdd FILL
XFILL_1_BUFX4_340 gnd vdd FILL
XFILL_5_DFFPOSX1_819 gnd vdd FILL
XFILL_1_BUFX4_351 gnd vdd FILL
XFILL_1_BUFX4_362 gnd vdd FILL
XFILL_1_BUFX4_373 gnd vdd FILL
XFILL_1_BUFX4_384 gnd vdd FILL
XFILL_0_BUFX2_131 gnd vdd FILL
XFILL_0_BUFX2_120 gnd vdd FILL
XFILL_2_OAI21X1_97 gnd vdd FILL
XFILL_0_BUFX2_153 gnd vdd FILL
XFILL_0_BUFX2_164 gnd vdd FILL
XFILL_0_BUFX2_142 gnd vdd FILL
XFILL_0_BUFX2_197 gnd vdd FILL
XFILL_0_BUFX2_186 gnd vdd FILL
XFILL_0_BUFX2_175 gnd vdd FILL
XFILL_1_DFFPOSX1_7 gnd vdd FILL
XFILL_4_DFFPOSX1_409 gnd vdd FILL
XFILL_2_OAI21X1_1292 gnd vdd FILL
XFILL_2_DFFPOSX1_860 gnd vdd FILL
XBUFX2_980 BUFX2_980/A gnd tid4_o[44] vdd BUFX2
XFILL_2_DFFPOSX1_882 gnd vdd FILL
XBUFX2_991 BUFX2_991/A gnd tid4_o[34] vdd BUFX2
XFILL_2_DFFPOSX1_871 gnd vdd FILL
XFILL_2_DFFPOSX1_893 gnd vdd FILL
XOAI21X1_305 INVX2_198/Y BUFX4_295/Y OAI21X1_305/C gnd OAI21X1_305/Y vdd OAI21X1
XOAI21X1_338 BUFX4_388/Y INVX2_15/Y NAND2X1_82/Y gnd OAI21X1_338/Y vdd OAI21X1
XOAI21X1_327 INVX2_7/Y BUFX4_303/Y OAI21X1_327/C gnd OAI21X1_327/Y vdd OAI21X1
XOAI21X1_316 BUFX4_131/Y BUFX4_30/Y BUFX2_1023/A gnd OAI21X1_317/C vdd OAI21X1
XOAI21X1_349 BUFX4_337/Y INVX4_8/Y NAND2X1_93/Y gnd OAI21X1_349/Y vdd OAI21X1
XFILL_21_11_1 gnd vdd FILL
XBUFX4_3 BUFX4_3/A gnd BUFX4_3/Y vdd BUFX4
XDFFPOSX1_230 BUFX2_917/A CLKBUF1_92/Y OAI21X1_77/Y gnd vdd DFFPOSX1
XDFFPOSX1_252 BUFX2_922/A CLKBUF1_43/Y OAI21X1_121/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_450 gnd vdd FILL
XDFFPOSX1_263 BUFX2_934/A CLKBUF1_73/Y OAI21X1_143/Y gnd vdd DFFPOSX1
XDFFPOSX1_241 BUFX2_910/A CLKBUF1_10/Y OAI21X1_99/Y gnd vdd DFFPOSX1
XDFFPOSX1_296 BUFX2_1003/A CLKBUF1_59/Y OAI21X1_209/Y gnd vdd DFFPOSX1
XDFFPOSX1_285 BUFX2_958/A CLKBUF1_43/Y OAI21X1_187/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_483 gnd vdd FILL
XFILL_1_DFFPOSX1_461 gnd vdd FILL
XNAND2X1_300 INVX2_46/A NOR2X1_95/Y gnd OAI21X1_639/A vdd NAND2X1
XDFFPOSX1_274 BUFX2_946/A CLKBUF1_4/Y OAI21X1_165/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_472 gnd vdd FILL
XNAND2X1_311 NOR2X1_5/A NOR2X1_105/A gnd NAND2X1_312/A vdd NAND2X1
XNAND2X1_333 OAI21X1_822/Y XNOR2X1_55/A gnd OAI21X1_824/A vdd NAND2X1
XFILL_3_NOR3X1_16 gnd vdd FILL
XNAND2X1_322 NOR2X1_19/Y INVX1_38/A gnd XNOR2X1_47/A vdd NAND2X1
XNAND2X1_344 INVX8_4/A bundle_i[25] gnd OAI21X1_850/C vdd NAND2X1
XFILL_1_DFFPOSX1_494 gnd vdd FILL
XNAND2X1_377 BUFX2_322/A BUFX4_184/Y gnd OAI21X1_883/C vdd NAND2X1
XNAND2X1_355 BUFX4_265/Y bundle_i[14] gnd OAI21X1_861/C vdd NAND2X1
XFILL_4_DFFPOSX1_932 gnd vdd FILL
XFILL_4_DFFPOSX1_921 gnd vdd FILL
XFILL_4_DFFPOSX1_910 gnd vdd FILL
XNAND2X1_366 BUFX4_262/Y bundle_i[3] gnd OAI21X1_872/C vdd NAND2X1
XFILL_4_DFFPOSX1_954 gnd vdd FILL
XFILL_4_DFFPOSX1_943 gnd vdd FILL
XFILL_4_DFFPOSX1_965 gnd vdd FILL
XNAND2X1_399 BUFX2_315/A BUFX4_189/Y gnd OAI21X1_905/C vdd NAND2X1
XNAND2X1_388 BUFX2_303/A BUFX4_206/Y gnd OAI21X1_894/C vdd NAND2X1
XFILL_0_INVX1_109 gnd vdd FILL
XFILL_4_DFFPOSX1_998 gnd vdd FILL
XFILL_4_DFFPOSX1_987 gnd vdd FILL
XFILL_4_DFFPOSX1_976 gnd vdd FILL
XFILL_1_BUFX2_811 gnd vdd FILL
XFILL_1_BUFX2_822 gnd vdd FILL
XFILL_1_BUFX2_855 gnd vdd FILL
XFILL_26_10_1 gnd vdd FILL
XINVX4_3 bundleStartMajId_i[54] gnd INVX4_3/Y vdd INVX4
XFILL_1_INVX2_77 gnd vdd FILL
XFILL_1_BUFX2_877 gnd vdd FILL
XFILL_1_BUFX2_866 gnd vdd FILL
XFILL_2_NOR3X1_8 gnd vdd FILL
XOAI21X1_850 INVX1_51/Y INVX8_4/A OAI21X1_850/C gnd OAI21X1_850/Y vdd OAI21X1
XFILL_3_DFFPOSX1_500 gnd vdd FILL
XFILL_3_DFFPOSX1_522 gnd vdd FILL
XFILL_3_DFFPOSX1_511 gnd vdd FILL
XOAI21X1_883 INVX1_84/Y BUFX4_184/Y OAI21X1_883/C gnd OAI21X1_883/Y vdd OAI21X1
XFILL_3_DFFPOSX1_544 gnd vdd FILL
XOAI21X1_861 INVX1_62/Y BUFX4_265/Y OAI21X1_861/C gnd OAI21X1_861/Y vdd OAI21X1
XFILL_1_BUFX2_899 gnd vdd FILL
XFILL_3_DFFPOSX1_555 gnd vdd FILL
XFILL_3_DFFPOSX1_533 gnd vdd FILL
XOAI21X1_872 INVX1_73/Y BUFX4_262/Y OAI21X1_872/C gnd OAI21X1_872/Y vdd OAI21X1
XOAI21X1_894 INVX1_95/Y BUFX4_206/Y OAI21X1_894/C gnd OAI21X1_894/Y vdd OAI21X1
XFILL_3_DFFPOSX1_588 gnd vdd FILL
XFILL_3_DFFPOSX1_566 gnd vdd FILL
XFILL_3_DFFPOSX1_577 gnd vdd FILL
XFILL_3_DFFPOSX1_599 gnd vdd FILL
XFILL_2_OAI21X1_582 gnd vdd FILL
XFILL_2_DFFPOSX1_112 gnd vdd FILL
XFILL_0_NAND2X1_607 gnd vdd FILL
XBUFX2_210 BUFX2_210/A gnd addr4_o[39] vdd BUFX2
XFILL_2_DFFPOSX1_101 gnd vdd FILL
XFILL_2_DFFPOSX1_134 gnd vdd FILL
XFILL_2_DFFPOSX1_145 gnd vdd FILL
XBUFX2_232 BUFX2_232/A gnd addr4_o[19] vdd BUFX2
XFILL_2_DFFPOSX1_123 gnd vdd FILL
XFILL_0_NAND2X1_618 gnd vdd FILL
XFILL_0_NAND3X1_60 gnd vdd FILL
XFILL_0_NAND2X1_629 gnd vdd FILL
XBUFX2_221 BUFX2_221/A gnd addr4_o[29] vdd BUFX2
XFILL_1_11_1 gnd vdd FILL
XBUFX2_243 BUFX2_243/A gnd addr4_o[9] vdd BUFX2
XFILL_2_DFFPOSX1_178 gnd vdd FILL
XFILL_2_DFFPOSX1_156 gnd vdd FILL
XFILL_2_DFFPOSX1_189 gnd vdd FILL
XBUFX2_254 BUFX2_254/A gnd addr4_o[56] vdd BUFX2
XBUFX2_276 INVX1_67/A gnd instr1_o[9] vdd BUFX2
XBUFX2_265 INVX1_57/A gnd instr1_o[19] vdd BUFX2
XBUFX2_287 INVX1_49/A gnd instr1_o[27] vdd BUFX2
XFILL_2_DFFPOSX1_167 gnd vdd FILL
XFILL_32_8_1 gnd vdd FILL
XBUFX2_298 BUFX2_298/A gnd instr2_o[18] vdd BUFX2
XFILL_31_3_0 gnd vdd FILL
XFILL_28_18_0 gnd vdd FILL
XFILL_5_DFFPOSX1_627 gnd vdd FILL
XFILL_5_DFFPOSX1_605 gnd vdd FILL
XFILL_5_DFFPOSX1_616 gnd vdd FILL
XFILL_1_BUFX4_170 gnd vdd FILL
XFILL_5_DFFPOSX1_649 gnd vdd FILL
XFILL_5_DFFPOSX1_638 gnd vdd FILL
XFILL_1_BUFX4_181 gnd vdd FILL
XFILL_1_BUFX4_192 gnd vdd FILL
XFILL_4_DFFPOSX1_217 gnd vdd FILL
XNAND3X1_6 AND2X2_7/A NOR2X1_11/Y NOR2X1_30/Y gnd NOR2X1_33/B vdd NAND3X1
XFILL_4_DFFPOSX1_206 gnd vdd FILL
XFILL_4_DFFPOSX1_239 gnd vdd FILL
XFILL_4_DFFPOSX1_228 gnd vdd FILL
XFILL_6_10_1 gnd vdd FILL
XFILL_2_CLKBUF1_32 gnd vdd FILL
XFILL_2_CLKBUF1_21 gnd vdd FILL
XFILL_2_CLKBUF1_10 gnd vdd FILL
XFILL_2_CLKBUF1_65 gnd vdd FILL
XFILL_2_CLKBUF1_43 gnd vdd FILL
XFILL_2_CLKBUF1_54 gnd vdd FILL
XFILL_2_CLKBUF1_98 gnd vdd FILL
XFILL_2_CLKBUF1_87 gnd vdd FILL
XFILL_2_CLKBUF1_76 gnd vdd FILL
XFILL_2_DFFPOSX1_690 gnd vdd FILL
XFILL_23_8_1 gnd vdd FILL
XFILL_1_BUFX2_107 gnd vdd FILL
XFILL_22_3_0 gnd vdd FILL
XOAI21X1_102 BUFX4_112/Y BUFX4_353/Y BUFX2_912/A gnd OAI21X1_103/C vdd OAI21X1
XOAI21X1_113 BUFX4_150/Y INVX2_166/Y OAI21X1_113/C gnd OAI21X1_113/Y vdd OAI21X1
XFILL_0_NOR2X1_150 gnd vdd FILL
XFILL_0_NOR2X1_161 gnd vdd FILL
XFILL_0_NOR2X1_172 gnd vdd FILL
XOAI21X1_124 BUFX4_4/A BUFX4_363/Y BUFX2_924/A gnd OAI21X1_125/C vdd OAI21X1
XFILL_0_NOR2X1_183 gnd vdd FILL
XOAI21X1_146 BUFX4_3/Y BUFX4_356/Y BUFX2_936/A gnd OAI21X1_147/C vdd OAI21X1
XOAI21X1_135 BUFX4_125/Y INVX2_177/Y OAI21X1_135/C gnd OAI21X1_135/Y vdd OAI21X1
XFILL_0_NOR2X1_194 gnd vdd FILL
XFILL_0_DFFPOSX1_1002 gnd vdd FILL
XFILL_0_DFFPOSX1_1013 gnd vdd FILL
XOAI21X1_179 BUFX4_178/Y INVX2_199/Y OAI21X1_179/C gnd OAI21X1_179/Y vdd OAI21X1
XOAI21X1_168 BUFX4_97/Y BUFX4_377/Y BUFX2_948/A gnd OAI21X1_169/C vdd OAI21X1
XFILL_0_DFFPOSX1_1024 gnd vdd FILL
XOAI21X1_157 BUFX4_124/Y INVX2_188/Y OAI21X1_157/C gnd OAI21X1_157/Y vdd OAI21X1
XFILL_1_DFFPOSX1_291 gnd vdd FILL
XFILL_1_DFFPOSX1_280 gnd vdd FILL
XNAND2X1_130 BUFX2_447/A BUFX4_328/Y gnd OAI21X1_386/C vdd NAND2X1
XNAND2X1_141 bundleStartMajId_i[61] bundleStartMajId_i[60] gnd NOR2X1_3/B vdd NAND2X1
XNAND2X1_152 BUFX2_518/A BUFX4_199/Y gnd OAI21X1_409/C vdd NAND2X1
XFILL_8_18_0 gnd vdd FILL
XFILL_4_DFFPOSX1_740 gnd vdd FILL
XFILL_0_XNOR2X1_17 gnd vdd FILL
XNAND2X1_174 bundleStartMajId_i[44] NOR2X1_12/Y gnd NAND2X1_177/B vdd NAND2X1
XNAND2X1_163 BUFX2_463/A BUFX4_215/Y gnd OAI21X1_421/C vdd NAND2X1
XFILL_5_4_0 gnd vdd FILL
XNAND2X1_185 bundleStartMajId_i[41] AND2X2_3/Y gnd XNOR2X1_9/A vdd NAND2X1
XFILL_6_9_1 gnd vdd FILL
XNAND2X1_196 XNOR2X1_11/A OAI21X1_442/Y gnd OAI21X1_443/A vdd NAND2X1
XFILL_4_DFFPOSX1_751 gnd vdd FILL
XFILL_1_OAI21X1_61 gnd vdd FILL
XFILL_4_DFFPOSX1_773 gnd vdd FILL
XFILL_4_DFFPOSX1_762 gnd vdd FILL
XFILL_0_XNOR2X1_39 gnd vdd FILL
XFILL_0_XNOR2X1_28 gnd vdd FILL
XFILL_1_OAI21X1_50 gnd vdd FILL
XFILL_1_OAI21X1_94 gnd vdd FILL
XFILL_1_OAI21X1_72 gnd vdd FILL
XFILL_12_16_1 gnd vdd FILL
XFILL_4_DFFPOSX1_784 gnd vdd FILL
XFILL_1_OAI21X1_83 gnd vdd FILL
XFILL_4_DFFPOSX1_795 gnd vdd FILL
XFILL_14_8_1 gnd vdd FILL
XFILL_0_DFFPOSX1_4 gnd vdd FILL
XFILL_13_3_0 gnd vdd FILL
XFILL_1_BUFX2_630 gnd vdd FILL
XFILL_1_BUFX2_663 gnd vdd FILL
XFILL_1_BUFX2_652 gnd vdd FILL
XFILL_0_BUFX4_204 gnd vdd FILL
XFILL_0_BUFX4_215 gnd vdd FILL
XFILL_3_DFFPOSX1_330 gnd vdd FILL
XFILL_0_BUFX4_248 gnd vdd FILL
XOAI21X1_1409 INVX1_219/Y INVX2_61/Y INVX2_62/Y gnd OAI21X1_1410/C vdd OAI21X1
XFILL_0_BUFX4_237 gnd vdd FILL
XFILL_1_BUFX2_674 gnd vdd FILL
XFILL_0_BUFX4_226 gnd vdd FILL
XFILL_1_OAI21X1_1629 gnd vdd FILL
XFILL_1_OAI21X1_1607 gnd vdd FILL
XFILL_3_DFFPOSX1_341 gnd vdd FILL
XOAI21X1_680 BUFX4_145/Y BUFX4_37/Y BUFX2_646/A gnd OAI21X1_681/C vdd OAI21X1
XFILL_0_BUFX4_259 gnd vdd FILL
XFILL_1_OAI21X1_1618 gnd vdd FILL
XNOR3X1_9 NOR3X1_9/A NOR3X1_9/B NOR3X1_9/C gnd NOR3X1_9/Y vdd NOR3X1
XOAI21X1_691 BUFX4_176/Y BUFX4_81/Y BUFX2_588/A gnd OAI21X1_692/C vdd OAI21X1
XFILL_3_DFFPOSX1_352 gnd vdd FILL
XFILL_3_DFFPOSX1_363 gnd vdd FILL
XFILL_3_DFFPOSX1_374 gnd vdd FILL
XFILL_3_DFFPOSX1_396 gnd vdd FILL
XFILL_3_DFFPOSX1_385 gnd vdd FILL
XFILL_0_OAI21X1_409 gnd vdd FILL
XFILL_0_INVX4_12 gnd vdd FILL
XFILL_3_DFFPOSX1_1006 gnd vdd FILL
XFILL_0_INVX4_34 gnd vdd FILL
XFILL_0_INVX4_23 gnd vdd FILL
XFILL_6_DFFPOSX1_845 gnd vdd FILL
XFILL_0_INVX4_45 gnd vdd FILL
XFILL_3_DFFPOSX1_1017 gnd vdd FILL
XFILL_6_DFFPOSX1_878 gnd vdd FILL
XFILL_6_DFFPOSX1_856 gnd vdd FILL
XFILL_17_15_1 gnd vdd FILL
XFILL_6_DFFPOSX1_867 gnd vdd FILL
XFILL_3_DFFPOSX1_1028 gnd vdd FILL
XXNOR2X1_41 INVX1_35/A INVX4_3/Y gnd XNOR2X1_41/Y vdd XNOR2X1
XFILL_5_3 gnd vdd FILL
XXNOR2X1_30 NOR2X1_68/Y bundleStartMajId_i[40] gnd XNOR2X1_30/Y vdd XNOR2X1
XXNOR2X1_74 INVX2_93/A bundleAddress_i[54] gnd XNOR2X1_74/Y vdd XNOR2X1
XFILL_6_DFFPOSX1_889 gnd vdd FILL
XXNOR2X1_63 XNOR2X1_63/A INVX4_37/Y gnd XNOR2X1_63/Y vdd XNOR2X1
XXNOR2X1_52 INVX4_31/A bundleStartMajId_i[22] gnd XNOR2X1_52/Y vdd XNOR2X1
XXNOR2X1_85 XNOR2X1_85/A bundleAddress_i[18] gnd XNOR2X1_85/Y vdd XNOR2X1
XXNOR2X1_96 XNOR2X1_96/A bundleAddress_i[39] gnd XNOR2X1_96/Y vdd XNOR2X1
XFILL_0_NAND2X1_404 gnd vdd FILL
XFILL_0_NAND2X1_415 gnd vdd FILL
XFILL_30_17_1 gnd vdd FILL
XFILL_1_XNOR2X1_8 gnd vdd FILL
XFILL_0_NAND2X1_426 gnd vdd FILL
XBUFX2_62 BUFX2_62/A gnd addr1_o[56] vdd BUFX2
XFILL_0_OAI21X1_1208 gnd vdd FILL
XBUFX2_40 BUFX2_40/A gnd addr1_o[19] vdd BUFX2
XFILL_0_OAI21X1_1219 gnd vdd FILL
XFILL_0_NAND2X1_448 gnd vdd FILL
XFILL_1_NAND2X1_608 gnd vdd FILL
XFILL_11_11_0 gnd vdd FILL
XFILL_0_NAND2X1_437 gnd vdd FILL
XFILL_0_NAND2X1_459 gnd vdd FILL
XBUFX2_51 BUFX2_51/A gnd addr1_o[9] vdd BUFX2
XBUFX2_73 BUFX2_73/A gnd addr2_o[47] vdd BUFX2
XBUFX2_84 BUFX2_84/A gnd addr2_o[37] vdd BUFX2
XFILL_0_DFFPOSX1_809 gnd vdd FILL
XBUFX2_95 BUFX2_95/A gnd addr2_o[27] vdd BUFX2
XFILL_5_DFFPOSX1_402 gnd vdd FILL
XFILL_5_DFFPOSX1_413 gnd vdd FILL
XFILL_5_DFFPOSX1_424 gnd vdd FILL
XFILL_5_DFFPOSX1_435 gnd vdd FILL
XFILL_5_DFFPOSX1_479 gnd vdd FILL
XFILL_5_DFFPOSX1_468 gnd vdd FILL
XFILL_5_DFFPOSX1_457 gnd vdd FILL
XFILL_5_DFFPOSX1_446 gnd vdd FILL
XFILL_1_BUFX4_40 gnd vdd FILL
XFILL_1_BUFX4_62 gnd vdd FILL
XFILL_1_BUFX4_51 gnd vdd FILL
XFILL_1_BUFX4_95 gnd vdd FILL
XFILL_1_BUFX4_84 gnd vdd FILL
XFILL_1_BUFX4_73 gnd vdd FILL
XFILL_0_AOI21X1_28 gnd vdd FILL
XFILL_0_AOI21X1_39 gnd vdd FILL
XFILL_0_AOI21X1_17 gnd vdd FILL
XFILL_0_OAI21X1_932 gnd vdd FILL
XFILL_2_CLKBUF1_8 gnd vdd FILL
XFILL_0_OAI21X1_910 gnd vdd FILL
XFILL_0_OAI21X1_921 gnd vdd FILL
XFILL_0_OAI21X1_965 gnd vdd FILL
XFILL_0_OAI21X1_954 gnd vdd FILL
XFILL_0_OAI21X1_943 gnd vdd FILL
XFILL_0_OAI21X1_998 gnd vdd FILL
XFILL_0_OAI21X1_976 gnd vdd FILL
XFILL_0_OAI21X1_987 gnd vdd FILL
XFILL_35_16_1 gnd vdd FILL
XFILL_16_10_0 gnd vdd FILL
XFILL_2_BUFX4_124 gnd vdd FILL
XFILL_2_BUFX4_157 gnd vdd FILL
XFILL_1_OR2X2_21 gnd vdd FILL
XFILL_1_OR2X2_10 gnd vdd FILL
XFILL_0_OAI21X1_1742 gnd vdd FILL
XFILL_0_OAI21X1_1731 gnd vdd FILL
XFILL_0_OAI21X1_1720 gnd vdd FILL
XFILL_0_OAI21X1_1786 gnd vdd FILL
XFILL_0_OAI21X1_1764 gnd vdd FILL
XFILL_0_OAI21X1_1753 gnd vdd FILL
XFILL_0_OAI21X1_1775 gnd vdd FILL
XFILL_0_OAI21X1_1797 gnd vdd FILL
XFILL_5_DFFPOSX1_980 gnd vdd FILL
XFILL_5_DFFPOSX1_991 gnd vdd FILL
XFILL_0_NOR2X1_15 gnd vdd FILL
XFILL_0_BUFX2_719 gnd vdd FILL
XAOI21X1_52 bundleAddress_i[18] XNOR2X1_85/A bundleAddress_i[17] gnd AOI21X1_52/Y
+ vdd AOI21X1
XAOI21X1_41 INVX1_195/Y INVX2_102/Y bundleAddress_i[14] gnd AOI21X1_41/Y vdd AOI21X1
XFILL_0_BUFX2_708 gnd vdd FILL
XFILL_0_NOR2X1_37 gnd vdd FILL
XFILL_0_NOR2X1_48 gnd vdd FILL
XAOI21X1_30 bundleStartMajId_i[54] INVX1_35/Y bundleStartMajId_i[53] gnd AOI21X1_30/Y
+ vdd AOI21X1
XFILL_0_NOR2X1_26 gnd vdd FILL
XAOI21X1_63 bundleAddress_i[12] NOR2X1_228/Y bundleAddress_i[11] gnd AOI21X1_63/Y
+ vdd AOI21X1
XFILL_0_NOR2X1_59 gnd vdd FILL
XOAI21X1_3 OAI21X1_4/A INVX2_3/Y OAI21X1_3/C gnd OAI21X1_3/Y vdd OAI21X1
XFILL_34_11_0 gnd vdd FILL
XXNOR2X1_100 INVX1_223/A INVX4_40/Y gnd XNOR2X1_100/Y vdd XNOR2X1
XBUFX4_316 BUFX4_386/A gnd BUFX4_316/Y vdd BUFX4
XBUFX4_305 BUFX4_310/A gnd BUFX4_305/Y vdd BUFX4
XBUFX4_327 BUFX4_388/A gnd OAI21X1_6/A vdd BUFX4
XBUFX4_349 BUFX4_380/A gnd BUFX4_349/Y vdd BUFX4
XFILL_4_DFFPOSX1_570 gnd vdd FILL
XBUFX4_338 BUFX4_384/A gnd OAI21X1_7/A vdd BUFX4
XFILL_4_DFFPOSX1_581 gnd vdd FILL
XFILL_4_DFFPOSX1_592 gnd vdd FILL
XFILL_1_BUFX2_460 gnd vdd FILL
XFILL_1_BUFX2_471 gnd vdd FILL
XOAI21X1_1228 INVX4_47/Y INVX2_60/Y INVX2_61/Y gnd OAI21X1_1229/C vdd OAI21X1
XOAI21X1_1217 NAND2X1_591/Y BUFX4_126/Y OAI21X1_1217/C gnd OAI21X1_1217/Y vdd OAI21X1
XFILL_1_OAI21X1_1415 gnd vdd FILL
XFILL_1_OAI21X1_1404 gnd vdd FILL
XOAI21X1_1206 NOR3X1_15/Y bundleAddress_i[0] BUFX4_243/Y gnd OAI21X1_1207/B vdd OAI21X1
XFILL_1_CLKBUF1_40 gnd vdd FILL
XOAI21X1_1239 INVX2_96/A INVX1_201/A OAI21X1_1239/C gnd OAI21X1_1241/A vdd OAI21X1
XFILL_1_OAI21X1_1437 gnd vdd FILL
XDFFPOSX1_818 BUFX2_67/A CLKBUF1_29/Y OAI21X1_1121/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1426 gnd vdd FILL
XFILL_3_DFFPOSX1_171 gnd vdd FILL
XFILL_3_DFFPOSX1_182 gnd vdd FILL
XDFFPOSX1_807 BUFX2_61/A CLKBUF1_30/Y OAI21X1_1099/Y gnd vdd DFFPOSX1
XFILL_1_CLKBUF1_73 gnd vdd FILL
XFILL_1_INVX8_2 gnd vdd FILL
XFILL_1_OAI21X1_1448 gnd vdd FILL
XFILL_3_DFFPOSX1_160 gnd vdd FILL
XFILL_1_CLKBUF1_51 gnd vdd FILL
XFILL_1_CLKBUF1_62 gnd vdd FILL
XDFFPOSX1_829 BUFX2_79/A CLKBUF1_34/Y OAI21X1_1138/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_228 gnd vdd FILL
XFILL_1_CLKBUF1_95 gnd vdd FILL
XFILL_1_OAI21X1_1459 gnd vdd FILL
XFILL_1_CLKBUF1_84 gnd vdd FILL
XFILL_0_OAI21X1_206 gnd vdd FILL
XFILL_0_OAI21X1_217 gnd vdd FILL
XFILL_3_DFFPOSX1_193 gnd vdd FILL
XFILL_0_OAI21X1_239 gnd vdd FILL
XFILL_6_DFFPOSX1_620 gnd vdd FILL
XFILL_6_DFFPOSX1_642 gnd vdd FILL
XFILL_6_DFFPOSX1_631 gnd vdd FILL
XFILL_6_DFFPOSX1_653 gnd vdd FILL
XFILL_37_7_1 gnd vdd FILL
XFILL_0_NAND2X1_201 gnd vdd FILL
XFILL_36_2_0 gnd vdd FILL
XFILL_1_NAND2X1_405 gnd vdd FILL
XFILL_0_NAND2X1_234 gnd vdd FILL
XFILL_0_NAND2X1_223 gnd vdd FILL
XFILL_0_NAND2X1_212 gnd vdd FILL
XFILL_0_OAI21X1_1005 gnd vdd FILL
XFILL_0_OAI21X1_1038 gnd vdd FILL
XFILL_1_NAND2X1_416 gnd vdd FILL
XFILL_0_NAND2X1_256 gnd vdd FILL
XFILL_0_DFFPOSX1_606 gnd vdd FILL
XFILL_0_NAND2X1_267 gnd vdd FILL
XFILL_0_OAI21X1_1016 gnd vdd FILL
XFILL_0_OAI21X1_1027 gnd vdd FILL
XFILL_0_NAND2X1_245 gnd vdd FILL
XFILL_0_DFFPOSX1_639 gnd vdd FILL
XFILL_0_OAI21X1_1049 gnd vdd FILL
XFILL_1_NAND2X1_449 gnd vdd FILL
XFILL_0_NAND2X1_289 gnd vdd FILL
XFILL_0_DFFPOSX1_617 gnd vdd FILL
XFILL_0_NAND2X1_278 gnd vdd FILL
XFILL_0_DFFPOSX1_628 gnd vdd FILL
XFILL_5_DFFPOSX1_210 gnd vdd FILL
XFILL_5_DFFPOSX1_232 gnd vdd FILL
XFILL_5_DFFPOSX1_254 gnd vdd FILL
XFILL_5_DFFPOSX1_243 gnd vdd FILL
XFILL_5_DFFPOSX1_221 gnd vdd FILL
XFILL_20_6_1 gnd vdd FILL
XFILL_5_DFFPOSX1_276 gnd vdd FILL
XFILL_5_DFFPOSX1_265 gnd vdd FILL
XFILL_5_DFFPOSX1_287 gnd vdd FILL
XFILL_5_DFFPOSX1_298 gnd vdd FILL
XFILL_0_OAI21X1_80 gnd vdd FILL
XFILL_0_OAI21X1_91 gnd vdd FILL
XOAI21X1_1740 BUFX4_170/Y BUFX4_32/Y BUFX2_752/A gnd OAI21X1_1741/C vdd OAI21X1
XOAI21X1_1751 INVX2_137/Y BUFX4_297/Y OAI21X1_1751/C gnd DFFPOSX1_88/D vdd OAI21X1
XOAI21X1_1762 BUFX4_123/Y BUFX4_47/Y BUFX2_764/A gnd OAI21X1_1763/C vdd OAI21X1
XOAI21X1_1784 BUFX4_326/Y INVX2_156/Y NAND2X1_725/Y gnd OAI21X1_1784/Y vdd OAI21X1
XOAI21X1_1773 INVX2_116/Y BUFX4_302/Y OAI21X1_1773/C gnd DFFPOSX1_99/D vdd OAI21X1
XFILL_1_OAI21X1_900 gnd vdd FILL
XOAI21X1_1795 BUFX4_368/Y INVX2_167/Y NAND2X1_736/Y gnd OAI21X1_1795/Y vdd OAI21X1
XFILL_1_OAI21X1_911 gnd vdd FILL
XFILL_1_OAI21X1_922 gnd vdd FILL
XFILL_0_OAI21X1_740 gnd vdd FILL
XFILL_1_OAI21X1_944 gnd vdd FILL
XFILL_1_OAI21X1_933 gnd vdd FILL
XFILL_0_OAI21X1_762 gnd vdd FILL
XFILL_0_OAI21X1_784 gnd vdd FILL
XFILL_0_OAI21X1_773 gnd vdd FILL
XFILL_0_OAI21X1_751 gnd vdd FILL
XFILL_1_OAI21X1_955 gnd vdd FILL
XFILL_0_OAI21X1_795 gnd vdd FILL
XFILL_1_OAI21X1_977 gnd vdd FILL
XFILL_1_OR2X2_7 gnd vdd FILL
XFILL_1_OAI21X1_966 gnd vdd FILL
XFILL_1_OAI21X1_988 gnd vdd FILL
XFILL_1_OAI21X1_999 gnd vdd FILL
XBUFX2_809 BUFX2_809/A gnd tid1_o[25] vdd BUFX2
XFILL_28_7_1 gnd vdd FILL
XFILL_3_7_1 gnd vdd FILL
XFILL_27_2_0 gnd vdd FILL
XFILL_2_2_0 gnd vdd FILL
XFILL_0_OAI21X1_1561 gnd vdd FILL
XFILL_0_OAI21X1_1550 gnd vdd FILL
XFILL_0_OAI21X1_1594 gnd vdd FILL
XFILL_0_OAI21X1_1583 gnd vdd FILL
XFILL_0_OAI21X1_1572 gnd vdd FILL
XFILL_11_6_1 gnd vdd FILL
XFILL_10_1_0 gnd vdd FILL
XFILL_0_BUFX2_505 gnd vdd FILL
XFILL_0_BUFX2_516 gnd vdd FILL
XFILL_20_17_0 gnd vdd FILL
XFILL_0_BUFX2_538 gnd vdd FILL
XFILL_0_BUFX2_527 gnd vdd FILL
XCLKBUF1_8 BUFX4_87/Y gnd CLKBUF1_8/Y vdd CLKBUF1
XFILL_0_BUFX2_549 gnd vdd FILL
XBUFX4_102 BUFX4_7/A gnd BUFX4_102/Y vdd BUFX4
XBUFX4_146 BUFX4_17/Y gnd BUFX4_146/Y vdd BUFX4
XFILL_19_7_1 gnd vdd FILL
XBUFX4_113 INVX8_4/Y gnd BUFX4_378/A vdd BUFX4
XBUFX4_135 BUFX4_13/Y gnd BUFX4_135/Y vdd BUFX4
XFILL_0_INVX1_13 gnd vdd FILL
XFILL_0_INVX1_24 gnd vdd FILL
XBUFX4_124 BUFX4_16/Y gnd BUFX4_124/Y vdd BUFX4
XFILL_0_INVX1_68 gnd vdd FILL
XFILL_4_CLKBUF1_39 gnd vdd FILL
XBUFX4_168 BUFX4_19/Y gnd BUFX4_168/Y vdd BUFX4
XFILL_2_OAI21X1_1666 gnd vdd FILL
XBUFX4_179 BUFX4_18/Y gnd BUFX4_179/Y vdd BUFX4
XNOR2X1_206 bundleAddress_i[14] INVX1_213/Y gnd NOR2X1_206/Y vdd NOR2X1
XBUFX4_157 BUFX4_15/Y gnd BUFX4_157/Y vdd BUFX4
XFILL_18_2_0 gnd vdd FILL
XFILL_0_INVX1_46 gnd vdd FILL
XFILL_1_AND2X2_5 gnd vdd FILL
XFILL_0_INVX1_57 gnd vdd FILL
XFILL_2_OAI21X1_1644 gnd vdd FILL
XFILL_0_INVX1_35 gnd vdd FILL
XFILL_4_CLKBUF1_28 gnd vdd FILL
XFILL_2_OAI21X1_1699 gnd vdd FILL
XNOR2X1_217 INVX2_61/Y INVX1_219/Y gnd NOR2X1_217/Y vdd NOR2X1
XFILL_0_INVX1_79 gnd vdd FILL
XNOR2X1_228 INVX4_44/Y OR2X2_21/A gnd NOR2X1_228/Y vdd NOR2X1
XFILL_25_16_0 gnd vdd FILL
XOAI21X1_1003 BUFX4_303/Y INVX1_156/Y OAI21X1_1003/C gnd OAI21X1_1003/Y vdd OAI21X1
XFILL_1_OAI21X1_1212 gnd vdd FILL
XOAI21X1_1036 BUFX4_322/Y INVX2_54/Y NAND2X1_402/Y gnd OAI21X1_1036/Y vdd OAI21X1
XFILL_1_OAI21X1_1223 gnd vdd FILL
XDFFPOSX1_604 BUFX2_637/A CLKBUF1_50/Y OAI21X1_824/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1201 gnd vdd FILL
XOAI21X1_1014 BUFX4_157/Y BUFX4_32/Y BUFX2_371/A gnd OAI21X1_1015/C vdd OAI21X1
XOAI21X1_1025 BUFX4_303/Y INVX1_167/Y OAI21X1_1025/C gnd OAI21X1_1025/Y vdd OAI21X1
XOAI21X1_1047 BUFX4_386/Y INVX4_33/Y NAND2X1_413/Y gnd OAI21X1_1047/Y vdd OAI21X1
XFILL_1_DFFPOSX1_813 gnd vdd FILL
XFILL_1_OAI21X1_1256 gnd vdd FILL
XFILL_1_OAI21X1_1234 gnd vdd FILL
XFILL_1_DFFPOSX1_824 gnd vdd FILL
XOAI21X1_1069 BUFX4_381/Y INVX2_75/Y NAND2X1_435/Y gnd OAI21X1_1069/Y vdd OAI21X1
XFILL_1_OAI21X1_1245 gnd vdd FILL
XDFFPOSX1_615 BUFX2_260/A CLKBUF1_67/Y BUFX4_284/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_802 gnd vdd FILL
XDFFPOSX1_648 BUFX2_293/A CLKBUF1_4/Y OAI21X1_876/Y gnd vdd DFFPOSX1
XDFFPOSX1_626 INVX1_55/A CLKBUF1_54/Y OAI21X1_854/Y gnd vdd DFFPOSX1
XDFFPOSX1_637 INVX1_66/A CLKBUF1_10/Y OAI21X1_865/Y gnd vdd DFFPOSX1
XOAI21X1_1058 OAI21X1_4/A INVX2_70/Y NAND2X1_424/Y gnd OAI21X1_1058/Y vdd OAI21X1
XFILL_1_DFFPOSX1_835 gnd vdd FILL
XFILL_1_OAI21X1_1289 gnd vdd FILL
XFILL_1_OAI21X1_1278 gnd vdd FILL
XFILL_1_OAI21X1_207 gnd vdd FILL
XFILL_1_DFFPOSX1_857 gnd vdd FILL
XFILL_1_OAI21X1_1267 gnd vdd FILL
XDFFPOSX1_659 BUFX2_296/A CLKBUF1_54/Y OAI21X1_887/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_846 gnd vdd FILL
XFILL_1_OAI21X1_229 gnd vdd FILL
XFILL_1_DFFPOSX1_879 gnd vdd FILL
XFILL_1_OAI21X1_218 gnd vdd FILL
XNAND2X1_707 BUFX2_699/A BUFX4_209/Y gnd NAND2X1_707/Y vdd NAND2X1
XFILL_1_DFFPOSX1_868 gnd vdd FILL
XNAND2X1_718 BUFX2_800/A BUFX4_365/Y gnd NAND2X1_718/Y vdd NAND2X1
XNAND2X1_729 BUFX2_783/A BUFX4_341/Y gnd NAND2X1_729/Y vdd NAND2X1
XFILL_6_DFFPOSX1_494 gnd vdd FILL
XFILL_1_NAND2X1_213 gnd vdd FILL
XFILL_1_NAND2X1_202 gnd vdd FILL
XFILL_0_DFFPOSX1_414 gnd vdd FILL
XFILL_1_NAND2X1_235 gnd vdd FILL
XFILL_0_DFFPOSX1_403 gnd vdd FILL
XFILL_0_17_0 gnd vdd FILL
XFILL_1_NAND2X1_246 gnd vdd FILL
XFILL_1_NAND2X1_279 gnd vdd FILL
XFILL_1_NAND2X1_268 gnd vdd FILL
XFILL_0_DFFPOSX1_447 gnd vdd FILL
XFILL_0_DFFPOSX1_425 gnd vdd FILL
XFILL_0_DFFPOSX1_436 gnd vdd FILL
XFILL_0_DFFPOSX1_458 gnd vdd FILL
XFILL_0_DFFPOSX1_469 gnd vdd FILL
XFILL_5_DFFPOSX1_1030 gnd vdd FILL
XFILL_3_DFFPOSX1_918 gnd vdd FILL
XFILL_3_DFFPOSX1_929 gnd vdd FILL
XFILL_3_DFFPOSX1_907 gnd vdd FILL
XDFFPOSX1_30 BUFX2_700/A CLKBUF1_99/Y DFFPOSX1_30/D gnd vdd DFFPOSX1
XDFFPOSX1_52 BUFX2_721/A CLKBUF1_31/Y DFFPOSX1_52/D gnd vdd DFFPOSX1
XDFFPOSX1_63 BUFX2_733/A CLKBUF1_47/Y DFFPOSX1_63/D gnd vdd DFFPOSX1
XDFFPOSX1_41 BUFX2_740/A CLKBUF1_58/Y DFFPOSX1_41/D gnd vdd DFFPOSX1
XOAI21X1_1581 BUFX4_322/Y INVX2_117/Y NAND2X1_650/Y gnd OAI21X1_1581/Y vdd OAI21X1
XDFFPOSX1_85 BUFX2_754/A CLKBUF1_27/Y DFFPOSX1_85/D gnd vdd DFFPOSX1
XOAI21X1_1592 BUFX4_366/Y INVX2_128/Y NAND2X1_661/Y gnd OAI21X1_1592/Y vdd OAI21X1
XDFFPOSX1_96 BUFX2_766/A CLKBUF1_64/Y DFFPOSX1_96/D gnd vdd DFFPOSX1
XOAI21X1_1570 OR2X2_21/Y INVX4_49/Y INVX2_92/Y gnd NAND2X1_647/B vdd OAI21X1
XDFFPOSX1_74 BUFX2_773/A CLKBUF1_56/Y DFFPOSX1_74/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1790 gnd vdd FILL
XFILL_1_OAI21X1_730 gnd vdd FILL
XFILL_1_OAI21X1_763 gnd vdd FILL
XFILL_0_OAI21X1_570 gnd vdd FILL
XFILL_2_OAI21X1_923 gnd vdd FILL
XFILL_0_OAI21X1_581 gnd vdd FILL
XFILL_1_OAI21X1_741 gnd vdd FILL
XFILL_0_OAI21X1_592 gnd vdd FILL
XFILL_1_OAI21X1_752 gnd vdd FILL
XFILL_2_OAI21X1_912 gnd vdd FILL
XFILL_1_OAI21X1_796 gnd vdd FILL
XFILL_1_OAI21X1_785 gnd vdd FILL
XBUFX4_19 INVX8_6/Y gnd BUFX4_19/Y vdd BUFX4
XFILL_1_OAI21X1_774 gnd vdd FILL
XFILL_5_16_0 gnd vdd FILL
XBUFX2_628 BUFX2_628/A gnd majID4_o[15] vdd BUFX2
XFILL_2_DFFPOSX1_519 gnd vdd FILL
XBUFX2_606 BUFX2_606/A gnd majID4_o[35] vdd BUFX2
XBUFX2_617 INVX1_42/A gnd majID4_o[25] vdd BUFX2
XFILL_2_DFFPOSX1_508 gnd vdd FILL
XFILL_0_CLKBUF1_70 gnd vdd FILL
XBUFX2_639 BUFX2_639/A gnd majID4_o[5] vdd BUFX2
XFILL_0_CLKBUF1_81 gnd vdd FILL
XFILL_0_CLKBUF1_92 gnd vdd FILL
XFILL_0_OAI21X1_1391 gnd vdd FILL
XFILL_0_OAI21X1_1380 gnd vdd FILL
XFILL_0_DFFPOSX1_970 gnd vdd FILL
XFILL_0_DFFPOSX1_981 gnd vdd FILL
XFILL_0_DFFPOSX1_992 gnd vdd FILL
XINVX2_102 INVX2_102/A gnd INVX2_102/Y vdd INVX2
XFILL_0_BUFX2_313 gnd vdd FILL
XFILL_0_BUFX2_302 gnd vdd FILL
XINVX2_113 is64Bit_i gnd INVX2_113/Y vdd INVX2
XINVX2_124 bundlePid_i[24] gnd INVX2_124/Y vdd INVX2
XINVX2_146 bundleTid_i[63] gnd OAI21X1_8/A vdd INVX2
XFILL_0_BUFX2_335 gnd vdd FILL
XINVX2_135 bundlePid_i[13] gnd INVX2_135/Y vdd INVX2
XFILL_1_DFFPOSX1_109 gnd vdd FILL
XFILL_0_BUFX2_357 gnd vdd FILL
XFILL_0_BUFX2_346 gnd vdd FILL
XFILL_0_BUFX2_324 gnd vdd FILL
XFILL_0_BUFX2_379 gnd vdd FILL
XINVX2_157 bundleTid_i[52] gnd INVX2_157/Y vdd INVX2
XINVX2_179 bundleTid_i[30] gnd INVX2_179/Y vdd INVX2
XINVX2_168 bundleTid_i[41] gnd INVX2_168/Y vdd INVX2
XFILL_0_BUFX2_368 gnd vdd FILL
XFILL_14_13_1 gnd vdd FILL
XFILL_34_5_1 gnd vdd FILL
XFILL_2_OAI21X1_1485 gnd vdd FILL
XFILL_33_0_0 gnd vdd FILL
XFILL_22_2 gnd vdd FILL
XOAI21X1_509 INVX1_24/A INVX2_10/Y INVX2_11/Y gnd OAI21X1_510/C vdd OAI21X1
XFILL_1_NAND3X1_20 gnd vdd FILL
XFILL_1_OAI21X1_1031 gnd vdd FILL
XFILL_1_OAI21X1_1020 gnd vdd FILL
XFILL_1_NAND3X1_64 gnd vdd FILL
XFILL_1_NAND3X1_42 gnd vdd FILL
XDFFPOSX1_412 BUFX2_445/A CLKBUF1_1/Y OAI21X1_384/Y gnd vdd DFFPOSX1
XFILL_1_NAND3X1_31 gnd vdd FILL
XFILL_1_NAND3X1_53 gnd vdd FILL
XDFFPOSX1_401 BUFX2_433/A CLKBUF1_90/Y OAI21X1_373/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1053 gnd vdd FILL
XFILL_1_OAI21X1_1042 gnd vdd FILL
XFILL_1_DFFPOSX1_632 gnd vdd FILL
XFILL_1_OAI21X1_1064 gnd vdd FILL
XFILL_1_DFFPOSX1_621 gnd vdd FILL
XFILL_1_DFFPOSX1_610 gnd vdd FILL
XDFFPOSX1_456 BUFX2_487/A CLKBUF1_1/Y OAI21X1_454/Y gnd vdd DFFPOSX1
XDFFPOSX1_445 BUFX2_475/A CLKBUF1_50/Y OAI21X1_437/Y gnd vdd DFFPOSX1
XDFFPOSX1_423 BUFX2_480/A CLKBUF1_94/Y OAI21X1_399/Y gnd vdd DFFPOSX1
XDFFPOSX1_434 BUFX2_463/A CLKBUF1_13/Y OAI21X1_421/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_654 gnd vdd FILL
XFILL_0_BUFX2_880 gnd vdd FILL
XFILL_0_BUFX2_891 gnd vdd FILL
XDFFPOSX1_478 BUFX2_511/A CLKBUF1_5/Y OAI21X1_490/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1097 gnd vdd FILL
XDFFPOSX1_489 BUFX2_566/A CLKBUF1_94/Y OAI21X1_515/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_643 gnd vdd FILL
XFILL_1_DFFPOSX1_665 gnd vdd FILL
XFILL_1_OAI21X1_1075 gnd vdd FILL
XDFFPOSX1_467 BUFX2_499/A CLKBUF1_48/Y OAI21X1_471/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1086 gnd vdd FILL
XFILL_1_DFFPOSX1_698 gnd vdd FILL
XNAND2X1_515 BUFX2_82/A BUFX4_220/Y gnd NAND2X1_515/Y vdd NAND2X1
XINVX1_190 INVX1_190/A gnd INVX1_190/Y vdd INVX1
XNAND2X1_526 bundleAddress_i[35] XNOR2X1_65/A gnd XNOR2X1_66/A vdd NAND2X1
XFILL_19_12_1 gnd vdd FILL
XFILL_1_DFFPOSX1_687 gnd vdd FILL
XFILL_1_DFFPOSX1_676 gnd vdd FILL
XNAND2X1_504 BUFX2_76/A BUFX4_186/Y gnd NAND2X1_504/Y vdd NAND2X1
XNAND2X1_559 BUFX2_107/A BUFX4_203/Y gnd NAND2X1_559/Y vdd NAND2X1
XNAND2X1_537 BUFX2_95/A OAI21X1_9/B gnd NAND2X1_537/Y vdd NAND2X1
XNAND2X1_548 BUFX2_101/A BUFX4_226/Y gnd NAND2X1_548/Y vdd NAND2X1
XFILL_6_DFFPOSX1_280 gnd vdd FILL
XFILL_6_DFFPOSX1_291 gnd vdd FILL
XFILL_32_14_1 gnd vdd FILL
XFILL_0_AND2X2_16 gnd vdd FILL
XFILL_25_5_1 gnd vdd FILL
XFILL_0_AND2X2_27 gnd vdd FILL
XFILL_0_5_1 gnd vdd FILL
XFILL_0_DFFPOSX1_211 gnd vdd FILL
XFILL_0_DFFPOSX1_200 gnd vdd FILL
XFILL_24_0_0 gnd vdd FILL
XFILL_0_DFFPOSX1_222 gnd vdd FILL
XFILL_0_DFFPOSX1_255 gnd vdd FILL
XFILL_0_DFFPOSX1_266 gnd vdd FILL
XFILL_0_DFFPOSX1_244 gnd vdd FILL
XFILL_0_DFFPOSX1_233 gnd vdd FILL
XFILL_0_DFFPOSX1_299 gnd vdd FILL
XFILL_0_DFFPOSX1_277 gnd vdd FILL
XFILL_0_DFFPOSX1_288 gnd vdd FILL
XFILL_3_DFFPOSX1_704 gnd vdd FILL
XFILL_3_DFFPOSX1_715 gnd vdd FILL
XFILL_3_CLKBUF1_14 gnd vdd FILL
XFILL_3_DFFPOSX1_737 gnd vdd FILL
XFILL_3_DFFPOSX1_726 gnd vdd FILL
XFILL_3_CLKBUF1_25 gnd vdd FILL
XFILL_3_DFFPOSX1_759 gnd vdd FILL
XFILL_3_DFFPOSX1_748 gnd vdd FILL
XFILL_3_CLKBUF1_47 gnd vdd FILL
XFILL_3_CLKBUF1_36 gnd vdd FILL
XFILL_3_CLKBUF1_58 gnd vdd FILL
XFILL_3_CLKBUF1_69 gnd vdd FILL
XFILL_37_13_1 gnd vdd FILL
XFILL_1_NOR2X1_121 gnd vdd FILL
XFILL_1_NOR2X1_110 gnd vdd FILL
XDFFPOSX1_990 BUFX2_243/A CLKBUF1_20/Y OAI21X1_1549/Y gnd vdd DFFPOSX1
XFILL_8_6_1 gnd vdd FILL
XFILL_1_OAI21X1_571 gnd vdd FILL
XFILL_2_OAI21X1_720 gnd vdd FILL
XFILL_1_NOR2X1_154 gnd vdd FILL
XFILL_1_OAI21X1_560 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XFILL_1_OAI21X1_582 gnd vdd FILL
XFILL_1_NOR2X1_187 gnd vdd FILL
XFILL_1_NOR2X1_198 gnd vdd FILL
XFILL_1_OAI21X1_593 gnd vdd FILL
XBUFX2_403 BUFX2_403/A gnd majID1_o[45] vdd BUFX2
XFILL_2_DFFPOSX1_316 gnd vdd FILL
XBUFX2_425 BUFX2_425/A gnd majID1_o[25] vdd BUFX2
XFILL_2_DFFPOSX1_327 gnd vdd FILL
XFILL_2_DFFPOSX1_338 gnd vdd FILL
XBUFX2_414 BUFX2_414/A gnd majID1_o[35] vdd BUFX2
XBUFX2_436 BUFX2_436/A gnd majID1_o[15] vdd BUFX2
XFILL_2_DFFPOSX1_305 gnd vdd FILL
XBUFX2_447 BUFX2_447/A gnd majID1_o[5] vdd BUFX2
XFILL_2_DFFPOSX1_349 gnd vdd FILL
XFILL_16_5_1 gnd vdd FILL
XBUFX2_469 BUFX2_469/A gnd majID2_o[61] vdd BUFX2
XBUFX2_458 INVX1_6/A gnd majID2_o[62] vdd BUFX2
XFILL_15_0_0 gnd vdd FILL
XFILL_5_DFFPOSX1_809 gnd vdd FILL
XFILL_1_BUFX4_330 gnd vdd FILL
XFILL_1_BUFX4_363 gnd vdd FILL
XFILL_1_BUFX4_352 gnd vdd FILL
XFILL_1_BUFX4_341 gnd vdd FILL
XFILL_1_BUFX4_374 gnd vdd FILL
XFILL_1_BUFX4_385 gnd vdd FILL
XFILL_2_OAI21X1_32 gnd vdd FILL
XFILL_0_BUFX2_110 gnd vdd FILL
XFILL_0_BUFX2_121 gnd vdd FILL
XFILL_2_OAI21X1_54 gnd vdd FILL
XFILL_0_BUFX2_132 gnd vdd FILL
XFILL_0_BUFX2_154 gnd vdd FILL
XFILL_0_BUFX2_143 gnd vdd FILL
XFILL_0_BUFX2_165 gnd vdd FILL
XFILL_0_BUFX2_198 gnd vdd FILL
XFILL_0_BUFX2_187 gnd vdd FILL
XFILL_0_BUFX2_176 gnd vdd FILL
XFILL_1_DFFPOSX1_8 gnd vdd FILL
XFILL_2_OAI21X1_1260 gnd vdd FILL
XFILL_2_OAI21X1_1282 gnd vdd FILL
XFILL_2_DFFPOSX1_850 gnd vdd FILL
XFILL_2_OAI21X1_1271 gnd vdd FILL
XFILL_2_DFFPOSX1_883 gnd vdd FILL
XFILL_2_DFFPOSX1_872 gnd vdd FILL
XFILL_2_OAI21X1_1293 gnd vdd FILL
XBUFX2_970 BUFX2_970/A gnd tid4_o[62] vdd BUFX2
XBUFX2_992 BUFX2_992/A gnd tid4_o[60] vdd BUFX2
XBUFX2_981 BUFX2_981/A gnd tid4_o[61] vdd BUFX2
XFILL_2_DFFPOSX1_861 gnd vdd FILL
XFILL_2_DFFPOSX1_894 gnd vdd FILL
XOAI21X1_306 BUFX4_178/Y BUFX4_50/Y BUFX2_1018/A gnd OAI21X1_307/C vdd OAI21X1
XOAI21X1_328 INVX4_1/Y BUFX4_321/Y NAND2X1_72/Y gnd OAI21X1_328/Y vdd OAI21X1
XOAI21X1_317 INVX2_2/Y BUFX4_299/Y OAI21X1_317/C gnd OAI21X1_317/Y vdd OAI21X1
XOAI21X1_339 BUFX4_387/Y INVX4_4/Y NAND2X1_83/Y gnd OAI21X1_339/Y vdd OAI21X1
XDFFPOSX1_220 BUFX2_893/A CLKBUF1_93/Y OAI21X1_64/Y gnd vdd DFFPOSX1
XDFFPOSX1_231 BUFX2_928/A CLKBUF1_45/Y OAI21X1_79/Y gnd vdd DFFPOSX1
XBUFX4_4 BUFX4_4/A gnd BUFX4_4/Y vdd BUFX4
XDFFPOSX1_242 BUFX2_911/A CLKBUF1_25/Y OAI21X1_101/Y gnd vdd DFFPOSX1
XDFFPOSX1_253 BUFX2_923/A CLKBUF1_35/Y OAI21X1_123/Y gnd vdd DFFPOSX1
XDFFPOSX1_264 BUFX2_935/A CLKBUF1_35/Y OAI21X1_145/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_440 gnd vdd FILL
XDFFPOSX1_275 BUFX2_947/A CLKBUF1_16/Y OAI21X1_167/Y gnd vdd DFFPOSX1
XNAND2X1_301 NOR2X1_96/B OAI21X1_639/A gnd OAI21X1_637/A vdd NAND2X1
XFILL_1_DFFPOSX1_484 gnd vdd FILL
XFILL_1_DFFPOSX1_462 gnd vdd FILL
XFILL_1_DFFPOSX1_451 gnd vdd FILL
XFILL_1_DFFPOSX1_473 gnd vdd FILL
XDFFPOSX1_297 BUFX2_1014/A CLKBUF1_81/Y OAI21X1_211/Y gnd vdd DFFPOSX1
XDFFPOSX1_286 BUFX2_959/A CLKBUF1_2/Y OAI21X1_189/Y gnd vdd DFFPOSX1
XNAND2X1_334 BUFX4_288/Y NOR3X1_11/C gnd OAI21X1_832/B vdd NAND2X1
XNAND2X1_345 BUFX4_261/Y bundle_i[24] gnd OAI21X1_851/C vdd NAND2X1
XFILL_3_NOR3X1_17 gnd vdd FILL
XNAND2X1_323 XNOR2X1_47/A OAI21X1_739/Y gnd OAI21X1_741/A vdd NAND2X1
XFILL_1_DFFPOSX1_495 gnd vdd FILL
XNAND2X1_312 NAND2X1_312/A INVX1_35/A gnd OAI21X1_683/A vdd NAND2X1
XNAND2X1_367 BUFX4_263/Y bundle_i[2] gnd OAI21X1_873/C vdd NAND2X1
XNAND2X1_378 BUFX2_323/A BUFX4_208/Y gnd OAI21X1_884/C vdd NAND2X1
XNAND2X1_356 INVX8_4/A bundle_i[13] gnd OAI21X1_862/C vdd NAND2X1
XFILL_4_DFFPOSX1_900 gnd vdd FILL
XFILL_4_DFFPOSX1_922 gnd vdd FILL
XFILL_4_DFFPOSX1_911 gnd vdd FILL
XFILL_4_DFFPOSX1_944 gnd vdd FILL
XFILL_4_DFFPOSX1_955 gnd vdd FILL
XFILL_4_DFFPOSX1_933 gnd vdd FILL
XNAND2X1_389 BUFX2_304/A BUFX4_228/Y gnd OAI21X1_895/C vdd NAND2X1
XFILL_4_DFFPOSX1_966 gnd vdd FILL
XFILL_4_DFFPOSX1_999 gnd vdd FILL
XFILL_4_DFFPOSX1_977 gnd vdd FILL
XFILL_4_DFFPOSX1_988 gnd vdd FILL
XFILL_1_BUFX2_801 gnd vdd FILL
XFILL_1_BUFX2_812 gnd vdd FILL
XFILL_1_BUFX2_845 gnd vdd FILL
XFILL_1_BUFX2_834 gnd vdd FILL
XINVX4_4 bundleStartMajId_i[52] gnd INVX4_4/Y vdd INVX4
XFILL_1_BUFX2_856 gnd vdd FILL
XOAI21X1_840 AOI21X1_35/Y OAI21X1_840/B OAI21X1_840/C gnd OAI21X1_840/Y vdd OAI21X1
XFILL_3_DFFPOSX1_512 gnd vdd FILL
XFILL_2_NOR3X1_9 gnd vdd FILL
XFILL_3_DFFPOSX1_501 gnd vdd FILL
XFILL_1_BUFX2_889 gnd vdd FILL
XOAI21X1_851 INVX1_52/Y BUFX4_261/Y OAI21X1_851/C gnd OAI21X1_851/Y vdd OAI21X1
XOAI21X1_873 INVX1_74/Y BUFX4_263/Y OAI21X1_873/C gnd OAI21X1_873/Y vdd OAI21X1
XOAI21X1_884 INVX1_85/Y BUFX4_208/Y OAI21X1_884/C gnd OAI21X1_884/Y vdd OAI21X1
XOAI21X1_862 INVX1_63/Y BUFX4_267/Y OAI21X1_862/C gnd OAI21X1_862/Y vdd OAI21X1
XFILL_3_DFFPOSX1_545 gnd vdd FILL
XFILL_3_DFFPOSX1_534 gnd vdd FILL
XFILL_3_DFFPOSX1_523 gnd vdd FILL
XFILL_3_DFFPOSX1_556 gnd vdd FILL
XFILL_3_DFFPOSX1_578 gnd vdd FILL
XFILL_3_DFFPOSX1_567 gnd vdd FILL
XFILL_3_DFFPOSX1_589 gnd vdd FILL
XOAI21X1_895 INVX1_96/Y BUFX4_228/Y OAI21X1_895/C gnd OAI21X1_895/Y vdd OAI21X1
XFILL_2_OAI21X1_583 gnd vdd FILL
XFILL_1_OAI21X1_390 gnd vdd FILL
XBUFX2_211 BUFX2_211/A gnd addr4_o[38] vdd BUFX2
XBUFX2_200 BUFX2_200/A gnd addr4_o[48] vdd BUFX2
XFILL_0_NAND2X1_608 gnd vdd FILL
XFILL_2_DFFPOSX1_102 gnd vdd FILL
XFILL_2_DFFPOSX1_113 gnd vdd FILL
XFILL_2_DFFPOSX1_124 gnd vdd FILL
XBUFX2_233 BUFX2_233/A gnd addr4_o[18] vdd BUFX2
XFILL_2_DFFPOSX1_135 gnd vdd FILL
XFILL_0_NAND2X1_619 gnd vdd FILL
XFILL_0_NAND3X1_50 gnd vdd FILL
XFILL_0_NAND3X1_61 gnd vdd FILL
XFILL_2_DFFPOSX1_146 gnd vdd FILL
XBUFX2_222 BUFX2_222/A gnd addr4_o[28] vdd BUFX2
XBUFX2_244 BUFX2_244/A gnd addr4_o[8] vdd BUFX2
XFILL_2_DFFPOSX1_157 gnd vdd FILL
XFILL_2_DFFPOSX1_179 gnd vdd FILL
XBUFX2_277 INVX1_68/A gnd instr1_o[8] vdd BUFX2
XFILL_2_DFFPOSX1_168 gnd vdd FILL
XBUFX2_255 BUFX2_255/A gnd addr4_o[55] vdd BUFX2
XBUFX2_266 INVX1_58/A gnd instr1_o[18] vdd BUFX2
XBUFX2_299 BUFX2_299/A gnd instr2_o[17] vdd BUFX2
XBUFX2_288 INVX1_50/A gnd instr1_o[26] vdd BUFX2
XFILL_31_3_1 gnd vdd FILL
XFILL_28_18_1 gnd vdd FILL
XFILL_5_DFFPOSX1_606 gnd vdd FILL
XFILL_5_DFFPOSX1_617 gnd vdd FILL
XFILL_5_DFFPOSX1_628 gnd vdd FILL
XFILL_5_DFFPOSX1_639 gnd vdd FILL
XFILL_1_BUFX4_171 gnd vdd FILL
XFILL_1_BUFX4_160 gnd vdd FILL
XFILL_1_BUFX4_182 gnd vdd FILL
XFILL_1_BUFX4_193 gnd vdd FILL
XFILL_22_14_0 gnd vdd FILL
XFILL_4_DFFPOSX1_218 gnd vdd FILL
XFILL_4_DFFPOSX1_207 gnd vdd FILL
XNAND3X1_7 AND2X2_7/Y NOR2X1_11/Y NOR2X1_30/Y gnd NOR3X1_2/C vdd NAND3X1
XFILL_4_DFFPOSX1_229 gnd vdd FILL
XFILL_2_CLKBUF1_11 gnd vdd FILL
XFILL_2_CLKBUF1_22 gnd vdd FILL
XFILL_2_BUFX4_317 gnd vdd FILL
XFILL_2_CLKBUF1_55 gnd vdd FILL
XFILL_2_CLKBUF1_44 gnd vdd FILL
XFILL_2_CLKBUF1_33 gnd vdd FILL
XFILL_2_CLKBUF1_66 gnd vdd FILL
XFILL_2_CLKBUF1_99 gnd vdd FILL
XFILL_2_CLKBUF1_88 gnd vdd FILL
XFILL_2_CLKBUF1_77 gnd vdd FILL
XFILL_2_DFFPOSX1_691 gnd vdd FILL
XFILL_2_DFFPOSX1_680 gnd vdd FILL
XFILL_22_3_1 gnd vdd FILL
XFILL_0_NOR2X1_140 gnd vdd FILL
XOAI21X1_103 BUFX4_132/Y INVX2_161/Y OAI21X1_103/C gnd OAI21X1_103/Y vdd OAI21X1
XFILL_27_13_0 gnd vdd FILL
XFILL_0_NOR2X1_151 gnd vdd FILL
XFILL_0_NOR2X1_162 gnd vdd FILL
XFILL_1_BUFX2_119 gnd vdd FILL
XFILL_0_NOR2X1_173 gnd vdd FILL
XOAI21X1_125 BUFX4_148/Y INVX2_172/Y OAI21X1_125/C gnd OAI21X1_125/Y vdd OAI21X1
XOAI21X1_114 BUFX4_8/Y BUFX4_368/Y BUFX2_919/A gnd OAI21X1_115/C vdd OAI21X1
XFILL_0_NOR2X1_184 gnd vdd FILL
XOAI21X1_147 BUFX4_150/Y INVX2_183/Y OAI21X1_147/C gnd OAI21X1_147/Y vdd OAI21X1
XFILL_0_NOR2X1_195 gnd vdd FILL
XFILL_0_DFFPOSX1_1003 gnd vdd FILL
XOAI21X1_136 BUFX4_102/Y OAI21X1_6/A BUFX2_931/A gnd OAI21X1_137/C vdd OAI21X1
XOAI21X1_158 BUFX4_11/A BUFX4_380/Y BUFX2_943/A gnd OAI21X1_159/C vdd OAI21X1
XFILL_0_DFFPOSX1_1014 gnd vdd FILL
XOAI21X1_169 BUFX4_148/Y INVX2_194/Y OAI21X1_169/C gnd OAI21X1_169/Y vdd OAI21X1
XFILL_0_DFFPOSX1_1025 gnd vdd FILL
XBUFX2_1 BUFX2_1/A gnd addr1_o[63] vdd BUFX2
XFILL_1_DFFPOSX1_281 gnd vdd FILL
XFILL_1_DFFPOSX1_292 gnd vdd FILL
XFILL_1_DFFPOSX1_270 gnd vdd FILL
XNAND2X1_131 BUFX2_448/A BUFX4_316/Y gnd OAI21X1_387/C vdd NAND2X1
XNAND2X1_142 BUFX2_480/A BUFX4_222/Y gnd OAI21X1_399/C vdd NAND2X1
XNAND2X1_120 BUFX2_436/A BUFX4_345/Y gnd OAI21X1_376/C vdd NAND2X1
XNAND2X1_153 BUFX2_519/A BUFX4_181/Y gnd OAI21X1_411/C vdd NAND2X1
XFILL_8_18_1 gnd vdd FILL
XFILL_0_XNOR2X1_18 gnd vdd FILL
XNAND2X1_175 OAI21X1_428/Y NAND2X1_177/B gnd OAI21X1_429/A vdd NAND2X1
XNAND2X1_186 AND2X2_4/Y AND2X2_5/Y gnd NOR2X1_16/A vdd NAND2X1
XNAND2X1_164 BUFX2_464/A BUFX4_215/Y gnd OAI21X1_422/C vdd NAND2X1
XFILL_5_4_1 gnd vdd FILL
XFILL_4_DFFPOSX1_730 gnd vdd FILL
XFILL_4_DFFPOSX1_741 gnd vdd FILL
XFILL_4_DFFPOSX1_752 gnd vdd FILL
XFILL_4_DFFPOSX1_774 gnd vdd FILL
XFILL_1_OAI21X1_51 gnd vdd FILL
XFILL_4_DFFPOSX1_763 gnd vdd FILL
XFILL_1_OAI21X1_40 gnd vdd FILL
XFILL_0_XNOR2X1_29 gnd vdd FILL
XNAND2X1_197 BUFX2_478/A BUFX4_214/Y gnd OAI21X1_443/C vdd NAND2X1
XFILL_1_OAI21X1_62 gnd vdd FILL
XFILL_1_OAI21X1_84 gnd vdd FILL
XFILL_1_OAI21X1_95 gnd vdd FILL
XFILL_1_OAI21X1_73 gnd vdd FILL
XFILL_2_14_0 gnd vdd FILL
XFILL_4_DFFPOSX1_785 gnd vdd FILL
XFILL_4_DFFPOSX1_796 gnd vdd FILL
XFILL_0_DFFPOSX1_5 gnd vdd FILL
XFILL_13_3_1 gnd vdd FILL
XINVX2_1 bundleTid_i[6] gnd INVX2_1/Y vdd INVX2
XFILL_0_BUFX4_205 gnd vdd FILL
XFILL_1_BUFX2_653 gnd vdd FILL
XFILL_1_BUFX2_642 gnd vdd FILL
XFILL_1_BUFX2_697 gnd vdd FILL
XFILL_0_BUFX4_216 gnd vdd FILL
XFILL_0_BUFX4_227 gnd vdd FILL
XFILL_0_BUFX4_249 gnd vdd FILL
XFILL_3_DFFPOSX1_331 gnd vdd FILL
XFILL_0_BUFX4_238 gnd vdd FILL
XAOI21X1_1 INVX2_42/Y NOR2X1_17/Y bundleStartMajId_i[36] gnd AOI21X1_1/Y vdd AOI21X1
XFILL_1_BUFX2_686 gnd vdd FILL
XFILL_3_DFFPOSX1_320 gnd vdd FILL
XFILL_3_DFFPOSX1_342 gnd vdd FILL
XFILL_1_OAI21X1_1608 gnd vdd FILL
XFILL_3_DFFPOSX1_353 gnd vdd FILL
XOAI21X1_681 OAI21X1_681/A BUFX4_290/Y OAI21X1_681/C gnd OAI21X1_681/Y vdd OAI21X1
XOAI21X1_692 OAI21X1_692/A BUFX4_302/Y OAI21X1_692/C gnd OAI21X1_692/Y vdd OAI21X1
XOAI21X1_670 BUFX4_135/Y BUFX4_49/Y BUFX2_619/A gnd OAI21X1_671/C vdd OAI21X1
XFILL_3_DFFPOSX1_364 gnd vdd FILL
XFILL_1_OAI21X1_1619 gnd vdd FILL
XFILL_3_DFFPOSX1_375 gnd vdd FILL
XFILL_3_DFFPOSX1_397 gnd vdd FILL
XFILL_3_DFFPOSX1_386 gnd vdd FILL
XFILL_6_DFFPOSX1_802 gnd vdd FILL
XFILL_6_DFFPOSX1_813 gnd vdd FILL
XFILL_6_DFFPOSX1_835 gnd vdd FILL
XFILL_6_DFFPOSX1_824 gnd vdd FILL
XFILL_0_INVX4_24 gnd vdd FILL
XFILL_0_INVX4_13 gnd vdd FILL
XFILL_0_INVX4_35 gnd vdd FILL
XFILL_3_DFFPOSX1_1018 gnd vdd FILL
XFILL_3_DFFPOSX1_1007 gnd vdd FILL
XFILL_0_INVX4_46 gnd vdd FILL
XFILL_3_DFFPOSX1_1029 gnd vdd FILL
XXNOR2X1_31 XNOR2X1_31/A INVX4_10/Y gnd XNOR2X1_31/Y vdd XNOR2X1
XXNOR2X1_20 NOR3X1_2/Y bundleStartMajId_i[18] gnd XNOR2X1_20/Y vdd XNOR2X1
XXNOR2X1_64 XNOR2X1_64/A bundleAddress_i[36] gnd XNOR2X1_64/Y vdd XNOR2X1
XXNOR2X1_75 XNOR2X1_75/A bundleAddress_i[53] gnd XNOR2X1_75/Y vdd XNOR2X1
XXNOR2X1_53 INVX2_53/A bundleStartMajId_i[14] gnd XNOR2X1_53/Y vdd XNOR2X1
XXNOR2X1_42 AND2X2_20/A bundleStartMajId_i[50] gnd XNOR2X1_42/Y vdd XNOR2X1
XFILL_7_13_0 gnd vdd FILL
XFILL_1_INVX2_171 gnd vdd FILL
XXNOR2X1_97 XNOR2X1_97/A INVX4_37/Y gnd XNOR2X1_97/Y vdd XNOR2X1
XXNOR2X1_86 NOR3X1_18/Y bundleAddress_i[12] gnd XNOR2X1_86/Y vdd XNOR2X1
XFILL_0_NAND2X1_405 gnd vdd FILL
XFILL_0_NAND2X1_416 gnd vdd FILL
XFILL_1_XNOR2X1_9 gnd vdd FILL
XBUFX2_63 BUFX2_63/A gnd addr1_o[55] vdd BUFX2
XFILL_0_OAI21X1_1209 gnd vdd FILL
XFILL_0_NAND2X1_449 gnd vdd FILL
XBUFX2_41 BUFX2_41/A gnd addr1_o[18] vdd BUFX2
XFILL_0_NAND2X1_427 gnd vdd FILL
XFILL_11_11_1 gnd vdd FILL
XBUFX2_52 BUFX2_52/A gnd addr1_o[8] vdd BUFX2
XFILL_1_NAND2X1_609 gnd vdd FILL
XBUFX2_30 BUFX2_30/A gnd addr1_o[28] vdd BUFX2
XFILL_0_NAND2X1_438 gnd vdd FILL
XBUFX2_85 BUFX2_85/A gnd addr2_o[36] vdd BUFX2
XBUFX2_74 BUFX2_74/A gnd addr2_o[46] vdd BUFX2
XBUFX2_96 BUFX2_96/A gnd addr2_o[26] vdd BUFX2
XFILL_5_DFFPOSX1_403 gnd vdd FILL
XFILL_5_DFFPOSX1_414 gnd vdd FILL
XFILL_5_DFFPOSX1_425 gnd vdd FILL
XFILL_5_DFFPOSX1_436 gnd vdd FILL
XFILL_5_DFFPOSX1_458 gnd vdd FILL
XFILL_5_DFFPOSX1_469 gnd vdd FILL
XFILL_5_DFFPOSX1_447 gnd vdd FILL
XFILL_1_BUFX4_63 gnd vdd FILL
XFILL_1_BUFX4_52 gnd vdd FILL
XFILL_1_BUFX4_41 gnd vdd FILL
XFILL_1_BUFX4_30 gnd vdd FILL
XFILL_1_BUFX4_85 gnd vdd FILL
XFILL_1_BUFX4_96 gnd vdd FILL
XFILL_1_BUFX4_74 gnd vdd FILL
XFILL_0_AOI21X1_18 gnd vdd FILL
XFILL_0_AOI21X1_29 gnd vdd FILL
XFILL_0_OAI21X1_900 gnd vdd FILL
XFILL_0_OAI21X1_933 gnd vdd FILL
XFILL_0_OAI21X1_911 gnd vdd FILL
XFILL_0_OAI21X1_922 gnd vdd FILL
XFILL_2_CLKBUF1_9 gnd vdd FILL
XFILL_0_OAI21X1_944 gnd vdd FILL
XFILL_0_OAI21X1_955 gnd vdd FILL
XFILL_0_OAI21X1_966 gnd vdd FILL
XFILL_0_OAI21X1_999 gnd vdd FILL
XFILL_0_OAI21X1_977 gnd vdd FILL
XFILL_0_OAI21X1_988 gnd vdd FILL
XFILL_16_10_1 gnd vdd FILL
XFILL_0_OAI21X1_1710 gnd vdd FILL
XFILL_1_OR2X2_11 gnd vdd FILL
XFILL_0_OAI21X1_1743 gnd vdd FILL
XFILL_0_OAI21X1_1732 gnd vdd FILL
XFILL_0_OAI21X1_1721 gnd vdd FILL
XFILL_0_OAI21X1_1754 gnd vdd FILL
XFILL_0_OAI21X1_1765 gnd vdd FILL
XFILL_0_OAI21X1_1776 gnd vdd FILL
XFILL_0_OAI21X1_1798 gnd vdd FILL
XFILL_0_OAI21X1_1787 gnd vdd FILL
XFILL_5_DFFPOSX1_981 gnd vdd FILL
XFILL_5_DFFPOSX1_970 gnd vdd FILL
XFILL_5_DFFPOSX1_992 gnd vdd FILL
XAOI21X1_53 bundleAddress_i[16] INVX1_212/Y bundleAddress_i[15] gnd AOI21X1_53/Y vdd
+ AOI21X1
XFILL_0_NOR2X1_38 gnd vdd FILL
XAOI21X1_20 bundleStartMajId_i[10] NOR2X1_95/Y bundleStartMajId_i[9] gnd AOI21X1_20/Y
+ vdd AOI21X1
XAOI21X1_31 bundleStartMajId_i[46] INVX1_36/Y bundleStartMajId_i[45] gnd AOI21X1_31/Y
+ vdd AOI21X1
XFILL_0_NOR2X1_27 gnd vdd FILL
XFILL_0_NOR2X1_16 gnd vdd FILL
XFILL_0_BUFX2_709 gnd vdd FILL
XAOI21X1_42 bundleAddress_i[8] NOR3X1_14/Y bundleAddress_i[7] gnd AOI21X1_42/Y vdd
+ AOI21X1
XFILL_0_NOR2X1_49 gnd vdd FILL
XAOI21X1_64 bundleAddress_i[8] INVX1_226/Y bundleAddress_i[7] gnd AOI21X1_64/Y vdd
+ AOI21X1
XOAI21X1_4 OAI21X1_4/A INVX2_4/Y OAI21X1_4/C gnd OAI21X1_4/Y vdd OAI21X1
XFILL_6_DFFPOSX1_109 gnd vdd FILL
XFILL_18_18_0 gnd vdd FILL
XFILL_34_11_1 gnd vdd FILL
XXNOR2X1_101 NAND3X1_65/Y INVX8_3/Y gnd XNOR2X1_101/Y vdd XNOR2X1
XFILL_2_OAI21X1_1804 gnd vdd FILL
XBUFX4_328 BUFX4_386/A gnd BUFX4_328/Y vdd BUFX4
XBUFX4_317 BUFX4_378/A gnd BUFX4_317/Y vdd BUFX4
XBUFX4_306 BUFX4_310/A gnd NOR2X1_96/B vdd BUFX4
XBUFX4_339 BUFX4_381/A gnd BUFX4_339/Y vdd BUFX4
XFILL_4_DFFPOSX1_582 gnd vdd FILL
XFILL_4_DFFPOSX1_560 gnd vdd FILL
XFILL_4_DFFPOSX1_571 gnd vdd FILL
XFILL_4_DFFPOSX1_593 gnd vdd FILL
XFILL_1_BUFX2_450 gnd vdd FILL
XFILL_1_BUFX2_461 gnd vdd FILL
XOAI21X1_1229 INVX4_47/Y NOR2X1_180/A OAI21X1_1229/C gnd OAI21X1_1231/A vdd OAI21X1
XOAI21X1_1218 INVX2_58/Y INVX1_183/A BUFX4_305/Y gnd OAI21X1_1220/A vdd OAI21X1
XFILL_1_OAI21X1_1405 gnd vdd FILL
XFILL_1_CLKBUF1_30 gnd vdd FILL
XOAI21X1_1207 AND2X2_25/Y OAI21X1_1207/B NAND2X1_589/Y gnd OAI21X1_1207/Y vdd OAI21X1
XFILL_1_BUFX2_494 gnd vdd FILL
XFILL_1_BUFX2_483 gnd vdd FILL
XDFFPOSX1_808 BUFX2_65/A CLKBUF1_17/Y OAI21X1_1100/Y gnd vdd DFFPOSX1
XFILL_3_DFFPOSX1_150 gnd vdd FILL
XFILL_1_CLKBUF1_74 gnd vdd FILL
XDFFPOSX1_819 BUFX2_68/A CLKBUF1_5/Y OAI21X1_1122/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1427 gnd vdd FILL
XFILL_1_OAI21X1_1416 gnd vdd FILL
XFILL_1_OAI21X1_1438 gnd vdd FILL
XFILL_1_CLKBUF1_63 gnd vdd FILL
XFILL_3_DFFPOSX1_161 gnd vdd FILL
XFILL_1_CLKBUF1_41 gnd vdd FILL
XFILL_3_DFFPOSX1_172 gnd vdd FILL
XFILL_1_INVX8_3 gnd vdd FILL
XFILL_1_CLKBUF1_52 gnd vdd FILL
XFILL_3_DFFPOSX1_194 gnd vdd FILL
XFILL_1_CLKBUF1_96 gnd vdd FILL
XFILL_3_DFFPOSX1_183 gnd vdd FILL
XFILL_0_OAI21X1_218 gnd vdd FILL
XFILL_1_CLKBUF1_85 gnd vdd FILL
XFILL_0_OAI21X1_207 gnd vdd FILL
XFILL_1_OAI21X1_1449 gnd vdd FILL
XFILL_0_OAI21X1_229 gnd vdd FILL
XFILL_3_1 gnd vdd FILL
XFILL_6_DFFPOSX1_687 gnd vdd FILL
XFILL_6_DFFPOSX1_676 gnd vdd FILL
XFILL_6_DFFPOSX1_698 gnd vdd FILL
XFILL_36_2_1 gnd vdd FILL
XFILL_1_NAND2X1_406 gnd vdd FILL
XFILL_0_NAND2X1_213 gnd vdd FILL
XFILL_0_NAND2X1_224 gnd vdd FILL
XFILL_0_NAND2X1_202 gnd vdd FILL
XFILL_0_OAI21X1_1028 gnd vdd FILL
XFILL_0_OAI21X1_1039 gnd vdd FILL
XFILL_1_NAND2X1_417 gnd vdd FILL
XFILL_0_OAI21X1_1006 gnd vdd FILL
XFILL_0_NAND2X1_257 gnd vdd FILL
XFILL_0_NAND2X1_235 gnd vdd FILL
XFILL_1_NAND2X1_428 gnd vdd FILL
XFILL_0_OAI21X1_1017 gnd vdd FILL
XFILL_0_NAND2X1_268 gnd vdd FILL
XFILL_0_NAND2X1_246 gnd vdd FILL
XFILL_1_NAND2X1_439 gnd vdd FILL
XFILL_0_DFFPOSX1_607 gnd vdd FILL
XFILL_0_NAND2X1_279 gnd vdd FILL
XFILL_0_DFFPOSX1_629 gnd vdd FILL
XFILL_0_DFFPOSX1_618 gnd vdd FILL
XFILL_5_DFFPOSX1_211 gnd vdd FILL
XFILL_5_DFFPOSX1_200 gnd vdd FILL
XFILL_5_DFFPOSX1_244 gnd vdd FILL
XFILL_5_DFFPOSX1_222 gnd vdd FILL
XFILL_5_DFFPOSX1_233 gnd vdd FILL
XFILL_5_DFFPOSX1_255 gnd vdd FILL
XFILL_5_DFFPOSX1_266 gnd vdd FILL
XFILL_5_DFFPOSX1_277 gnd vdd FILL
XFILL_5_DFFPOSX1_299 gnd vdd FILL
XFILL_5_DFFPOSX1_288 gnd vdd FILL
XFILL_0_OAI21X1_81 gnd vdd FILL
XOAI21X1_1730 BUFX4_137/Y BUFX4_53/Y BUFX2_747/A gnd OAI21X1_1731/C vdd OAI21X1
XOAI21X1_1741 INVX2_132/Y BUFX4_301/Y OAI21X1_1741/C gnd DFFPOSX1_83/D vdd OAI21X1
XFILL_0_OAI21X1_92 gnd vdd FILL
XFILL_0_OAI21X1_70 gnd vdd FILL
XOAI21X1_1763 INVX2_143/Y BUFX4_293/Y OAI21X1_1763/C gnd DFFPOSX1_94/D vdd OAI21X1
XOAI21X1_1752 BUFX4_151/Y BUFX4_70/Y BUFX2_759/A gnd OAI21X1_1753/C vdd OAI21X1
XOAI21X1_1774 BUFX4_334/Y OAI21X1_8/A NAND2X1_715/Y gnd OAI21X1_1774/Y vdd OAI21X1
XOAI21X1_1785 BUFX4_363/Y INVX2_157/Y NAND2X1_726/Y gnd OAI21X1_1785/Y vdd OAI21X1
XOAI21X1_1796 BUFX4_375/Y INVX2_168/Y NAND2X1_737/Y gnd OAI21X1_1796/Y vdd OAI21X1
XFILL_0_OAI21X1_741 gnd vdd FILL
XFILL_0_OAI21X1_730 gnd vdd FILL
XFILL_1_OAI21X1_901 gnd vdd FILL
XFILL_1_OAI21X1_912 gnd vdd FILL
XFILL_1_OAI21X1_945 gnd vdd FILL
XFILL_0_OAI21X1_763 gnd vdd FILL
XFILL_1_OAI21X1_923 gnd vdd FILL
XFILL_0_OAI21X1_774 gnd vdd FILL
XFILL_0_OAI21X1_752 gnd vdd FILL
XFILL_1_OAI21X1_934 gnd vdd FILL
XFILL_1_OAI21X1_978 gnd vdd FILL
XFILL_1_OAI21X1_956 gnd vdd FILL
XFILL_0_OAI21X1_796 gnd vdd FILL
XFILL_0_OAI21X1_785 gnd vdd FILL
XFILL_1_OR2X2_8 gnd vdd FILL
XFILL_1_OAI21X1_967 gnd vdd FILL
XFILL_1_OAI21X1_989 gnd vdd FILL
XFILL_27_2_1 gnd vdd FILL
XFILL_2_2_1 gnd vdd FILL
XFILL_0_OAI21X1_1540 gnd vdd FILL
XFILL_0_OAI21X1_1551 gnd vdd FILL
XFILL_0_OAI21X1_1584 gnd vdd FILL
XFILL_0_OAI21X1_1573 gnd vdd FILL
XFILL_0_OAI21X1_1562 gnd vdd FILL
XFILL_0_OAI21X1_1595 gnd vdd FILL
XFILL_10_1_1 gnd vdd FILL
XFILL_0_BUFX2_506 gnd vdd FILL
XFILL_0_BUFX2_517 gnd vdd FILL
XFILL_0_BUFX2_539 gnd vdd FILL
XFILL_0_BUFX2_528 gnd vdd FILL
XFILL_20_17_1 gnd vdd FILL
XCLKBUF1_9 BUFX4_84/Y gnd CLKBUF1_9/Y vdd CLKBUF1
XBUFX4_103 BUFX4_11/A gnd BUFX4_103/Y vdd BUFX4
XBUFX4_136 BUFX4_18/Y gnd BUFX4_136/Y vdd BUFX4
XBUFX4_125 BUFX4_18/Y gnd BUFX4_125/Y vdd BUFX4
XBUFX4_114 INVX8_4/Y gnd BUFX4_388/A vdd BUFX4
XFILL_0_INVX1_14 gnd vdd FILL
XFILL_0_INVX1_25 gnd vdd FILL
XFILL_4_CLKBUF1_29 gnd vdd FILL
XBUFX4_147 BUFX4_19/Y gnd BUFX4_147/Y vdd BUFX4
XNOR2X1_207 INVX1_195/A NOR2X1_207/B gnd AND2X2_32/B vdd NOR2X1
XFILL_18_2_1 gnd vdd FILL
XFILL_1_AND2X2_6 gnd vdd FILL
XFILL_0_INVX1_36 gnd vdd FILL
XFILL_4_CLKBUF1_18 gnd vdd FILL
XBUFX4_169 BUFX4_16/Y gnd BUFX4_169/Y vdd BUFX4
XFILL_0_INVX1_58 gnd vdd FILL
XFILL_0_INVX1_47 gnd vdd FILL
XBUFX4_158 BUFX4_16/Y gnd BUFX4_158/Y vdd BUFX4
XFILL_4_DFFPOSX1_390 gnd vdd FILL
XFILL_0_INVX1_69 gnd vdd FILL
XNOR2X1_218 INVX2_63/Y NOR2X1_220/B gnd INVX2_108/A vdd NOR2X1
XNOR2X1_229 INVX4_48/Y OR2X2_21/A gnd NOR2X1_229/Y vdd NOR2X1
XFILL_30_9_0 gnd vdd FILL
XFILL_25_16_1 gnd vdd FILL
XOAI21X1_1004 BUFX4_154/Y BUFX4_51/Y BUFX2_365/A gnd OAI21X1_1005/C vdd OAI21X1
XFILL_1_OAI21X1_1213 gnd vdd FILL
XFILL_1_BUFX2_291 gnd vdd FILL
XDFFPOSX1_605 BUFX2_638/A CLKBUF1_19/Y OAI21X1_826/Y gnd vdd DFFPOSX1
XOAI21X1_1037 BUFX4_376/Y INVX2_55/Y NAND2X1_403/Y gnd OAI21X1_1037/Y vdd OAI21X1
XFILL_1_OAI21X1_1202 gnd vdd FILL
XOAI21X1_1015 BUFX4_294/Y INVX1_162/Y OAI21X1_1015/C gnd OAI21X1_1015/Y vdd OAI21X1
XOAI21X1_1026 BUFX4_153/Y BUFX4_69/Y BUFX2_377/A gnd OAI21X1_1027/C vdd OAI21X1
XFILL_1_DFFPOSX1_814 gnd vdd FILL
XFILL_1_OAI21X1_1257 gnd vdd FILL
XOAI21X1_1048 BUFX4_386/Y INVX2_64/Y NAND2X1_414/Y gnd OAI21X1_1048/Y vdd OAI21X1
XFILL_1_OAI21X1_1224 gnd vdd FILL
XFILL_1_OAI21X1_1235 gnd vdd FILL
XFILL_1_OAI21X1_1246 gnd vdd FILL
XDFFPOSX1_627 INVX1_56/A CLKBUF1_67/Y OAI21X1_855/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_803 gnd vdd FILL
XDFFPOSX1_616 INVX1_45/A CLKBUF1_82/Y OAI21X1_844/Y gnd vdd DFFPOSX1
XDFFPOSX1_638 INVX1_67/A CLKBUF1_82/Y OAI21X1_866/Y gnd vdd DFFPOSX1
XOAI21X1_1059 BUFX4_326/Y INVX1_174/Y NAND2X1_425/Y gnd OAI21X1_1059/Y vdd OAI21X1
XFILL_1_OAI21X1_208 gnd vdd FILL
XFILL_1_DFFPOSX1_825 gnd vdd FILL
XDFFPOSX1_649 BUFX2_294/A CLKBUF1_64/Y OAI21X1_877/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_836 gnd vdd FILL
XFILL_1_OAI21X1_1279 gnd vdd FILL
XFILL_1_DFFPOSX1_858 gnd vdd FILL
XFILL_1_OAI21X1_1268 gnd vdd FILL
XFILL_1_DFFPOSX1_847 gnd vdd FILL
XNAND2X1_719 BUFX2_811/A BUFX4_385/Y gnd NAND2X1_719/Y vdd NAND2X1
XNAND2X1_708 BUFX2_700/A BUFX4_227/Y gnd NAND2X1_708/Y vdd NAND2X1
XFILL_1_OAI21X1_219 gnd vdd FILL
XFILL_1_DFFPOSX1_869 gnd vdd FILL
XFILL_6_DFFPOSX1_462 gnd vdd FILL
XFILL_6_DFFPOSX1_451 gnd vdd FILL
XFILL_6_DFFPOSX1_440 gnd vdd FILL
XFILL_6_DFFPOSX1_484 gnd vdd FILL
XFILL_6_DFFPOSX1_473 gnd vdd FILL
XFILL_1_NAND2X1_214 gnd vdd FILL
XFILL_1_NAND2X1_203 gnd vdd FILL
XFILL_0_DFFPOSX1_415 gnd vdd FILL
XFILL_0_DFFPOSX1_404 gnd vdd FILL
XFILL_0_17_1 gnd vdd FILL
XFILL_1_NAND2X1_258 gnd vdd FILL
XFILL_1_NAND2X1_269 gnd vdd FILL
XFILL_0_DFFPOSX1_426 gnd vdd FILL
XFILL_0_DFFPOSX1_448 gnd vdd FILL
XFILL_0_DFFPOSX1_437 gnd vdd FILL
XFILL_0_DFFPOSX1_459 gnd vdd FILL
XFILL_21_9_0 gnd vdd FILL
XFILL_5_DFFPOSX1_1020 gnd vdd FILL
XFILL_5_DFFPOSX1_1031 gnd vdd FILL
XFILL_3_DFFPOSX1_919 gnd vdd FILL
XFILL_24_11_0 gnd vdd FILL
XFILL_3_DFFPOSX1_908 gnd vdd FILL
XDFFPOSX1_20 BUFX2_689/A CLKBUF1_11/Y DFFPOSX1_20/D gnd vdd DFFPOSX1
XDFFPOSX1_53 BUFX2_722/A CLKBUF1_95/Y DFFPOSX1_53/D gnd vdd DFFPOSX1
XDFFPOSX1_31 BUFX2_701/A CLKBUF1_2/Y DFFPOSX1_31/D gnd vdd DFFPOSX1
XDFFPOSX1_42 BUFX2_741/A CLKBUF1_41/Y DFFPOSX1_42/D gnd vdd DFFPOSX1
XOAI21X1_1582 BUFX4_316/Y INVX2_118/Y NAND2X1_651/Y gnd OAI21X1_1582/Y vdd OAI21X1
XDFFPOSX1_75 BUFX2_774/A CLKBUF1_93/Y DFFPOSX1_75/D gnd vdd DFFPOSX1
XOAI21X1_1571 BUFX4_128/Y BUFX4_45/Y BUFX2_252/A gnd OAI21X1_1572/C vdd OAI21X1
XDFFPOSX1_64 BUFX2_734/A CLKBUF1_22/Y DFFPOSX1_64/D gnd vdd DFFPOSX1
XDFFPOSX1_86 BUFX2_755/A CLKBUF1_73/Y DFFPOSX1_86/D gnd vdd DFFPOSX1
XOAI21X1_1593 BUFX4_376/Y INVX2_129/Y NAND2X1_662/Y gnd OAI21X1_1593/Y vdd OAI21X1
XOAI21X1_1560 NAND2X1_646/Y BUFX4_297/Y OAI21X1_1560/C gnd OAI21X1_1560/Y vdd OAI21X1
XFILL_1_OAI21X1_1791 gnd vdd FILL
XFILL_1_OAI21X1_1780 gnd vdd FILL
XDFFPOSX1_97 BUFX2_767/A CLKBUF1_26/Y DFFPOSX1_97/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_720 gnd vdd FILL
XFILL_1_OAI21X1_764 gnd vdd FILL
XFILL_0_OAI21X1_571 gnd vdd FILL
XFILL_0_OAI21X1_582 gnd vdd FILL
XFILL_1_OAI21X1_731 gnd vdd FILL
XFILL_1_OAI21X1_742 gnd vdd FILL
XFILL_1_OAI21X1_753 gnd vdd FILL
XFILL_0_OAI21X1_560 gnd vdd FILL
XFILL_1_OAI21X1_786 gnd vdd FILL
XFILL_1_OAI21X1_797 gnd vdd FILL
XFILL_1_OAI21X1_775 gnd vdd FILL
XFILL_0_OAI21X1_593 gnd vdd FILL
XFILL_5_16_1 gnd vdd FILL
XBUFX2_618 BUFX2_618/A gnd majID4_o[24] vdd BUFX2
XFILL_2_DFFPOSX1_509 gnd vdd FILL
XBUFX2_607 BUFX2_607/A gnd majID4_o[34] vdd BUFX2
XFILL_0_CLKBUF1_60 gnd vdd FILL
XBUFX2_629 BUFX2_629/A gnd majID4_o[14] vdd BUFX2
XFILL_0_CLKBUF1_82 gnd vdd FILL
XFILL_0_CLKBUF1_71 gnd vdd FILL
XFILL_0_CLKBUF1_93 gnd vdd FILL
XFILL_29_10_0 gnd vdd FILL
XFILL_1_NAND2X1_770 gnd vdd FILL
XFILL_0_OAI21X1_1392 gnd vdd FILL
XFILL_0_OAI21X1_1381 gnd vdd FILL
XFILL_0_DFFPOSX1_960 gnd vdd FILL
XFILL_12_9_0 gnd vdd FILL
XFILL_0_OAI21X1_1370 gnd vdd FILL
XFILL_0_DFFPOSX1_982 gnd vdd FILL
XFILL_0_DFFPOSX1_993 gnd vdd FILL
XFILL_0_DFFPOSX1_971 gnd vdd FILL
XINVX2_103 INVX2_103/A gnd NOR3X1_12/B vdd INVX2
XINVX2_114 bundlePid_i[2] gnd INVX2_114/Y vdd INVX2
XFILL_0_BUFX2_314 gnd vdd FILL
XFILL_0_BUFX2_303 gnd vdd FILL
XINVX2_125 bundlePid_i[23] gnd INVX2_125/Y vdd INVX2
XFILL_0_BUFX2_325 gnd vdd FILL
XFILL_0_BUFX2_336 gnd vdd FILL
XINVX2_136 bundlePid_i[12] gnd INVX2_136/Y vdd INVX2
XFILL_0_BUFX2_347 gnd vdd FILL
XINVX2_147 bundleTid_i[62] gnd OAI21X1_9/A vdd INVX2
XINVX2_158 bundleTid_i[51] gnd INVX2_158/Y vdd INVX2
XFILL_0_BUFX2_358 gnd vdd FILL
XINVX2_169 bundleTid_i[40] gnd INVX2_169/Y vdd INVX2
XFILL_0_BUFX2_369 gnd vdd FILL
XFILL_4_11_0 gnd vdd FILL
XFILL_33_0_1 gnd vdd FILL
XFILL_0_INVX1_1 gnd vdd FILL
XFILL_22_3 gnd vdd FILL
XFILL_1_NAND3X1_10 gnd vdd FILL
XFILL_1_NAND3X1_21 gnd vdd FILL
XFILL_1_OAI21X1_1032 gnd vdd FILL
XFILL_1_OAI21X1_1021 gnd vdd FILL
XDFFPOSX1_413 BUFX2_446/A CLKBUF1_29/Y OAI21X1_385/Y gnd vdd DFFPOSX1
XFILL_1_NAND3X1_54 gnd vdd FILL
XFILL_1_NAND3X1_32 gnd vdd FILL
XDFFPOSX1_402 BUFX2_434/A CLKBUF1_80/Y OAI21X1_374/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1010 gnd vdd FILL
XFILL_1_NAND3X1_43 gnd vdd FILL
XFILL_1_OAI21X1_1043 gnd vdd FILL
XFILL_1_DFFPOSX1_633 gnd vdd FILL
XFILL_1_OAI21X1_1065 gnd vdd FILL
XFILL_1_DFFPOSX1_600 gnd vdd FILL
XFILL_1_OAI21X1_1054 gnd vdd FILL
XFILL_0_BUFX2_870 gnd vdd FILL
XFILL_1_DFFPOSX1_611 gnd vdd FILL
XFILL_1_NAND3X1_65 gnd vdd FILL
XFILL_1_DFFPOSX1_622 gnd vdd FILL
XDFFPOSX1_424 BUFX2_491/A CLKBUF1_75/Y OAI21X1_401/Y gnd vdd DFFPOSX1
XDFFPOSX1_435 BUFX2_464/A CLKBUF1_13/Y OAI21X1_422/Y gnd vdd DFFPOSX1
XDFFPOSX1_446 BUFX2_476/A CLKBUF1_33/Y OAI21X1_439/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_881 gnd vdd FILL
XFILL_1_DFFPOSX1_655 gnd vdd FILL
XDFFPOSX1_479 BUFX2_512/A CLKBUF1_29/Y OAI21X1_492/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1098 gnd vdd FILL
XDFFPOSX1_468 BUFX2_500/A CLKBUF1_72/Y OAI21X1_473/Y gnd vdd DFFPOSX1
XDFFPOSX1_457 BUFX2_488/A CLKBUF1_9/Y OAI21X1_455/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_892 gnd vdd FILL
XFILL_1_DFFPOSX1_644 gnd vdd FILL
XFILL_1_DFFPOSX1_666 gnd vdd FILL
XFILL_1_OAI21X1_1076 gnd vdd FILL
XFILL_1_OAI21X1_1087 gnd vdd FILL
XFILL_1_DFFPOSX1_688 gnd vdd FILL
XNAND2X1_516 BUFX2_83/A BUFX4_229/Y gnd NAND2X1_516/Y vdd NAND2X1
XINVX1_191 BUFX2_90/A gnd INVX1_191/Y vdd INVX1
XNAND2X1_527 bundleAddress_i[34] INVX2_98/Y gnd NOR2X1_145/A vdd NAND2X1
XINVX1_180 bundleAddress_i[6] gnd INVX1_180/Y vdd INVX1
XNAND2X1_505 bundleAddress_i[44] bundleAddress_i[43] gnd OR2X2_18/A vdd NAND2X1
XFILL_1_DFFPOSX1_677 gnd vdd FILL
XFILL_1_DFFPOSX1_699 gnd vdd FILL
XNAND2X1_549 bundleAddress_i[21] NOR2X1_160/Y gnd INVX1_194/A vdd NAND2X1
XNAND2X1_538 BUFX2_96/A INVX8_1/A gnd NAND2X1_538/Y vdd NAND2X1
XFILL_9_10_0 gnd vdd FILL
XFILL_0_INVX2_90 gnd vdd FILL
XFILL_0_AND2X2_17 gnd vdd FILL
XFILL_0_AND2X2_28 gnd vdd FILL
XFILL_10_17_0 gnd vdd FILL
XFILL_0_DFFPOSX1_212 gnd vdd FILL
XFILL_0_DFFPOSX1_201 gnd vdd FILL
XFILL_24_0_1 gnd vdd FILL
XFILL_0_DFFPOSX1_223 gnd vdd FILL
XFILL_0_DFFPOSX1_245 gnd vdd FILL
XFILL_0_DFFPOSX1_234 gnd vdd FILL
XFILL_0_DFFPOSX1_256 gnd vdd FILL
XFILL_0_DFFPOSX1_278 gnd vdd FILL
XFILL_0_DFFPOSX1_289 gnd vdd FILL
XFILL_0_DFFPOSX1_267 gnd vdd FILL
XFILL_3_DFFPOSX1_705 gnd vdd FILL
XFILL_3_DFFPOSX1_716 gnd vdd FILL
XFILL_3_DFFPOSX1_727 gnd vdd FILL
XFILL_3_DFFPOSX1_738 gnd vdd FILL
XFILL_3_CLKBUF1_15 gnd vdd FILL
XFILL_3_DFFPOSX1_749 gnd vdd FILL
XFILL_3_CLKBUF1_26 gnd vdd FILL
XFILL_3_CLKBUF1_48 gnd vdd FILL
XFILL_3_CLKBUF1_37 gnd vdd FILL
XFILL_3_CLKBUF1_59 gnd vdd FILL
XOAI21X1_1390 BUFX4_168/Y BUFX4_36/Y BUFX2_216/A gnd OAI21X1_1391/C vdd OAI21X1
XFILL_1_NOR2X1_100 gnd vdd FILL
XFILL_1_NOR2X1_122 gnd vdd FILL
XDFFPOSX1_980 BUFX2_232/A CLKBUF1_68/Y OAI21X1_1517/Y gnd vdd DFFPOSX1
XDFFPOSX1_991 BUFX2_244/A CLKBUF1_20/Y OAI21X1_1552/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_390 gnd vdd FILL
XFILL_1_OAI21X1_550 gnd vdd FILL
XFILL_7_1_1 gnd vdd FILL
XFILL_1_OAI21X1_561 gnd vdd FILL
XFILL_1_OAI21X1_572 gnd vdd FILL
XFILL_1_OAI21X1_583 gnd vdd FILL
XFILL_2_OAI21X1_776 gnd vdd FILL
XFILL_2_NAND3X1_8 gnd vdd FILL
XFILL_1_NOR2X1_188 gnd vdd FILL
XFILL_1_OAI21X1_594 gnd vdd FILL
XFILL_15_16_0 gnd vdd FILL
XFILL_2_DFFPOSX1_306 gnd vdd FILL
XFILL_2_DFFPOSX1_328 gnd vdd FILL
XBUFX2_404 BUFX2_404/A gnd majID1_o[44] vdd BUFX2
XFILL_2_DFFPOSX1_317 gnd vdd FILL
XBUFX2_426 BUFX2_426/A gnd majID1_o[24] vdd BUFX2
XBUFX2_415 BUFX2_415/A gnd majID1_o[34] vdd BUFX2
XBUFX2_448 BUFX2_448/A gnd majID1_o[4] vdd BUFX2
XFILL_2_DFFPOSX1_339 gnd vdd FILL
XBUFX2_437 BUFX2_437/A gnd majID1_o[14] vdd BUFX2
XBUFX2_459 BUFX2_459/A gnd majID2_o[53] vdd BUFX2
XFILL_15_0_1 gnd vdd FILL
XFILL_1_BUFX4_331 gnd vdd FILL
XFILL_1_BUFX4_320 gnd vdd FILL
XFILL_1_BUFX4_353 gnd vdd FILL
XFILL_1_BUFX4_342 gnd vdd FILL
XFILL_1_BUFX4_364 gnd vdd FILL
XFILL_1_BUFX4_386 gnd vdd FILL
XFILL_1_BUFX4_375 gnd vdd FILL
XFILL_0_DFFPOSX1_790 gnd vdd FILL
XFILL_0_BUFX2_122 gnd vdd FILL
XFILL_0_BUFX2_111 gnd vdd FILL
XFILL_2_OAI21X1_77 gnd vdd FILL
XFILL_0_BUFX2_100 gnd vdd FILL
XFILL_0_BUFX2_133 gnd vdd FILL
XFILL_0_BUFX2_155 gnd vdd FILL
XFILL_0_BUFX2_144 gnd vdd FILL
XFILL_0_BUFX2_199 gnd vdd FILL
XFILL_0_BUFX2_188 gnd vdd FILL
XFILL_0_BUFX2_166 gnd vdd FILL
XFILL_0_BUFX2_177 gnd vdd FILL
XFILL_1_DFFPOSX1_9 gnd vdd FILL
XFILL_33_17_0 gnd vdd FILL
XFILL_35_8_0 gnd vdd FILL
XFILL_2_DFFPOSX1_840 gnd vdd FILL
XFILL_2_DFFPOSX1_851 gnd vdd FILL
XFILL_2_OAI21X1_1283 gnd vdd FILL
XFILL_2_DFFPOSX1_884 gnd vdd FILL
XBUFX2_982 BUFX2_982/A gnd tid4_o[43] vdd BUFX2
XFILL_2_DFFPOSX1_873 gnd vdd FILL
XBUFX2_960 BUFX2_960/A gnd tid3_o[4] vdd BUFX2
XBUFX2_971 BUFX2_971/A gnd tid4_o[53] vdd BUFX2
XFILL_2_DFFPOSX1_862 gnd vdd FILL
XBUFX2_993 BUFX2_993/A gnd tid4_o[33] vdd BUFX2
XFILL_2_DFFPOSX1_895 gnd vdd FILL
XOAI21X1_307 INVX2_199/Y BUFX4_301/Y OAI21X1_307/C gnd OAI21X1_307/Y vdd OAI21X1
XOAI21X1_329 INVX2_8/Y BUFX4_321/Y NAND2X1_73/Y gnd OAI21X1_329/Y vdd OAI21X1
XOAI21X1_318 BUFX4_169/Y BUFX4_80/A BUFX2_1024/A gnd OAI21X1_319/C vdd OAI21X1
XDFFPOSX1_221 BUFX2_894/A CLKBUF1_47/Y OAI21X1_65/Y gnd vdd DFFPOSX1
XBUFX4_5 BUFX4_6/A gnd BUFX4_5/Y vdd BUFX4
XDFFPOSX1_210 BUFX2_882/A CLKBUF1_4/Y OAI21X1_54/Y gnd vdd DFFPOSX1
XDFFPOSX1_232 BUFX2_939/A CLKBUF1_74/Y OAI21X1_81/Y gnd vdd DFFPOSX1
XDFFPOSX1_254 BUFX2_924/A CLKBUF1_3/Y OAI21X1_125/Y gnd vdd DFFPOSX1
XDFFPOSX1_243 BUFX2_912/A CLKBUF1_12/Y OAI21X1_103/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_430 gnd vdd FILL
XFILL_1_DFFPOSX1_441 gnd vdd FILL
XFILL_38_16_0 gnd vdd FILL
XDFFPOSX1_276 BUFX2_948/A CLKBUF1_14/Y OAI21X1_169/Y gnd vdd DFFPOSX1
XDFFPOSX1_265 BUFX2_936/A CLKBUF1_70/Y OAI21X1_147/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_463 gnd vdd FILL
XNAND2X1_302 INVX1_21/Y NOR2X1_95/Y gnd OR2X2_12/A vdd NAND2X1
XDFFPOSX1_298 BUFX2_1025/A CLKBUF1_60/Y OAI21X1_213/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_452 gnd vdd FILL
XDFFPOSX1_287 BUFX2_960/A CLKBUF1_51/Y OAI21X1_191/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_474 gnd vdd FILL
XNAND2X1_335 bundleStartMajId_i[3] NOR3X1_10/Y gnd OAI21X1_839/A vdd NAND2X1
XFILL_3_NOR3X1_18 gnd vdd FILL
XNAND2X1_324 NOR2X1_105/Y NOR2X1_30/Y gnd OR2X2_15/A vdd NAND2X1
XFILL_1_DFFPOSX1_485 gnd vdd FILL
XNAND2X1_313 AND2X2_12/Y AND2X2_20/A gnd OAI21X1_698/C vdd NAND2X1
XFILL_1_DFFPOSX1_496 gnd vdd FILL
XNAND2X1_346 BUFX4_263/Y bundle_i[23] gnd OAI21X1_852/C vdd NAND2X1
XFILL_4_DFFPOSX1_901 gnd vdd FILL
XFILL_4_DFFPOSX1_923 gnd vdd FILL
XNAND2X1_357 BUFX4_261/Y bundle_i[12] gnd OAI21X1_863/C vdd NAND2X1
XNAND2X1_368 BUFX4_268/Y bundle_i[1] gnd OAI21X1_874/C vdd NAND2X1
XFILL_4_DFFPOSX1_912 gnd vdd FILL
XFILL_4_DFFPOSX1_945 gnd vdd FILL
XFILL_4_DFFPOSX1_934 gnd vdd FILL
XFILL_4_DFFPOSX1_956 gnd vdd FILL
XNAND2X1_379 BUFX2_324/A BUFX4_232/Y gnd OAI21X1_885/C vdd NAND2X1
XFILL_4_DFFPOSX1_967 gnd vdd FILL
XFILL_4_DFFPOSX1_978 gnd vdd FILL
XFILL_4_DFFPOSX1_989 gnd vdd FILL
XFILL_26_8_0 gnd vdd FILL
XFILL_1_8_0 gnd vdd FILL
XFILL_0_XNOR2X1_1 gnd vdd FILL
XFILL_1_BUFX2_824 gnd vdd FILL
XINVX4_5 bundleStartMajId_i[51] gnd INVX4_5/Y vdd INVX4
XFILL_1_BUFX2_835 gnd vdd FILL
XFILL_1_BUFX2_868 gnd vdd FILL
XFILL_1_BUFX2_879 gnd vdd FILL
XOAI21X1_830 OAI21X1_830/A BUFX4_289/Y OAI21X1_830/C gnd OAI21X1_830/Y vdd OAI21X1
XOAI21X1_841 BUFX4_155/Y BUFX4_61/Y BUFX2_645/A gnd OAI21X1_843/C vdd OAI21X1
XFILL_3_DFFPOSX1_513 gnd vdd FILL
XFILL_3_DFFPOSX1_502 gnd vdd FILL
XFILL_3_DFFPOSX1_546 gnd vdd FILL
XOAI21X1_852 INVX1_53/Y BUFX4_265/Y OAI21X1_852/C gnd OAI21X1_852/Y vdd OAI21X1
XFILL_3_DFFPOSX1_535 gnd vdd FILL
XFILL_3_DFFPOSX1_524 gnd vdd FILL
XOAI21X1_874 INVX1_75/Y BUFX4_268/Y OAI21X1_874/C gnd OAI21X1_874/Y vdd OAI21X1
XOAI21X1_863 INVX1_64/Y BUFX4_267/Y OAI21X1_863/C gnd OAI21X1_863/Y vdd OAI21X1
XOAI21X1_885 INVX1_86/Y BUFX4_232/Y OAI21X1_885/C gnd OAI21X1_885/Y vdd OAI21X1
XOAI21X1_896 INVX1_97/Y BUFX4_184/Y OAI21X1_896/C gnd OAI21X1_896/Y vdd OAI21X1
XFILL_3_DFFPOSX1_568 gnd vdd FILL
XFILL_3_DFFPOSX1_579 gnd vdd FILL
XFILL_3_DFFPOSX1_557 gnd vdd FILL
XFILL_9_9_0 gnd vdd FILL
XFILL_1_OAI21X1_380 gnd vdd FILL
XFILL_1_CLKBUF1_1 gnd vdd FILL
XFILL_1_OAI21X1_391 gnd vdd FILL
XBUFX2_201 BUFX2_201/A gnd addr4_o[47] vdd BUFX2
XFILL_2_DFFPOSX1_103 gnd vdd FILL
XFILL_2_DFFPOSX1_114 gnd vdd FILL
XFILL_2_DFFPOSX1_125 gnd vdd FILL
XBUFX2_212 BUFX2_212/A gnd addr4_o[37] vdd BUFX2
XFILL_2_DFFPOSX1_136 gnd vdd FILL
XBUFX2_234 BUFX2_234/A gnd addr4_o[17] vdd BUFX2
XFILL_0_NAND3X1_40 gnd vdd FILL
XFILL_0_NAND3X1_62 gnd vdd FILL
XFILL_17_8_0 gnd vdd FILL
XFILL_0_NAND3X1_51 gnd vdd FILL
XFILL_0_NAND2X1_609 gnd vdd FILL
XBUFX2_223 BUFX2_223/A gnd addr4_o[27] vdd BUFX2
XBUFX2_278 INVX1_69/A gnd instr1_o[7] vdd BUFX2
XBUFX2_267 INVX1_59/A gnd instr1_o[17] vdd BUFX2
XFILL_2_DFFPOSX1_147 gnd vdd FILL
XBUFX2_256 BUFX2_256/A gnd addr4_o[54] vdd BUFX2
XFILL_2_DFFPOSX1_158 gnd vdd FILL
XFILL_2_DFFPOSX1_169 gnd vdd FILL
XBUFX2_245 BUFX2_245/A gnd addr4_o[7] vdd BUFX2
XBUFX2_289 INVX1_51/A gnd instr1_o[25] vdd BUFX2
XFILL_5_DFFPOSX1_607 gnd vdd FILL
XFILL_5_DFFPOSX1_618 gnd vdd FILL
XFILL_1_BUFX4_172 gnd vdd FILL
XFILL_1_BUFX4_150 gnd vdd FILL
XFILL_1_BUFX4_161 gnd vdd FILL
XFILL_5_DFFPOSX1_629 gnd vdd FILL
XFILL_1_BUFX4_183 gnd vdd FILL
XFILL_1_BUFX4_194 gnd vdd FILL
XFILL_22_14_1 gnd vdd FILL
XFILL_4_DFFPOSX1_208 gnd vdd FILL
XNAND3X1_8 bundleStartMajId_i[23] bundleStartMajId_i[22] bundleStartMajId_i[21] gnd
+ NOR3X1_3/A vdd NAND3X1
XFILL_4_DFFPOSX1_219 gnd vdd FILL
XFILL_2_CLKBUF1_12 gnd vdd FILL
XFILL_2_CLKBUF1_23 gnd vdd FILL
XFILL_2_CLKBUF1_45 gnd vdd FILL
XFILL_2_CLKBUF1_34 gnd vdd FILL
XFILL_2_CLKBUF1_56 gnd vdd FILL
XFILL_2_CLKBUF1_67 gnd vdd FILL
XFILL_2_CLKBUF1_89 gnd vdd FILL
XFILL_2_CLKBUF1_78 gnd vdd FILL
XFILL_2_DFFPOSX1_670 gnd vdd FILL
XFILL_2_DFFPOSX1_692 gnd vdd FILL
XFILL_2_DFFPOSX1_681 gnd vdd FILL
XBUFX2_790 BUFX2_790/A gnd tid1_o[43] vdd BUFX2
XFILL_0_NOR2X1_130 gnd vdd FILL
XFILL_27_13_1 gnd vdd FILL
XOAI21X1_104 BUFX4_108/Y BUFX4_334/Y BUFX2_913/A gnd OAI21X1_105/C vdd OAI21X1
XFILL_0_NOR2X1_163 gnd vdd FILL
XFILL_0_NOR2X1_152 gnd vdd FILL
XFILL_0_NOR2X1_141 gnd vdd FILL
XFILL_1_BUFX2_109 gnd vdd FILL
XOAI21X1_126 BUFX4_11/A BUFX4_332/Y BUFX2_925/A gnd OAI21X1_127/C vdd OAI21X1
XOAI21X1_115 BUFX4_136/Y INVX2_167/Y OAI21X1_115/C gnd OAI21X1_115/Y vdd OAI21X1
XFILL_0_NOR2X1_185 gnd vdd FILL
XFILL_0_NOR2X1_196 gnd vdd FILL
XFILL_0_NOR2X1_174 gnd vdd FILL
XOAI21X1_137 BUFX4_173/Y INVX2_178/Y OAI21X1_137/C gnd OAI21X1_137/Y vdd OAI21X1
XOAI21X1_159 BUFX4_172/Y INVX2_189/Y OAI21X1_159/C gnd OAI21X1_159/Y vdd OAI21X1
XOAI21X1_148 BUFX4_11/A BUFX4_322/Y BUFX2_937/A gnd OAI21X1_149/C vdd OAI21X1
XFILL_0_DFFPOSX1_1004 gnd vdd FILL
XFILL_0_DFFPOSX1_1026 gnd vdd FILL
XFILL_0_DFFPOSX1_1015 gnd vdd FILL
XBUFX2_2 BUFX2_2/A gnd addr1_o[62] vdd BUFX2
XFILL_1_DFFPOSX1_282 gnd vdd FILL
XFILL_1_DFFPOSX1_271 gnd vdd FILL
XNAND2X1_110 BUFX2_425/A BUFX4_351/Y gnd OAI21X1_366/C vdd NAND2X1
XFILL_1_DFFPOSX1_260 gnd vdd FILL
XNAND2X1_132 BUFX2_450/A BUFX4_351/Y gnd OAI21X1_388/C vdd NAND2X1
XNAND2X1_121 BUFX2_437/A BUFX4_323/Y gnd OAI21X1_377/C vdd NAND2X1
XNAND2X1_143 bundleStartMajId_i[59] NOR2X1_3/Y gnd INVX1_8/A vdd NAND2X1
XFILL_1_DFFPOSX1_293 gnd vdd FILL
XNAND2X1_176 BUFX2_468/A BUFX4_224/Y gnd OAI21X1_429/C vdd NAND2X1
XNAND2X1_187 NOR2X1_16/Y NOR2X1_11/Y gnd NOR3X1_1/C vdd NAND2X1
XNAND2X1_154 BUFX2_520/A BUFX4_181/Y gnd OAI21X1_412/C vdd NAND2X1
XFILL_4_DFFPOSX1_720 gnd vdd FILL
XFILL_4_DFFPOSX1_731 gnd vdd FILL
XNAND2X1_165 bundleStartMajId_i[51] bundleStartMajId_i[48] gnd NOR2X1_10/A vdd NAND2X1
XFILL_1_OAI21X1_52 gnd vdd FILL
XFILL_4_DFFPOSX1_742 gnd vdd FILL
XFILL_1_OAI21X1_41 gnd vdd FILL
XFILL_4_DFFPOSX1_753 gnd vdd FILL
XFILL_1_OAI21X1_30 gnd vdd FILL
XFILL_0_XNOR2X1_19 gnd vdd FILL
XNAND2X1_198 BUFX2_479/A BUFX4_214/Y gnd OAI21X1_444/C vdd NAND2X1
XFILL_4_DFFPOSX1_764 gnd vdd FILL
XFILL_1_OAI21X1_85 gnd vdd FILL
XFILL_4_DFFPOSX1_775 gnd vdd FILL
XFILL_1_OAI21X1_74 gnd vdd FILL
XFILL_1_OAI21X1_63 gnd vdd FILL
XFILL_4_DFFPOSX1_786 gnd vdd FILL
XFILL_4_DFFPOSX1_797 gnd vdd FILL
XFILL_2_14_1 gnd vdd FILL
XFILL_1_OAI21X1_96 gnd vdd FILL
XFILL_0_DFFPOSX1_6 gnd vdd FILL
XFILL_1_BUFX2_621 gnd vdd FILL
XFILL_1_BUFX2_643 gnd vdd FILL
XFILL_1_BUFX2_632 gnd vdd FILL
XINVX2_2 bundleTid_i[5] gnd INVX2_2/Y vdd INVX2
XFILL_0_BUFX4_206 gnd vdd FILL
XFILL_1_BUFX2_665 gnd vdd FILL
XFILL_1_BUFX2_687 gnd vdd FILL
XFILL_3_DFFPOSX1_321 gnd vdd FILL
XFILL_3_DFFPOSX1_310 gnd vdd FILL
XFILL_0_BUFX4_239 gnd vdd FILL
XFILL_0_BUFX4_228 gnd vdd FILL
XFILL_1_BUFX2_676 gnd vdd FILL
XOAI21X1_660 BUFX4_131/Y BUFX4_61/Y BUFX2_586/A gnd OAI21X1_661/C vdd OAI21X1
XFILL_0_BUFX4_217 gnd vdd FILL
XFILL_1_OAI21X1_1609 gnd vdd FILL
XAOI21X1_2 bundleStartMajId_i[33] NOR3X1_1/Y INVX2_24/Y gnd AOI21X1_2/Y vdd AOI21X1
XFILL_3_DFFPOSX1_343 gnd vdd FILL
XOAI21X1_671 XNOR2X1_40/Y BUFX4_302/Y OAI21X1_671/C gnd OAI21X1_671/Y vdd OAI21X1
XFILL_3_DFFPOSX1_354 gnd vdd FILL
XFILL_3_DFFPOSX1_332 gnd vdd FILL
XOAI21X1_693 AND2X2_19/A bundleStartMajId_i[51] BUFX4_285/Y gnd OAI21X1_695/B vdd
+ OAI21X1
XOAI21X1_682 BUFX4_167/Y BUFX4_33/Y BUFX2_647/A gnd OAI21X1_683/C vdd OAI21X1
XFILL_3_DFFPOSX1_398 gnd vdd FILL
XFILL_3_DFFPOSX1_365 gnd vdd FILL
XFILL_3_DFFPOSX1_376 gnd vdd FILL
XFILL_3_DFFPOSX1_387 gnd vdd FILL
XFILL_0_INVX4_25 gnd vdd FILL
XFILL_0_INVX4_14 gnd vdd FILL
XFILL_0_INVX4_36 gnd vdd FILL
XFILL_3_DFFPOSX1_1019 gnd vdd FILL
XFILL_0_INVX4_47 gnd vdd FILL
XXNOR2X1_21 XNOR2X1_21/A INVX2_34/Y gnd XNOR2X1_21/Y vdd XNOR2X1
XXNOR2X1_32 NOR2X1_70/B INVX4_11/Y gnd XNOR2X1_32/Y vdd XNOR2X1
XFILL_6_DFFPOSX1_869 gnd vdd FILL
XFILL_3_DFFPOSX1_1008 gnd vdd FILL
XFILL_6_DFFPOSX1_858 gnd vdd FILL
XXNOR2X1_10 NOR2X1_17/Y bundleStartMajId_i[38] gnd XNOR2X1_10/Y vdd XNOR2X1
XXNOR2X1_65 XNOR2X1_65/A bundleAddress_i[35] gnd XNOR2X1_65/Y vdd XNOR2X1
XXNOR2X1_43 INVX1_36/A INVX4_7/Y gnd XNOR2X1_43/Y vdd XNOR2X1
XXNOR2X1_54 NOR3X1_8/Y bundleStartMajId_i[10] gnd XNOR2X1_54/Y vdd XNOR2X1
XFILL_7_13_1 gnd vdd FILL
XXNOR2X1_76 INVX1_201/A INVX4_33/Y gnd XNOR2X1_76/Y vdd XNOR2X1
XXNOR2X1_98 XNOR2X1_98/A INVX2_72/Y gnd XNOR2X1_98/Y vdd XNOR2X1
XFILL_2_OAI21X1_381 gnd vdd FILL
XXNOR2X1_87 XNOR2X1_87/A bundleAddress_i[10] gnd XNOR2X1_87/Y vdd XNOR2X1
XFILL_0_NAND2X1_417 gnd vdd FILL
XFILL_0_NAND2X1_406 gnd vdd FILL
XBUFX2_20 BUFX2_20/A gnd addr1_o[37] vdd BUFX2
XBUFX2_42 BUFX2_42/A gnd addr1_o[17] vdd BUFX2
XFILL_0_NAND2X1_428 gnd vdd FILL
XBUFX2_53 BUFX2_53/A gnd addr1_o[7] vdd BUFX2
XFILL_0_NAND2X1_439 gnd vdd FILL
XBUFX2_31 BUFX2_31/A gnd addr1_o[27] vdd BUFX2
XBUFX2_64 BUFX2_64/A gnd addr1_o[54] vdd BUFX2
XBUFX2_86 BUFX2_86/A gnd addr2_o[35] vdd BUFX2
XBUFX2_75 BUFX2_75/A gnd addr2_o[45] vdd BUFX2
XFILL_32_6_0 gnd vdd FILL
XBUFX2_97 BUFX2_97/A gnd addr2_o[25] vdd BUFX2
XFILL_5_DFFPOSX1_415 gnd vdd FILL
XFILL_5_DFFPOSX1_404 gnd vdd FILL
XFILL_5_DFFPOSX1_426 gnd vdd FILL
XFILL_5_DFFPOSX1_459 gnd vdd FILL
XFILL_1_BUFX4_20 gnd vdd FILL
XFILL_5_DFFPOSX1_448 gnd vdd FILL
XFILL_5_DFFPOSX1_437 gnd vdd FILL
XFILL_1_BUFX4_42 gnd vdd FILL
XFILL_1_BUFX4_53 gnd vdd FILL
XFILL_1_BUFX4_31 gnd vdd FILL
XFILL_1_BUFX4_97 gnd vdd FILL
XFILL_1_BUFX4_75 gnd vdd FILL
XFILL_1_BUFX4_64 gnd vdd FILL
XFILL_1_BUFX4_86 gnd vdd FILL
XFILL_0_AOI21X1_19 gnd vdd FILL
XFILL_0_OAI21X1_923 gnd vdd FILL
XFILL_0_OAI21X1_901 gnd vdd FILL
XFILL_0_OAI21X1_912 gnd vdd FILL
XFILL_0_OAI21X1_956 gnd vdd FILL
XFILL_0_OAI21X1_945 gnd vdd FILL
XFILL_0_OAI21X1_934 gnd vdd FILL
XFILL_0_OAI21X1_978 gnd vdd FILL
XFILL_0_OAI21X1_967 gnd vdd FILL
XFILL_0_OAI21X1_989 gnd vdd FILL
XFILL_2_BUFX4_137 gnd vdd FILL
XFILL_0_OAI21X1_1700 gnd vdd FILL
XFILL_1_OR2X2_12 gnd vdd FILL
XFILL_0_OAI21X1_1711 gnd vdd FILL
XFILL_0_OAI21X1_1733 gnd vdd FILL
XFILL_0_OAI21X1_1722 gnd vdd FILL
XFILL_0_OAI21X1_1755 gnd vdd FILL
XFILL_0_OAI21X1_1744 gnd vdd FILL
XFILL_0_OAI21X1_1766 gnd vdd FILL
XFILL_23_6_0 gnd vdd FILL
XFILL_0_OAI21X1_1777 gnd vdd FILL
XFILL_0_OAI21X1_1788 gnd vdd FILL
XFILL_0_OAI21X1_1799 gnd vdd FILL
XFILL_5_DFFPOSX1_982 gnd vdd FILL
XFILL_5_DFFPOSX1_960 gnd vdd FILL
XAOI21X1_10 INVX1_30/Y NOR2X1_80/Y INVX4_18/Y gnd AOI21X1_10/Y vdd AOI21X1
XFILL_5_DFFPOSX1_971 gnd vdd FILL
XAOI21X1_21 INVX2_46/A NOR2X1_95/Y bundleStartMajId_i[8] gnd AOI21X1_21/Y vdd AOI21X1
XAOI21X1_32 INVX1_12/A NOR2X1_109/Y bundleStartMajId_i[37] gnd AOI21X1_32/Y vdd AOI21X1
XFILL_0_NOR2X1_28 gnd vdd FILL
XFILL_0_NOR2X1_39 gnd vdd FILL
XFILL_5_DFFPOSX1_993 gnd vdd FILL
XFILL_0_NOR2X1_17 gnd vdd FILL
XAOI21X1_43 INVX2_104/A NOR3X1_14/Y bundleAddress_i[6] gnd AOI21X1_43/Y vdd AOI21X1
XAOI21X1_54 bundleAddress_i[14] INVX1_213/Y bundleAddress_i[13] gnd AOI21X1_54/Y vdd
+ AOI21X1
XAOI21X1_65 bundleAddress_i[4] INVX2_112/Y bundleAddress_i[3] gnd AOI21X1_65/Y vdd
+ AOI21X1
XOAI21X1_5 OAI21X1_5/A INVX2_5/Y OAI21X1_5/C gnd OAI21X1_5/Y vdd OAI21X1
XFILL_18_18_1 gnd vdd FILL
XXNOR2X1_102 INVX2_110/A bundleAddress_i[20] gnd XNOR2X1_102/Y vdd XNOR2X1
XFILL_6_7_0 gnd vdd FILL
XBUFX4_318 BUFX4_381/A gnd BUFX4_318/Y vdd BUFX4
XBUFX4_307 BUFX4_310/A gnd MUX2X1_2/S vdd BUFX4
XBUFX4_329 BUFX4_376/A gnd BUFX4_329/Y vdd BUFX4
XFILL_4_DFFPOSX1_550 gnd vdd FILL
XFILL_4_DFFPOSX1_572 gnd vdd FILL
XFILL_4_DFFPOSX1_561 gnd vdd FILL
XFILL_4_DFFPOSX1_583 gnd vdd FILL
XFILL_4_DFFPOSX1_594 gnd vdd FILL
XFILL_12_14_0 gnd vdd FILL
XFILL_14_6_0 gnd vdd FILL
XFILL_1_BUFX2_1030 gnd vdd FILL
XFILL_1_BUFX2_440 gnd vdd FILL
XOAI21X1_1208 BUFX4_104/Y BUFX4_336/Y BUFX2_129/A gnd OAI21X1_1209/C vdd OAI21X1
XOAI21X1_1219 BUFX4_2/Y BUFX4_382/Y BUFX2_174/A gnd OAI21X1_1220/C vdd OAI21X1
XFILL_1_OAI21X1_1406 gnd vdd FILL
XFILL_1_CLKBUF1_31 gnd vdd FILL
XFILL_1_CLKBUF1_20 gnd vdd FILL
XFILL_1_BUFX2_473 gnd vdd FILL
XFILL_1_BUFX2_484 gnd vdd FILL
XOAI21X1_490 XNOR2X1_23/Y BUFX4_231/Y OAI21X1_490/C gnd OAI21X1_490/Y vdd OAI21X1
XFILL_1_CLKBUF1_42 gnd vdd FILL
XFILL_1_OAI21X1_1417 gnd vdd FILL
XFILL_1_OAI21X1_1428 gnd vdd FILL
XFILL_1_CLKBUF1_64 gnd vdd FILL
XFILL_3_DFFPOSX1_173 gnd vdd FILL
XDFFPOSX1_809 BUFX2_66/A CLKBUF1_78/Y OAI21X1_1101/Y gnd vdd DFFPOSX1
XFILL_3_DFFPOSX1_151 gnd vdd FILL
XFILL_1_INVX8_4 gnd vdd FILL
XFILL_1_OAI21X1_1439 gnd vdd FILL
XFILL_3_DFFPOSX1_162 gnd vdd FILL
XFILL_3_DFFPOSX1_140 gnd vdd FILL
XFILL_1_CLKBUF1_53 gnd vdd FILL
XFILL_0_OAI21X1_208 gnd vdd FILL
XFILL_1_CLKBUF1_86 gnd vdd FILL
XFILL_0_OAI21X1_219 gnd vdd FILL
XFILL_3_DFFPOSX1_195 gnd vdd FILL
XFILL_1_CLKBUF1_97 gnd vdd FILL
XFILL_3_DFFPOSX1_184 gnd vdd FILL
XFILL_1_CLKBUF1_75 gnd vdd FILL
XFILL_6_DFFPOSX1_611 gnd vdd FILL
XFILL_6_DFFPOSX1_633 gnd vdd FILL
XFILL_6_DFFPOSX1_644 gnd vdd FILL
XFILL_6_DFFPOSX1_622 gnd vdd FILL
XFILL_6_DFFPOSX1_655 gnd vdd FILL
XFILL_17_13_0 gnd vdd FILL
XFILL_6_DFFPOSX1_666 gnd vdd FILL
XFILL_30_15_0 gnd vdd FILL
XFILL_0_NAND2X1_214 gnd vdd FILL
XFILL_0_NAND2X1_225 gnd vdd FILL
XFILL_0_NAND2X1_203 gnd vdd FILL
XFILL_0_OAI21X1_1029 gnd vdd FILL
XFILL_1_NAND2X1_407 gnd vdd FILL
XFILL_1_NAND2X1_418 gnd vdd FILL
XFILL_0_OAI21X1_1007 gnd vdd FILL
XFILL_1_NAND2X1_429 gnd vdd FILL
XFILL_0_NAND2X1_258 gnd vdd FILL
XFILL_0_NAND2X1_236 gnd vdd FILL
XFILL_0_OAI21X1_1018 gnd vdd FILL
XFILL_0_NAND2X1_247 gnd vdd FILL
XFILL_38_1 gnd vdd FILL
XFILL_0_DFFPOSX1_608 gnd vdd FILL
XFILL_0_NAND2X1_269 gnd vdd FILL
XFILL_0_DFFPOSX1_619 gnd vdd FILL
XFILL_5_DFFPOSX1_201 gnd vdd FILL
XFILL_5_DFFPOSX1_245 gnd vdd FILL
XFILL_5_DFFPOSX1_212 gnd vdd FILL
XFILL_5_DFFPOSX1_234 gnd vdd FILL
XFILL_5_DFFPOSX1_223 gnd vdd FILL
XFILL_5_DFFPOSX1_278 gnd vdd FILL
XFILL_5_DFFPOSX1_267 gnd vdd FILL
XFILL_5_DFFPOSX1_256 gnd vdd FILL
XFILL_5_DFFPOSX1_289 gnd vdd FILL
XFILL_0_OAI21X1_60 gnd vdd FILL
XOAI21X1_1742 BUFX4_126/Y BUFX4_29/Y BUFX2_753/A gnd OAI21X1_1743/C vdd OAI21X1
XOAI21X1_1731 INVX2_127/Y BUFX4_293/Y OAI21X1_1731/C gnd DFFPOSX1_78/D vdd OAI21X1
XFILL_0_OAI21X1_93 gnd vdd FILL
XFILL_0_OAI21X1_71 gnd vdd FILL
XFILL_0_OAI21X1_82 gnd vdd FILL
XOAI21X1_1720 BUFX4_139/Y BUFX4_73/Y BUFX2_772/A gnd OAI21X1_1721/C vdd OAI21X1
XOAI21X1_1764 BUFX4_149/Y BUFX4_44/Y BUFX2_765/A gnd OAI21X1_1765/C vdd OAI21X1
XOAI21X1_1753 INVX2_138/Y BUFX4_296/Y OAI21X1_1753/C gnd DFFPOSX1_89/D vdd OAI21X1
XOAI21X1_1775 BUFX4_343/Y OAI21X1_9/A NAND2X1_716/Y gnd OAI21X1_1775/Y vdd OAI21X1
XOAI21X1_1786 BUFX4_322/Y INVX2_158/Y NAND2X1_727/Y gnd OAI21X1_1786/Y vdd OAI21X1
XOAI21X1_1797 BUFX4_375/Y INVX2_169/Y NAND2X1_738/Y gnd OAI21X1_1797/Y vdd OAI21X1
XFILL_0_OAI21X1_731 gnd vdd FILL
XFILL_0_OAI21X1_720 gnd vdd FILL
XFILL_1_OAI21X1_902 gnd vdd FILL
XFILL_1_OAI21X1_913 gnd vdd FILL
XFILL_1_OAI21X1_924 gnd vdd FILL
XFILL_0_OAI21X1_764 gnd vdd FILL
XFILL_0_OAI21X1_775 gnd vdd FILL
XFILL_0_OAI21X1_742 gnd vdd FILL
XFILL_0_OAI21X1_753 gnd vdd FILL
XFILL_1_OAI21X1_935 gnd vdd FILL
XFILL_1_OAI21X1_946 gnd vdd FILL
XFILL_1_OAI21X1_957 gnd vdd FILL
XFILL_1_OAI21X1_979 gnd vdd FILL
XFILL_1_OAI21X1_968 gnd vdd FILL
XFILL_35_14_0 gnd vdd FILL
XFILL_0_OAI21X1_786 gnd vdd FILL
XFILL_0_OAI21X1_797 gnd vdd FILL
XFILL_1_OR2X2_9 gnd vdd FILL
XFILL_2_NAND3X1_25 gnd vdd FILL
XFILL_0_OAI21X1_1530 gnd vdd FILL
XFILL_0_NAND2X1_770 gnd vdd FILL
XFILL_2_BUFX4_7 gnd vdd FILL
XFILL_0_OAI21X1_1541 gnd vdd FILL
XFILL_0_OAI21X1_1552 gnd vdd FILL
XFILL_0_OAI21X1_1574 gnd vdd FILL
XFILL_0_OAI21X1_1563 gnd vdd FILL
XFILL_0_OAI21X1_1585 gnd vdd FILL
XFILL_0_OAI21X1_1596 gnd vdd FILL
XFILL_5_DFFPOSX1_790 gnd vdd FILL
XFILL_0_BUFX2_518 gnd vdd FILL
XFILL_0_BUFX2_529 gnd vdd FILL
XFILL_0_BUFX2_507 gnd vdd FILL
XBUFX4_137 BUFX4_14/Y gnd BUFX4_137/Y vdd BUFX4
XBUFX4_126 BUFX4_18/Y gnd BUFX4_126/Y vdd BUFX4
XFILL_2_OAI21X1_1613 gnd vdd FILL
XBUFX4_115 INVX8_4/Y gnd BUFX4_376/A vdd BUFX4
XBUFX4_104 BUFX4_95/A gnd BUFX4_104/Y vdd BUFX4
XFILL_0_INVX1_15 gnd vdd FILL
XBUFX4_148 BUFX4_15/Y gnd BUFX4_148/Y vdd BUFX4
XBUFX4_159 BUFX4_15/Y gnd BUFX4_159/Y vdd BUFX4
XFILL_4_CLKBUF1_19 gnd vdd FILL
XFILL_0_INVX1_37 gnd vdd FILL
XFILL_1_AND2X2_7 gnd vdd FILL
XFILL_0_INVX1_26 gnd vdd FILL
XFILL_0_INVX1_48 gnd vdd FILL
XFILL_4_DFFPOSX1_391 gnd vdd FILL
XFILL_4_DFFPOSX1_380 gnd vdd FILL
XFILL_0_INVX1_59 gnd vdd FILL
XFILL_2_OAI21X1_1679 gnd vdd FILL
XNOR2X1_219 INVX2_66/Y INVX1_220/A gnd INVX1_221/A vdd NOR2X1
XNOR2X1_208 NOR3X1_12/B NOR2X1_211/B gnd XNOR2X1_87/A vdd NOR2X1
XFILL_30_9_1 gnd vdd FILL
XFILL_1_BUFX2_270 gnd vdd FILL
XFILL_1_BUFX2_281 gnd vdd FILL
XFILL_1_OAI21X1_1214 gnd vdd FILL
XFILL_1_OAI21X1_1203 gnd vdd FILL
XOAI21X1_1016 BUFX4_133/Y BUFX4_27/Y BUFX2_372/A gnd OAI21X1_1017/C vdd OAI21X1
XFILL_1_BUFX2_292 gnd vdd FILL
XOAI21X1_1027 BUFX4_302/Y INVX1_168/Y OAI21X1_1027/C gnd OAI21X1_1027/Y vdd OAI21X1
XOAI21X1_1005 BUFX4_303/Y INVX1_157/Y OAI21X1_1005/C gnd OAI21X1_1005/Y vdd OAI21X1
XFILL_1_DFFPOSX1_815 gnd vdd FILL
XOAI21X1_1038 INVX4_32/Y BUFX4_353/Y NAND2X1_404/Y gnd OAI21X1_1038/Y vdd OAI21X1
XDFFPOSX1_639 INVX1_68/A CLKBUF1_96/Y OAI21X1_867/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1236 gnd vdd FILL
XFILL_1_OAI21X1_1225 gnd vdd FILL
XOAI21X1_1049 BUFX4_340/Y INVX2_65/Y NAND2X1_415/Y gnd OAI21X1_1049/Y vdd OAI21X1
XFILL_1_OAI21X1_1247 gnd vdd FILL
XDFFPOSX1_606 BUFX2_639/A CLKBUF1_5/Y OAI21X1_830/Y gnd vdd DFFPOSX1
XDFFPOSX1_617 INVX1_46/A CLKBUF1_87/Y OAI21X1_845/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_804 gnd vdd FILL
XDFFPOSX1_628 INVX1_57/A CLKBUF1_71/Y OAI21X1_856/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1258 gnd vdd FILL
XFILL_1_DFFPOSX1_837 gnd vdd FILL
XFILL_1_OAI21X1_1269 gnd vdd FILL
XFILL_1_DFFPOSX1_848 gnd vdd FILL
XFILL_1_DFFPOSX1_826 gnd vdd FILL
XFILL_1_OAI21X1_209 gnd vdd FILL
XNAND2X1_709 BUFX2_701/A BUFX4_190/Y gnd NAND2X1_709/Y vdd NAND2X1
XFILL_1_DFFPOSX1_859 gnd vdd FILL
XFILL_37_5_0 gnd vdd FILL
XFILL_1_NAND2X1_204 gnd vdd FILL
XFILL_0_DFFPOSX1_405 gnd vdd FILL
XFILL_1_NAND2X1_237 gnd vdd FILL
XFILL_1_NAND2X1_226 gnd vdd FILL
XFILL_0_DFFPOSX1_416 gnd vdd FILL
XFILL_0_DFFPOSX1_427 gnd vdd FILL
XFILL_0_DFFPOSX1_438 gnd vdd FILL
XFILL_0_DFFPOSX1_449 gnd vdd FILL
XFILL_21_9_1 gnd vdd FILL
XFILL_20_4_0 gnd vdd FILL
XFILL_5_DFFPOSX1_1010 gnd vdd FILL
XFILL_5_DFFPOSX1_1032 gnd vdd FILL
XFILL_5_DFFPOSX1_1021 gnd vdd FILL
XFILL_24_11_1 gnd vdd FILL
XFILL_3_DFFPOSX1_909 gnd vdd FILL
XDFFPOSX1_10 BUFX2_709/A CLKBUF1_41/Y DFFPOSX1_10/D gnd vdd DFFPOSX1
XDFFPOSX1_21 BUFX2_690/A CLKBUF1_95/Y DFFPOSX1_21/D gnd vdd DFFPOSX1
XDFFPOSX1_32 BUFX2_702/A CLKBUF1_101/Y DFFPOSX1_32/D gnd vdd DFFPOSX1
XDFFPOSX1_43 BUFX2_742/A CLKBUF1_93/Y DFFPOSX1_43/D gnd vdd DFFPOSX1
XDFFPOSX1_54 BUFX2_723/A CLKBUF1_78/Y DFFPOSX1_54/D gnd vdd DFFPOSX1
XOAI21X1_1550 BUFX4_139/Y BUFX4_68/Y BUFX2_244/A gnd OAI21X1_1552/C vdd OAI21X1
XDFFPOSX1_76 BUFX2_775/A CLKBUF1_17/Y DFFPOSX1_76/D gnd vdd DFFPOSX1
XOAI21X1_1583 BUFX4_349/Y INVX2_119/Y NAND2X1_652/Y gnd OAI21X1_1583/Y vdd OAI21X1
XOAI21X1_1572 NAND2X1_647/Y BUFX4_297/Y OAI21X1_1572/C gnd OAI21X1_1572/Y vdd OAI21X1
XDFFPOSX1_87 BUFX2_756/A CLKBUF1_19/Y DFFPOSX1_87/D gnd vdd DFFPOSX1
XOAI21X1_1561 BUFX4_141/Y BUFX4_58/Y BUFX2_248/A gnd OAI21X1_1563/C vdd OAI21X1
XDFFPOSX1_65 BUFX2_735/A CLKBUF1_69/Y DFFPOSX1_65/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1770 gnd vdd FILL
XOAI21X1_1594 BUFX4_363/Y INVX2_130/Y NAND2X1_663/Y gnd OAI21X1_1594/Y vdd OAI21X1
XFILL_1_OAI21X1_1792 gnd vdd FILL
XFILL_1_OAI21X1_1781 gnd vdd FILL
XFILL_1_OAI21X1_710 gnd vdd FILL
XFILL_1_OAI21X1_721 gnd vdd FILL
XDFFPOSX1_98 BUFX2_769/A CLKBUF1_6/Y DFFPOSX1_98/D gnd vdd DFFPOSX1
XFILL_0_OAI21X1_583 gnd vdd FILL
XFILL_1_OAI21X1_732 gnd vdd FILL
XFILL_1_OAI21X1_743 gnd vdd FILL
XFILL_0_OAI21X1_550 gnd vdd FILL
XFILL_1_OAI21X1_754 gnd vdd FILL
XFILL_0_OAI21X1_561 gnd vdd FILL
XFILL_0_OAI21X1_572 gnd vdd FILL
XFILL_1_OAI21X1_765 gnd vdd FILL
XFILL_1_OAI21X1_776 gnd vdd FILL
XFILL_1_OAI21X1_787 gnd vdd FILL
XFILL_0_OAI21X1_594 gnd vdd FILL
XFILL_1_OAI21X1_798 gnd vdd FILL
XFILL_28_5_0 gnd vdd FILL
XBUFX2_608 BUFX2_608/A gnd majID4_o[60] vdd BUFX2
XBUFX2_619 BUFX2_619/A gnd majID4_o[59] vdd BUFX2
XFILL_3_5_0 gnd vdd FILL
XFILL_0_CLKBUF1_61 gnd vdd FILL
XFILL_0_CLKBUF1_72 gnd vdd FILL
XFILL_0_CLKBUF1_50 gnd vdd FILL
XFILL_0_CLKBUF1_83 gnd vdd FILL
XFILL_0_CLKBUF1_94 gnd vdd FILL
XFILL_1_NAND2X1_760 gnd vdd FILL
XFILL_0_OAI21X1_1360 gnd vdd FILL
XFILL_29_10_1 gnd vdd FILL
XFILL_0_DFFPOSX1_950 gnd vdd FILL
XFILL_0_OAI21X1_1393 gnd vdd FILL
XFILL_0_DFFPOSX1_961 gnd vdd FILL
XFILL_0_OAI21X1_1382 gnd vdd FILL
XFILL_0_OAI21X1_1371 gnd vdd FILL
XFILL_0_DFFPOSX1_983 gnd vdd FILL
XFILL_0_DFFPOSX1_994 gnd vdd FILL
XFILL_0_DFFPOSX1_972 gnd vdd FILL
XFILL_12_9_1 gnd vdd FILL
XFILL_11_4_0 gnd vdd FILL
XINVX2_104 INVX2_104/A gnd INVX2_104/Y vdd INVX2
XFILL_0_BUFX2_304 gnd vdd FILL
XINVX2_126 bundlePid_i[22] gnd INVX2_126/Y vdd INVX2
XFILL_0_BUFX2_348 gnd vdd FILL
XINVX2_137 bundlePid_i[11] gnd INVX2_137/Y vdd INVX2
XFILL_0_BUFX2_326 gnd vdd FILL
XFILL_0_BUFX2_315 gnd vdd FILL
XINVX2_115 bundlePid_i[1] gnd INVX2_115/Y vdd INVX2
XFILL_0_BUFX2_337 gnd vdd FILL
XFILL_0_BUFX2_359 gnd vdd FILL
XINVX2_148 bundleTid_i[61] gnd INVX2_148/Y vdd INVX2
XINVX2_159 bundleTid_i[50] gnd INVX2_159/Y vdd INVX2
XFILL_2_OAI21X1_1432 gnd vdd FILL
XFILL_2_OAI21X1_1410 gnd vdd FILL
XFILL_19_5_0 gnd vdd FILL
XFILL_4_11_1 gnd vdd FILL
XFILL_2_NOR3X1_10 gnd vdd FILL
XFILL_0_INVX1_2 gnd vdd FILL
XFILL_1_NAND3X1_11 gnd vdd FILL
XFILL_1_OAI21X1_1022 gnd vdd FILL
XFILL_1_NAND3X1_55 gnd vdd FILL
XFILL_1_NAND3X1_33 gnd vdd FILL
XDFFPOSX1_403 BUFX2_435/A CLKBUF1_22/Y OAI21X1_375/Y gnd vdd DFFPOSX1
XFILL_1_NAND3X1_22 gnd vdd FILL
XFILL_1_NAND3X1_44 gnd vdd FILL
XFILL_1_OAI21X1_1000 gnd vdd FILL
XFILL_1_OAI21X1_1011 gnd vdd FILL
XFILL_0_BUFX2_860 gnd vdd FILL
XDFFPOSX1_414 BUFX2_447/A CLKBUF1_11/Y OAI21X1_386/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1033 gnd vdd FILL
XFILL_1_OAI21X1_1044 gnd vdd FILL
XFILL_1_NAND3X1_66 gnd vdd FILL
XFILL_1_OAI21X1_1055 gnd vdd FILL
XFILL_1_DFFPOSX1_601 gnd vdd FILL
XFILL_1_DFFPOSX1_612 gnd vdd FILL
XFILL_1_DFFPOSX1_623 gnd vdd FILL
XDFFPOSX1_447 BUFX2_477/A CLKBUF1_33/Y OAI21X1_441/Y gnd vdd DFFPOSX1
XDFFPOSX1_425 BUFX2_502/A CLKBUF1_66/Y OAI21X1_404/Y gnd vdd DFFPOSX1
XDFFPOSX1_436 BUFX2_465/A CLKBUF1_18/Y OAI21X1_424/Y gnd vdd DFFPOSX1
XINVX1_170 bundle_i[98] gnd INVX1_170/Y vdd INVX1
XFILL_0_BUFX2_893 gnd vdd FILL
XFILL_1_DFFPOSX1_645 gnd vdd FILL
XFILL_1_DFFPOSX1_634 gnd vdd FILL
XFILL_1_DFFPOSX1_656 gnd vdd FILL
XFILL_0_BUFX2_871 gnd vdd FILL
XFILL_1_OAI21X1_1066 gnd vdd FILL
XDFFPOSX1_458 BUFX2_489/A CLKBUF1_29/Y OAI21X1_456/Y gnd vdd DFFPOSX1
XDFFPOSX1_469 BUFX2_501/A CLKBUF1_22/Y OAI21X1_475/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1099 gnd vdd FILL
XFILL_1_OAI21X1_1088 gnd vdd FILL
XFILL_0_BUFX2_882 gnd vdd FILL
XFILL_1_OAI21X1_1077 gnd vdd FILL
XINVX1_192 INVX1_192/A gnd INVX1_192/Y vdd INVX1
XNAND2X1_517 bundleAddress_i[39] XNOR2X1_62/A gnd XNOR2X1_63/A vdd NAND2X1
XINVX1_181 bundleAddress_i[3] gnd INVX1_181/Y vdd INVX1
XFILL_1_DFFPOSX1_678 gnd vdd FILL
XFILL_1_DFFPOSX1_667 gnd vdd FILL
XFILL_1_DFFPOSX1_689 gnd vdd FILL
XNAND2X1_506 BUFX2_78/A BUFX4_192/Y gnd NAND2X1_506/Y vdd NAND2X1
XFILL_6_DFFPOSX1_271 gnd vdd FILL
XNAND2X1_528 bundleAddress_i[33] NOR2X1_146/B gnd NOR2X1_148/B vdd NAND2X1
XNAND2X1_539 bundleAddress_i[27] XNOR2X1_68/A gnd XNOR2X1_69/A vdd NAND2X1
XFILL_6_DFFPOSX1_260 gnd vdd FILL
XFILL_9_10_1 gnd vdd FILL
XFILL_6_DFFPOSX1_282 gnd vdd FILL
XFILL_6_DFFPOSX1_293 gnd vdd FILL
XFILL_0_INVX2_91 gnd vdd FILL
XFILL_0_INVX2_80 gnd vdd FILL
XFILL_0_AND2X2_29 gnd vdd FILL
XFILL_10_17_1 gnd vdd FILL
XFILL_0_AND2X2_18 gnd vdd FILL
XFILL_0_DFFPOSX1_202 gnd vdd FILL
XFILL_0_DFFPOSX1_213 gnd vdd FILL
XFILL_0_DFFPOSX1_246 gnd vdd FILL
XFILL_0_DFFPOSX1_235 gnd vdd FILL
XFILL_0_DFFPOSX1_224 gnd vdd FILL
XFILL_0_DFFPOSX1_257 gnd vdd FILL
XFILL_0_DFFPOSX1_279 gnd vdd FILL
XFILL_0_DFFPOSX1_268 gnd vdd FILL
XFILL_3_DFFPOSX1_728 gnd vdd FILL
XFILL_3_DFFPOSX1_706 gnd vdd FILL
XFILL_3_DFFPOSX1_717 gnd vdd FILL
XFILL_3_CLKBUF1_16 gnd vdd FILL
XFILL_3_CLKBUF1_27 gnd vdd FILL
XFILL_3_CLKBUF1_49 gnd vdd FILL
XFILL_3_DFFPOSX1_739 gnd vdd FILL
XFILL_3_CLKBUF1_38 gnd vdd FILL
XOAI21X1_1391 NOR2X1_123/Y BUFX4_291/Y OAI21X1_1391/C gnd OAI21X1_1391/Y vdd OAI21X1
XOAI21X1_1380 INVX1_217/A INVX1_218/Y BUFX4_310/Y gnd OAI21X1_1381/B vdd OAI21X1
XDFFPOSX1_981 BUFX2_233/A CLKBUF1_30/Y OAI21X1_1521/Y gnd vdd DFFPOSX1
XFILL_1_NOR2X1_112 gnd vdd FILL
XDFFPOSX1_970 BUFX2_221/A CLKBUF1_85/Y OAI21X1_1484/Y gnd vdd DFFPOSX1
XDFFPOSX1_992 BUFX2_245/A CLKBUF1_20/Y OAI21X1_1555/Y gnd vdd DFFPOSX1
XFILL_1_NOR2X1_134 gnd vdd FILL
XFILL_2_OAI21X1_733 gnd vdd FILL
XFILL_0_OAI21X1_380 gnd vdd FILL
XFILL_1_OAI21X1_540 gnd vdd FILL
XFILL_0_OAI21X1_391 gnd vdd FILL
XFILL_1_NOR2X1_156 gnd vdd FILL
XFILL_1_OAI21X1_551 gnd vdd FILL
XFILL_1_OAI21X1_562 gnd vdd FILL
XFILL_1_OAI21X1_584 gnd vdd FILL
XFILL_1_NOR2X1_167 gnd vdd FILL
XFILL_1_OAI21X1_595 gnd vdd FILL
XFILL_1_OAI21X1_573 gnd vdd FILL
XFILL_15_16_1 gnd vdd FILL
XFILL_2_DFFPOSX1_318 gnd vdd FILL
XFILL_2_DFFPOSX1_307 gnd vdd FILL
XFILL_2_DFFPOSX1_329 gnd vdd FILL
XBUFX2_416 BUFX2_416/A gnd majID1_o[60] vdd BUFX2
XBUFX2_405 BUFX2_405/A gnd majID1_o[61] vdd BUFX2
XBUFX2_427 BUFX2_427/A gnd majID1_o[59] vdd BUFX2
XBUFX2_438 BUFX2_438/A gnd majID1_o[58] vdd BUFX2
XBUFX2_449 BUFX2_449/A gnd majID1_o[57] vdd BUFX2
XFILL_1_BUFX4_310 gnd vdd FILL
XFILL_1_BUFX4_321 gnd vdd FILL
XFILL_1_BUFX4_332 gnd vdd FILL
XFILL_1_NAND2X1_590 gnd vdd FILL
XFILL_1_BUFX4_365 gnd vdd FILL
XFILL_0_OAI21X1_1190 gnd vdd FILL
XFILL_1_BUFX4_343 gnd vdd FILL
XFILL_1_BUFX4_354 gnd vdd FILL
XFILL_0_DFFPOSX1_791 gnd vdd FILL
XFILL_1_BUFX4_376 gnd vdd FILL
XFILL_1_BUFX4_387 gnd vdd FILL
XFILL_0_DFFPOSX1_780 gnd vdd FILL
XFILL_2_OAI21X1_45 gnd vdd FILL
XFILL_0_BUFX2_112 gnd vdd FILL
XFILL_2_OAI21X1_67 gnd vdd FILL
XFILL_0_BUFX2_101 gnd vdd FILL
XFILL_0_BUFX2_134 gnd vdd FILL
XFILL_0_BUFX2_156 gnd vdd FILL
XFILL_0_BUFX2_123 gnd vdd FILL
XFILL_0_BUFX2_145 gnd vdd FILL
XFILL_0_BUFX2_167 gnd vdd FILL
XFILL_0_BUFX2_189 gnd vdd FILL
XFILL_0_BUFX2_178 gnd vdd FILL
XFILL_33_17_1 gnd vdd FILL
XFILL_14_11_0 gnd vdd FILL
XFILL_35_8_1 gnd vdd FILL
XFILL_2_DFFPOSX1_841 gnd vdd FILL
XFILL_2_DFFPOSX1_830 gnd vdd FILL
XFILL_2_DFFPOSX1_874 gnd vdd FILL
XBUFX2_961 BUFX2_961/A gnd tid3_o[57] vdd BUFX2
XFILL_34_3_0 gnd vdd FILL
XBUFX2_972 BUFX2_972/A gnd tid4_o[52] vdd BUFX2
XBUFX2_983 BUFX2_983/A gnd tid4_o[42] vdd BUFX2
XFILL_2_DFFPOSX1_852 gnd vdd FILL
XBUFX2_950 BUFX2_950/A gnd tid3_o[58] vdd BUFX2
XFILL_2_DFFPOSX1_863 gnd vdd FILL
XBUFX2_994 BUFX2_994/A gnd tid4_o[32] vdd BUFX2
XFILL_2_DFFPOSX1_885 gnd vdd FILL
XFILL_2_DFFPOSX1_896 gnd vdd FILL
XOAI21X1_308 BUFX4_151/Y BUFX4_43/Y BUFX2_1019/A gnd OAI21X1_309/C vdd OAI21X1
XOAI21X1_319 INVX2_3/Y INVX8_2/A OAI21X1_319/C gnd OAI21X1_319/Y vdd OAI21X1
XDFFPOSX1_211 BUFX2_883/A CLKBUF1_93/Y OAI21X1_55/Y gnd vdd DFFPOSX1
XDFFPOSX1_200 BUFX2_871/A CLKBUF1_16/Y OAI21X1_44/Y gnd vdd DFFPOSX1
XBUFX4_6 BUFX4_6/A gnd BUFX4_6/Y vdd BUFX4
XFILL_2_AOI21X1_3 gnd vdd FILL
XDFFPOSX1_222 BUFX2_895/A CLKBUF1_15/Y OAI21X1_66/Y gnd vdd DFFPOSX1
XDFFPOSX1_255 BUFX2_925/A CLKBUF1_32/Y OAI21X1_127/Y gnd vdd DFFPOSX1
XDFFPOSX1_244 BUFX2_913/A CLKBUF1_47/Y OAI21X1_105/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_431 gnd vdd FILL
XFILL_1_DFFPOSX1_420 gnd vdd FILL
XDFFPOSX1_233 BUFX2_950/A CLKBUF1_37/Y OAI21X1_83/Y gnd vdd DFFPOSX1
XFILL_38_16_1 gnd vdd FILL
XFILL_0_BUFX2_690 gnd vdd FILL
XDFFPOSX1_266 BUFX2_937/A CLKBUF1_8/Y OAI21X1_149/Y gnd vdd DFFPOSX1
XDFFPOSX1_277 BUFX2_949/A CLKBUF1_40/Y OAI21X1_171/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_442 gnd vdd FILL
XFILL_1_DFFPOSX1_453 gnd vdd FILL
XFILL_1_DFFPOSX1_464 gnd vdd FILL
XDFFPOSX1_288 BUFX2_962/A CLKBUF1_2/Y OAI21X1_193/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_475 gnd vdd FILL
XNAND2X1_303 bundleStartMajId_i[6] NOR2X1_97/Y gnd OAI21X1_645/A vdd NAND2X1
XNAND2X1_336 INVX2_38/Y NOR3X1_11/C gnd NAND2X1_337/B vdd NAND2X1
XDFFPOSX1_299 BUFX2_1030/A CLKBUF1_26/Y OAI21X1_215/Y gnd vdd DFFPOSX1
XFILL_19_10_0 gnd vdd FILL
XNAND2X1_325 OAI21X1_748/Y OR2X2_15/Y gnd OAI21X1_750/A vdd NAND2X1
XFILL_1_DFFPOSX1_486 gnd vdd FILL
XFILL_1_DFFPOSX1_497 gnd vdd FILL
XNAND2X1_314 INVX4_6/Y OAI21X1_698/C gnd OAI21X1_701/C vdd NAND2X1
XNAND2X1_358 BUFX4_263/Y bundle_i[11] gnd OAI21X1_864/C vdd NAND2X1
XFILL_4_DFFPOSX1_902 gnd vdd FILL
XNAND2X1_369 BUFX4_268/Y bundle_i[0] gnd OAI21X1_875/C vdd NAND2X1
XNAND2X1_347 BUFX4_262/Y bundle_i[22] gnd OAI21X1_853/C vdd NAND2X1
XFILL_4_DFFPOSX1_913 gnd vdd FILL
XFILL_4_DFFPOSX1_946 gnd vdd FILL
XNOR3X1_10 NOR3X1_4/A INVX1_44/Y NOR3X1_8/C gnd NOR3X1_10/Y vdd NOR3X1
XFILL_4_DFFPOSX1_935 gnd vdd FILL
XFILL_4_DFFPOSX1_924 gnd vdd FILL
XFILL_32_12_0 gnd vdd FILL
XFILL_4_DFFPOSX1_968 gnd vdd FILL
XFILL_4_DFFPOSX1_979 gnd vdd FILL
XFILL_4_DFFPOSX1_957 gnd vdd FILL
XFILL_26_8_1 gnd vdd FILL
XFILL_25_3_0 gnd vdd FILL
XFILL_1_8_1 gnd vdd FILL
XFILL_0_3_0 gnd vdd FILL
XFILL_1_INVX2_36 gnd vdd FILL
XFILL_1_BUFX2_803 gnd vdd FILL
XFILL_0_XNOR2X1_2 gnd vdd FILL
XFILL_1_BUFX2_814 gnd vdd FILL
XFILL_1_BUFX2_825 gnd vdd FILL
XINVX4_6 bundleStartMajId_i[48] gnd INVX4_6/Y vdd INVX4
XFILL_1_BUFX2_869 gnd vdd FILL
XFILL_1_BUFX2_847 gnd vdd FILL
XFILL_1_BUFX2_858 gnd vdd FILL
XOAI21X1_831 BUFX4_171/Y BUFX4_77/Y BUFX2_640/A gnd OAI21X1_832/C vdd OAI21X1
XOAI21X1_842 NOR3X1_11/Y bundleStartMajId_i[0] BUFX4_288/Y gnd OAI21X1_843/A vdd OAI21X1
XFILL_3_DFFPOSX1_503 gnd vdd FILL
XOAI21X1_820 NAND3X1_33/Y INVX2_46/Y INVX2_36/Y gnd OAI21X1_820/Y vdd OAI21X1
XOAI21X1_864 INVX1_65/Y BUFX4_263/Y OAI21X1_864/C gnd OAI21X1_864/Y vdd OAI21X1
XFILL_3_DFFPOSX1_547 gnd vdd FILL
XFILL_3_DFFPOSX1_525 gnd vdd FILL
XFILL_3_DFFPOSX1_536 gnd vdd FILL
XFILL_3_DFFPOSX1_514 gnd vdd FILL
XOAI21X1_875 INVX1_76/Y BUFX4_268/Y OAI21X1_875/C gnd OAI21X1_875/Y vdd OAI21X1
XOAI21X1_853 INVX1_54/Y INVX8_4/A OAI21X1_853/C gnd OAI21X1_853/Y vdd OAI21X1
XFILL_3_DFFPOSX1_569 gnd vdd FILL
XOAI21X1_897 INVX1_98/Y BUFX4_189/Y OAI21X1_897/C gnd OAI21X1_897/Y vdd OAI21X1
XOAI21X1_886 INVX1_87/Y BUFX4_186/Y OAI21X1_886/C gnd OAI21X1_886/Y vdd OAI21X1
XFILL_3_DFFPOSX1_558 gnd vdd FILL
XFILL_37_11_0 gnd vdd FILL
XFILL_8_4_0 gnd vdd FILL
XFILL_9_9_1 gnd vdd FILL
XFILL_1_OAI21X1_370 gnd vdd FILL
XFILL_1_OAI21X1_381 gnd vdd FILL
XFILL_1_OAI21X1_392 gnd vdd FILL
XFILL_2_OAI21X1_563 gnd vdd FILL
XFILL_1_CLKBUF1_2 gnd vdd FILL
XBUFX2_202 BUFX2_202/A gnd addr4_o[46] vdd BUFX2
XFILL_2_DFFPOSX1_104 gnd vdd FILL
XFILL_2_DFFPOSX1_126 gnd vdd FILL
XFILL_2_DFFPOSX1_115 gnd vdd FILL
XFILL_2_DFFPOSX1_137 gnd vdd FILL
XBUFX2_213 BUFX2_213/A gnd addr4_o[36] vdd BUFX2
XFILL_0_NAND3X1_63 gnd vdd FILL
XFILL_0_NAND3X1_52 gnd vdd FILL
XBUFX2_235 BUFX2_235/A gnd addr4_o[16] vdd BUFX2
XFILL_0_NAND3X1_41 gnd vdd FILL
XFILL_0_NAND3X1_30 gnd vdd FILL
XBUFX2_224 BUFX2_224/A gnd addr4_o[26] vdd BUFX2
XFILL_2_DFFPOSX1_148 gnd vdd FILL
XFILL_17_8_1 gnd vdd FILL
XFILL_16_3_0 gnd vdd FILL
XBUFX2_268 INVX1_60/A gnd instr1_o[16] vdd BUFX2
XBUFX2_257 BUFX2_257/A gnd enable1_o vdd BUFX2
XFILL_2_DFFPOSX1_159 gnd vdd FILL
XBUFX2_246 INVX1_227/A gnd addr4_o[6] vdd BUFX2
XBUFX2_279 INVX1_70/A gnd instr1_o[6] vdd BUFX2
XFILL_5_DFFPOSX1_608 gnd vdd FILL
XFILL_5_DFFPOSX1_619 gnd vdd FILL
XFILL_1_BUFX4_140 gnd vdd FILL
XFILL_1_BUFX4_151 gnd vdd FILL
XFILL_1_BUFX4_162 gnd vdd FILL
XFILL_1_BUFX4_173 gnd vdd FILL
XFILL_1_BUFX4_184 gnd vdd FILL
XFILL_1_BUFX4_195 gnd vdd FILL
XFILL_2_OAI21X1_6 gnd vdd FILL
XFILL_4_DFFPOSX1_209 gnd vdd FILL
XNAND3X1_9 bundleStartMajId_i[18] bundleStartMajId_i[17] bundleStartMajId_i[16] gnd
+ NOR3X1_3/C vdd NAND3X1
XFILL_2_CLKBUF1_13 gnd vdd FILL
XFILL_2_CLKBUF1_57 gnd vdd FILL
XFILL_2_CLKBUF1_35 gnd vdd FILL
XFILL_2_CLKBUF1_24 gnd vdd FILL
XFILL_2_CLKBUF1_46 gnd vdd FILL
XFILL_2_CLKBUF1_68 gnd vdd FILL
XFILL_2_OAI21X1_1070 gnd vdd FILL
XFILL_2_CLKBUF1_79 gnd vdd FILL
XFILL_2_OAI21X1_1092 gnd vdd FILL
XBUFX2_780 BUFX2_780/A gnd tid1_o[52] vdd BUFX2
XBUFX2_791 BUFX2_791/A gnd tid1_o[42] vdd BUFX2
XFILL_2_DFFPOSX1_660 gnd vdd FILL
XFILL_2_DFFPOSX1_693 gnd vdd FILL
XFILL_2_DFFPOSX1_671 gnd vdd FILL
XFILL_2_DFFPOSX1_682 gnd vdd FILL
XFILL_0_NOR2X1_131 gnd vdd FILL
XFILL_0_NOR2X1_120 gnd vdd FILL
XFILL_0_NOR2X1_164 gnd vdd FILL
XFILL_0_NOR2X1_142 gnd vdd FILL
XFILL_0_NOR2X1_153 gnd vdd FILL
XOAI21X1_138 BUFX4_100/Y BUFX4_329/Y BUFX2_932/A gnd OAI21X1_139/C vdd OAI21X1
XOAI21X1_127 BUFX4_123/Y INVX2_173/Y OAI21X1_127/C gnd OAI21X1_127/Y vdd OAI21X1
XOAI21X1_105 BUFX4_147/Y INVX2_162/Y OAI21X1_105/C gnd OAI21X1_105/Y vdd OAI21X1
XOAI21X1_116 BUFX4_1/Y BUFX4_348/Y BUFX2_920/A gnd OAI21X1_117/C vdd OAI21X1
XFILL_0_NOR2X1_175 gnd vdd FILL
XFILL_0_NOR2X1_197 gnd vdd FILL
XFILL_0_NOR2X1_186 gnd vdd FILL
XFILL_0_DFFPOSX1_1027 gnd vdd FILL
XFILL_0_DFFPOSX1_1005 gnd vdd FILL
XOAI21X1_149 BUFX4_137/Y INVX2_184/Y OAI21X1_149/C gnd OAI21X1_149/Y vdd OAI21X1
XFILL_0_DFFPOSX1_1016 gnd vdd FILL
XBUFX2_3 BUFX2_3/A gnd addr1_o[53] vdd BUFX2
XFILL_1_DFFPOSX1_250 gnd vdd FILL
XFILL_1_DFFPOSX1_261 gnd vdd FILL
XFILL_1_DFFPOSX1_272 gnd vdd FILL
XFILL_1_DFFPOSX1_283 gnd vdd FILL
XNAND2X1_100 BUFX2_414/A OAI21X1_2/A gnd OAI21X1_356/C vdd NAND2X1
XNAND2X1_122 BUFX2_439/A BUFX4_323/Y gnd OAI21X1_378/C vdd NAND2X1
XNAND2X1_111 BUFX2_426/A BUFX4_325/Y gnd OAI21X1_367/C vdd NAND2X1
XFILL_1_DFFPOSX1_294 gnd vdd FILL
XNAND2X1_144 BUFX2_491/A BUFX4_199/Y gnd OAI21X1_401/C vdd NAND2X1
XNAND2X1_133 BUFX2_451/A BUFX4_337/Y gnd OAI21X1_389/C vdd NAND2X1
XFILL_4_DFFPOSX1_710 gnd vdd FILL
XFILL_4_DFFPOSX1_721 gnd vdd FILL
XNAND2X1_155 bundleStartMajId_i[54] bundleStartMajId_i[53] gnd OR2X2_1/A vdd NAND2X1
XNAND2X1_166 bundleStartMajId_i[50] bundleStartMajId_i[49] gnd NOR2X1_10/B vdd NAND2X1
XNAND2X1_177 INVX2_20/Y NAND2X1_177/B gnd OAI21X1_430/C vdd NAND2X1
XFILL_1_OAI21X1_42 gnd vdd FILL
XFILL_1_OAI21X1_20 gnd vdd FILL
XFILL_4_DFFPOSX1_754 gnd vdd FILL
XFILL_1_OAI21X1_31 gnd vdd FILL
XFILL_4_DFFPOSX1_743 gnd vdd FILL
XNAND2X1_199 bundleStartMajId_i[39] bundleStartMajId_i[36] gnd OR2X2_4/B vdd NAND2X1
XFILL_4_DFFPOSX1_732 gnd vdd FILL
XNAND2X1_188 BUFX2_474/A BUFX4_214/Y gnd OAI21X1_436/C vdd NAND2X1
XFILL_4_DFFPOSX1_765 gnd vdd FILL
XFILL_1_OAI21X1_64 gnd vdd FILL
XFILL_1_OAI21X1_53 gnd vdd FILL
XFILL_4_DFFPOSX1_776 gnd vdd FILL
XFILL_1_OAI21X1_75 gnd vdd FILL
XFILL_4_DFFPOSX1_787 gnd vdd FILL
XFILL_1_OAI21X1_86 gnd vdd FILL
XFILL_4_DFFPOSX1_798 gnd vdd FILL
XFILL_1_OAI21X1_97 gnd vdd FILL
XFILL_0_DFFPOSX1_7 gnd vdd FILL
XFILL_1_BUFX2_611 gnd vdd FILL
XFILL_1_BUFX2_600 gnd vdd FILL
XFILL_1_BUFX2_655 gnd vdd FILL
XFILL_1_BUFX2_622 gnd vdd FILL
XINVX2_3 bundleTid_i[4] gnd INVX2_3/Y vdd INVX2
XFILL_0_BUFX4_207 gnd vdd FILL
XFILL_3_DFFPOSX1_322 gnd vdd FILL
XFILL_0_BUFX4_218 gnd vdd FILL
XFILL_0_BUFX4_229 gnd vdd FILL
XOAI21X1_650 BUFX4_3/A BUFX4_356/Y BUFX2_578/A gnd OAI21X1_651/C vdd OAI21X1
XFILL_3_DFFPOSX1_311 gnd vdd FILL
XFILL_23_17_0 gnd vdd FILL
XFILL_3_DFFPOSX1_300 gnd vdd FILL
XFILL_1_BUFX2_666 gnd vdd FILL
XFILL_3_DFFPOSX1_333 gnd vdd FILL
XFILL_1_BUFX2_699 gnd vdd FILL
XAOI21X1_3 INVX2_46/A INVX1_20/Y bundleStartMajId_i[8] gnd AOI21X1_3/Y vdd AOI21X1
XFILL_3_DFFPOSX1_355 gnd vdd FILL
XOAI21X1_683 OAI21X1_683/A BUFX4_299/Y OAI21X1_683/C gnd OAI21X1_683/Y vdd OAI21X1
XFILL_3_DFFPOSX1_344 gnd vdd FILL
XOAI21X1_672 INVX2_52/Y INVX2_11/Y INVX2_12/Y gnd OAI21X1_673/C vdd OAI21X1
XOAI21X1_661 BUFX4_299/Y NOR2X1_2/Y OAI21X1_661/C gnd OAI21X1_661/Y vdd OAI21X1
XFILL_3_DFFPOSX1_388 gnd vdd FILL
XOAI21X1_694 BUFX4_122/Y BUFX4_76/Y BUFX2_589/A gnd OAI21X1_695/C vdd OAI21X1
XFILL_3_DFFPOSX1_377 gnd vdd FILL
XFILL_3_DFFPOSX1_366 gnd vdd FILL
XFILL_3_DFFPOSX1_399 gnd vdd FILL
XFILL_6_DFFPOSX1_815 gnd vdd FILL
XFILL_0_INVX4_26 gnd vdd FILL
XFILL_6_DFFPOSX1_837 gnd vdd FILL
XFILL_6_DFFPOSX1_804 gnd vdd FILL
XFILL_6_DFFPOSX1_826 gnd vdd FILL
XFILL_0_INVX4_15 gnd vdd FILL
XFILL_0_INVX4_37 gnd vdd FILL
XFILL_0_INVX4_48 gnd vdd FILL
XXNOR2X1_22 INVX1_20/A INVX4_24/Y gnd XNOR2X1_22/Y vdd XNOR2X1
XFILL_6_DFFPOSX1_848 gnd vdd FILL
XFILL_3_DFFPOSX1_1009 gnd vdd FILL
XXNOR2X1_11 XNOR2X1_11/A INVX4_14/Y gnd XNOR2X1_11/Y vdd XNOR2X1
XXNOR2X1_66 XNOR2X1_66/A INVX4_38/Y gnd XNOR2X1_66/Y vdd XNOR2X1
XXNOR2X1_55 XNOR2X1_55/A INVX4_25/Y gnd XNOR2X1_55/Y vdd XNOR2X1
XXNOR2X1_33 NOR2X1_72/Y bundleStartMajId_i[34] gnd XNOR2X1_33/Y vdd XNOR2X1
XXNOR2X1_44 INVX1_37/A INVX4_8/Y gnd XNOR2X1_44/Y vdd XNOR2X1
XXNOR2X1_77 INVX1_200/A bundleAddress_i[48] gnd XNOR2X1_77/Y vdd XNOR2X1
XFILL_1_INVX2_184 gnd vdd FILL
XXNOR2X1_99 XNOR2X1_99/A INVX4_39/Y gnd XNOR2X1_99/Y vdd XNOR2X1
XFILL_2_OAI21X1_371 gnd vdd FILL
XXNOR2X1_88 XNOR2X1_88/A bundleAddress_i[4] gnd XNOR2X1_88/Y vdd XNOR2X1
XBUFX2_10 BUFX2_10/A gnd addr1_o[46] vdd BUFX2
XFILL_0_NAND2X1_407 gnd vdd FILL
XINVX1_90 bundle_i[50] gnd INVX1_90/Y vdd INVX1
XBUFX2_21 BUFX2_21/A gnd addr1_o[36] vdd BUFX2
XFILL_0_NAND2X1_418 gnd vdd FILL
XFILL_0_NAND2X1_429 gnd vdd FILL
XBUFX2_43 BUFX2_43/A gnd addr1_o[16] vdd BUFX2
XBUFX2_54 BUFX2_54/A gnd addr1_o[6] vdd BUFX2
XBUFX2_32 BUFX2_32/A gnd addr1_o[26] vdd BUFX2
XBUFX2_65 BUFX2_65/A gnd addr2_o[63] vdd BUFX2
XBUFX2_87 BUFX2_87/A gnd addr2_o[34] vdd BUFX2
XBUFX2_76 BUFX2_76/A gnd addr2_o[44] vdd BUFX2
XFILL_32_6_1 gnd vdd FILL
XBUFX2_98 BUFX2_98/A gnd addr2_o[24] vdd BUFX2
XFILL_31_1_0 gnd vdd FILL
XFILL_28_16_0 gnd vdd FILL
XFILL_5_DFFPOSX1_416 gnd vdd FILL
XFILL_5_DFFPOSX1_405 gnd vdd FILL
XFILL_5_DFFPOSX1_427 gnd vdd FILL
XFILL_1_BUFX4_10 gnd vdd FILL
XFILL_5_DFFPOSX1_449 gnd vdd FILL
XFILL_5_DFFPOSX1_438 gnd vdd FILL
XFILL_1_BUFX4_43 gnd vdd FILL
XFILL_1_BUFX4_32 gnd vdd FILL
XFILL_1_BUFX4_54 gnd vdd FILL
XFILL_1_BUFX4_21 gnd vdd FILL
XFILL_1_BUFX4_65 gnd vdd FILL
XFILL_1_BUFX4_87 gnd vdd FILL
XFILL_1_BUFX4_76 gnd vdd FILL
XFILL_1_BUFX4_98 gnd vdd FILL
XFILL_0_OAI21X1_924 gnd vdd FILL
XNOR2X1_1 bundleStartMajId_i[63] bundleStartMajId_i[62] gnd NOR2X1_2/A vdd NOR2X1
XFILL_0_OAI21X1_902 gnd vdd FILL
XFILL_0_OAI21X1_913 gnd vdd FILL
XFILL_0_OAI21X1_957 gnd vdd FILL
XFILL_0_OAI21X1_935 gnd vdd FILL
XFILL_0_OAI21X1_946 gnd vdd FILL
XFILL_0_OAI21X1_979 gnd vdd FILL
XFILL_0_OAI21X1_968 gnd vdd FILL
XFILL_2_BUFX4_105 gnd vdd FILL
XFILL_3_17_0 gnd vdd FILL
XFILL_0_OAI21X1_1701 gnd vdd FILL
XFILL_1_OR2X2_13 gnd vdd FILL
XFILL_0_OAI21X1_1712 gnd vdd FILL
XFILL_0_OAI21X1_1734 gnd vdd FILL
XFILL_0_OAI21X1_1723 gnd vdd FILL
XFILL_0_OAI21X1_1756 gnd vdd FILL
XFILL_0_OAI21X1_1745 gnd vdd FILL
XFILL_0_OAI21X1_1767 gnd vdd FILL
XFILL_23_6_1 gnd vdd FILL
XFILL_2_DFFPOSX1_490 gnd vdd FILL
XFILL_0_OAI21X1_1778 gnd vdd FILL
XFILL_0_OAI21X1_1789 gnd vdd FILL
XFILL_22_1_0 gnd vdd FILL
XFILL_5_DFFPOSX1_950 gnd vdd FILL
XFILL_5_DFFPOSX1_961 gnd vdd FILL
XFILL_5_DFFPOSX1_983 gnd vdd FILL
XFILL_5_DFFPOSX1_972 gnd vdd FILL
XAOI21X1_22 bundleStartMajId_i[7] OR2X2_12/A BUFX4_155/Y gnd AOI21X1_23/A vdd AOI21X1
XFILL_5_DFFPOSX1_994 gnd vdd FILL
XAOI21X1_44 bundleAddress_i[4] NOR2X1_174/B bundleAddress_i[3] gnd AOI21X1_44/Y vdd
+ AOI21X1
XAOI21X1_11 bundleStartMajId_i[23] NAND3X1_20/Y BUFX4_155/Y gnd AOI21X1_12/A vdd AOI21X1
XAOI21X1_33 bundleStartMajId_i[33] INVX1_40/Y INVX2_24/Y gnd AOI21X1_33/Y vdd AOI21X1
XFILL_0_NOR2X1_29 gnd vdd FILL
XFILL_0_NOR2X1_18 gnd vdd FILL
XAOI21X1_66 INVX1_199/A INVX2_112/Y bundleAddress_i[2] gnd AOI21X1_66/Y vdd AOI21X1
XAOI21X1_55 bundleAddress_i[12] NOR3X1_18/Y bundleAddress_i[11] gnd AOI21X1_55/Y vdd
+ AOI21X1
XOAI21X1_6 OAI21X1_6/A INVX2_6/Y OAI21X1_6/C gnd OAI21X1_6/Y vdd OAI21X1
XFILL_8_16_0 gnd vdd FILL
XXNOR2X1_103 OR2X2_21/A INVX4_44/Y gnd XNOR2X1_103/Y vdd XNOR2X1
XBUFX4_319 BUFX4_385/A gnd BUFX4_319/Y vdd BUFX4
XFILL_4_DFFPOSX1_540 gnd vdd FILL
XBUFX4_308 BUFX4_310/A gnd BUFX4_308/Y vdd BUFX4
XFILL_5_2_0 gnd vdd FILL
XFILL_6_7_1 gnd vdd FILL
XFILL_2_OAI21X1_1817 gnd vdd FILL
XFILL_4_DFFPOSX1_551 gnd vdd FILL
XFILL_4_DFFPOSX1_573 gnd vdd FILL
XFILL_4_DFFPOSX1_562 gnd vdd FILL
XFILL_4_DFFPOSX1_595 gnd vdd FILL
XFILL_4_DFFPOSX1_584 gnd vdd FILL
XFILL_12_14_1 gnd vdd FILL
XFILL_1_BUFX2_1020 gnd vdd FILL
XFILL_14_6_1 gnd vdd FILL
XFILL_13_1_0 gnd vdd FILL
XFILL_1_BUFX2_452 gnd vdd FILL
XFILL_1_BUFX2_463 gnd vdd FILL
XFILL_3_DFFPOSX1_130 gnd vdd FILL
XOAI21X1_1209 BUFX4_148/Y INVX2_54/Y OAI21X1_1209/C gnd OAI21X1_1209/Y vdd OAI21X1
XFILL_1_CLKBUF1_21 gnd vdd FILL
XFILL_1_CLKBUF1_10 gnd vdd FILL
XFILL_1_BUFX2_474 gnd vdd FILL
XFILL_1_BUFX2_496 gnd vdd FILL
XFILL_1_CLKBUF1_65 gnd vdd FILL
XFILL_1_INVX8_5 gnd vdd FILL
XFILL_1_CLKBUF1_32 gnd vdd FILL
XFILL_1_OAI21X1_1418 gnd vdd FILL
XFILL_1_CLKBUF1_43 gnd vdd FILL
XFILL_1_OAI21X1_1407 gnd vdd FILL
XFILL_1_OAI21X1_1429 gnd vdd FILL
XOAI21X1_491 INVX1_22/A NOR2X1_99/B BUFX4_240/Y gnd OAI21X1_492/B vdd OAI21X1
XFILL_3_DFFPOSX1_163 gnd vdd FILL
XFILL_3_DFFPOSX1_152 gnd vdd FILL
XFILL_1_CLKBUF1_54 gnd vdd FILL
XFILL_3_DFFPOSX1_141 gnd vdd FILL
XOAI21X1_480 INVX1_20/Y OAI21X1_480/B OAI21X1_480/C gnd OAI21X1_480/Y vdd OAI21X1
XFILL_0_OAI21X1_209 gnd vdd FILL
XFILL_1_CLKBUF1_98 gnd vdd FILL
XFILL_3_DFFPOSX1_185 gnd vdd FILL
XFILL_1_CLKBUF1_87 gnd vdd FILL
XFILL_3_DFFPOSX1_196 gnd vdd FILL
XFILL_3_DFFPOSX1_174 gnd vdd FILL
XFILL_1_CLKBUF1_76 gnd vdd FILL
XFILL_6_DFFPOSX1_601 gnd vdd FILL
XFILL_17_13_1 gnd vdd FILL
XFILL_6_DFFPOSX1_689 gnd vdd FILL
XFILL_30_15_1 gnd vdd FILL
XFILL_0_NAND2X1_215 gnd vdd FILL
XFILL_0_NAND2X1_204 gnd vdd FILL
XFILL_1_NAND2X1_419 gnd vdd FILL
XFILL_0_NAND2X1_237 gnd vdd FILL
XFILL_0_OAI21X1_1019 gnd vdd FILL
XFILL_0_NAND2X1_259 gnd vdd FILL
XFILL_0_NAND2X1_226 gnd vdd FILL
XFILL_0_OAI21X1_1008 gnd vdd FILL
XFILL_0_NAND2X1_248 gnd vdd FILL
XFILL_0_DFFPOSX1_609 gnd vdd FILL
XFILL_5_DFFPOSX1_202 gnd vdd FILL
XFILL_5_DFFPOSX1_213 gnd vdd FILL
XFILL_5_DFFPOSX1_235 gnd vdd FILL
XFILL_5_DFFPOSX1_224 gnd vdd FILL
XFILL_5_DFFPOSX1_246 gnd vdd FILL
XFILL_5_DFFPOSX1_268 gnd vdd FILL
XFILL_5_DFFPOSX1_257 gnd vdd FILL
XFILL_5_DFFPOSX1_279 gnd vdd FILL
XFILL_0_OAI21X1_50 gnd vdd FILL
XOAI21X1_1710 BUFX4_165/Y BUFX4_34/Y BUFX2_745/A gnd OAI21X1_1711/C vdd OAI21X1
XFILL_0_OAI21X1_61 gnd vdd FILL
XFILL_0_OAI21X1_72 gnd vdd FILL
XOAI21X1_1732 BUFX4_151/Y BUFX4_49/Y BUFX2_748/A gnd OAI21X1_1733/C vdd OAI21X1
XFILL_0_OAI21X1_83 gnd vdd FILL
XOAI21X1_1721 INVX2_122/Y BUFX4_303/Y OAI21X1_1721/C gnd DFFPOSX1_73/D vdd OAI21X1
XOAI21X1_1743 INVX2_133/Y BUFX4_290/Y OAI21X1_1743/C gnd DFFPOSX1_84/D vdd OAI21X1
XFILL_0_OAI21X1_94 gnd vdd FILL
XOAI21X1_1754 BUFX4_159/Y BUFX4_65/Y BUFX2_760/A gnd OAI21X1_1755/C vdd OAI21X1
XOAI21X1_1765 INVX2_144/Y BUFX4_291/Y OAI21X1_1765/C gnd DFFPOSX1_95/D vdd OAI21X1
XOAI21X1_1798 BUFX4_361/Y INVX2_170/Y NAND2X1_739/Y gnd OAI21X1_1798/Y vdd OAI21X1
XFILL_0_OAI21X1_710 gnd vdd FILL
XFILL_0_OAI21X1_732 gnd vdd FILL
XFILL_0_OAI21X1_721 gnd vdd FILL
XFILL_1_OAI21X1_903 gnd vdd FILL
XOAI21X1_1776 BUFX4_337/Y INVX2_148/Y NAND2X1_717/Y gnd OAI21X1_1776/Y vdd OAI21X1
XOAI21X1_1787 BUFX4_320/Y INVX2_159/Y NAND2X1_728/Y gnd OAI21X1_1787/Y vdd OAI21X1
XFILL_1_OAI21X1_914 gnd vdd FILL
XFILL_1_OAI21X1_936 gnd vdd FILL
XFILL_1_OAI21X1_925 gnd vdd FILL
XFILL_0_OAI21X1_765 gnd vdd FILL
XFILL_0_OAI21X1_743 gnd vdd FILL
XFILL_0_OAI21X1_754 gnd vdd FILL
XFILL_1_OAI21X1_969 gnd vdd FILL
XFILL_0_OAI21X1_798 gnd vdd FILL
XFILL_0_OAI21X1_776 gnd vdd FILL
XFILL_0_OAI21X1_787 gnd vdd FILL
XFILL_1_OAI21X1_958 gnd vdd FILL
XFILL_1_OAI21X1_947 gnd vdd FILL
XFILL_35_14_1 gnd vdd FILL
XFILL_2_NAND3X1_15 gnd vdd FILL
XFILL_0_NAND2X1_760 gnd vdd FILL
XFILL_0_NAND2X1_771 gnd vdd FILL
XFILL_0_OAI21X1_1520 gnd vdd FILL
XFILL_0_OAI21X1_1531 gnd vdd FILL
XFILL_0_OAI21X1_1542 gnd vdd FILL
XFILL_0_OAI21X1_1575 gnd vdd FILL
XFILL_0_OAI21X1_1564 gnd vdd FILL
XFILL_0_OAI21X1_1553 gnd vdd FILL
XFILL_0_OAI21X1_1597 gnd vdd FILL
XFILL_0_OAI21X1_1586 gnd vdd FILL
XFILL_5_DFFPOSX1_791 gnd vdd FILL
XFILL_5_DFFPOSX1_780 gnd vdd FILL
XFILL_0_BUFX2_519 gnd vdd FILL
XFILL_0_BUFX2_508 gnd vdd FILL
XBUFX4_127 BUFX4_19/Y gnd BUFX4_127/Y vdd BUFX4
XBUFX4_116 INVX8_4/Y gnd BUFX4_386/A vdd BUFX4
XBUFX4_105 BUFX4_1/A gnd BUFX4_105/Y vdd BUFX4
XFILL_0_INVX1_16 gnd vdd FILL
XFILL_2_OAI21X1_1647 gnd vdd FILL
XBUFX4_149 BUFX4_19/Y gnd BUFX4_149/Y vdd BUFX4
XFILL_2_OAI21X1_1625 gnd vdd FILL
XBUFX4_138 BUFX4_15/Y gnd BUFX4_138/Y vdd BUFX4
XFILL_4_DFFPOSX1_381 gnd vdd FILL
XFILL_0_INVX1_27 gnd vdd FILL
XFILL_0_INVX1_38 gnd vdd FILL
XFILL_1_AND2X2_8 gnd vdd FILL
XFILL_0_INVX1_49 gnd vdd FILL
XFILL_4_DFFPOSX1_370 gnd vdd FILL
XFILL_4_DFFPOSX1_392 gnd vdd FILL
XNOR2X1_209 bundleAddress_i[8] INVX1_215/Y gnd NOR2X1_209/Y vdd NOR2X1
XFILL_1_BUFX2_271 gnd vdd FILL
XFILL_1_BUFX2_260 gnd vdd FILL
XOAI21X1_1028 BUFX4_164/Y BUFX4_64/Y BUFX2_378/A gnd OAI21X1_1029/C vdd OAI21X1
XOAI21X1_1006 BUFX4_151/Y BUFX4_49/Y BUFX2_366/A gnd OAI21X1_1007/C vdd OAI21X1
XFILL_1_OAI21X1_1204 gnd vdd FILL
XOAI21X1_1017 BUFX4_295/Y INVX1_163/Y OAI21X1_1017/C gnd OAI21X1_1017/Y vdd OAI21X1
XFILL_1_OAI21X1_1215 gnd vdd FILL
XFILL_1_OAI21X1_1237 gnd vdd FILL
XOAI21X1_1039 BUFX4_312/Y INVX2_56/Y NAND2X1_405/Y gnd OAI21X1_1039/Y vdd OAI21X1
XFILL_1_OAI21X1_1226 gnd vdd FILL
XFILL_1_OAI21X1_1248 gnd vdd FILL
XDFFPOSX1_607 BUFX2_640/A CLKBUF1_19/Y OAI21X1_832/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_805 gnd vdd FILL
XDFFPOSX1_629 INVX1_58/A CLKBUF1_82/Y OAI21X1_857/Y gnd vdd DFFPOSX1
XDFFPOSX1_618 INVX1_47/A CLKBUF1_81/Y OAI21X1_846/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_816 gnd vdd FILL
XFILL_1_OAI21X1_1259 gnd vdd FILL
XFILL_1_DFFPOSX1_838 gnd vdd FILL
XFILL_1_DFFPOSX1_849 gnd vdd FILL
XFILL_1_DFFPOSX1_827 gnd vdd FILL
XFILL_6_DFFPOSX1_442 gnd vdd FILL
XFILL_6_DFFPOSX1_453 gnd vdd FILL
XFILL_6_DFFPOSX1_486 gnd vdd FILL
XFILL_6_DFFPOSX1_464 gnd vdd FILL
XFILL_6_DFFPOSX1_475 gnd vdd FILL
XFILL_6_DFFPOSX1_497 gnd vdd FILL
XFILL_37_5_1 gnd vdd FILL
XFILL_36_0_0 gnd vdd FILL
XFILL_0_DFFPOSX1_406 gnd vdd FILL
XFILL_1_NAND2X1_238 gnd vdd FILL
XFILL_1_NAND2X1_216 gnd vdd FILL
XFILL_1_NAND3X1_1 gnd vdd FILL
XFILL_0_DFFPOSX1_439 gnd vdd FILL
XFILL_0_DFFPOSX1_428 gnd vdd FILL
XFILL_0_DFFPOSX1_417 gnd vdd FILL
XFILL_5_DFFPOSX1_1000 gnd vdd FILL
XFILL_20_4_1 gnd vdd FILL
XFILL_5_DFFPOSX1_1011 gnd vdd FILL
XFILL_5_DFFPOSX1_1022 gnd vdd FILL
XDFFPOSX1_11 BUFX2_710/A CLKBUF1_93/Y DFFPOSX1_11/D gnd vdd DFFPOSX1
XDFFPOSX1_44 BUFX2_743/A CLKBUF1_42/Y DFFPOSX1_44/D gnd vdd DFFPOSX1
XDFFPOSX1_22 BUFX2_691/A CLKBUF1_73/Y DFFPOSX1_22/D gnd vdd DFFPOSX1
XOAI21X1_1540 BUFX4_160/Y BUFX4_80/Y BUFX2_241/A gnd OAI21X1_1542/C vdd OAI21X1
XDFFPOSX1_33 BUFX2_703/A CLKBUF1_38/Y DFFPOSX1_33/D gnd vdd DFFPOSX1
XDFFPOSX1_77 BUFX2_776/A CLKBUF1_95/Y DFFPOSX1_77/D gnd vdd DFFPOSX1
XOAI21X1_1584 BUFX4_311/Y INVX2_120/Y NAND2X1_653/Y gnd OAI21X1_1584/Y vdd OAI21X1
XOAI21X1_1573 BUFX4_162/Y BUFX4_39/Y BUFX2_253/A gnd OAI21X1_1574/C vdd OAI21X1
XFILL_1_OAI21X1_1760 gnd vdd FILL
XDFFPOSX1_55 BUFX2_724/A CLKBUF1_45/Y DFFPOSX1_55/D gnd vdd DFFPOSX1
XOAI21X1_1562 INVX2_112/A INVX2_90/Y BUFX4_284/Y gnd OAI21X1_1563/B vdd OAI21X1
XOAI21X1_1551 INVX1_226/A INVX4_45/Y BUFX4_286/Y gnd OAI21X1_1552/B vdd OAI21X1
XDFFPOSX1_66 BUFX2_737/A CLKBUF1_75/Y DFFPOSX1_66/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1793 gnd vdd FILL
XOAI21X1_1595 BUFX4_313/Y INVX2_131/Y NAND2X1_664/Y gnd OAI21X1_1595/Y vdd OAI21X1
XFILL_1_OAI21X1_711 gnd vdd FILL
XDFFPOSX1_88 BUFX2_758/A CLKBUF1_40/Y DFFPOSX1_88/D gnd vdd DFFPOSX1
XFILL_0_OAI21X1_540 gnd vdd FILL
XFILL_1_OAI21X1_1782 gnd vdd FILL
XFILL_1_OAI21X1_1771 gnd vdd FILL
XDFFPOSX1_99 BUFX2_770/A CLKBUF1_66/Y DFFPOSX1_99/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_700 gnd vdd FILL
XFILL_1_OAI21X1_744 gnd vdd FILL
XFILL_1_OAI21X1_733 gnd vdd FILL
XFILL_1_OAI21X1_755 gnd vdd FILL
XFILL_1_OAI21X1_722 gnd vdd FILL
XFILL_0_OAI21X1_551 gnd vdd FILL
XFILL_0_OAI21X1_573 gnd vdd FILL
XFILL_0_OAI21X1_562 gnd vdd FILL
XFILL_0_OAI21X1_584 gnd vdd FILL
XFILL_1_OAI21X1_766 gnd vdd FILL
XFILL_0_OAI21X1_595 gnd vdd FILL
XFILL_1_OAI21X1_777 gnd vdd FILL
XFILL_1_OAI21X1_788 gnd vdd FILL
XFILL_2_OAI21X1_959 gnd vdd FILL
XFILL_1_OAI21X1_799 gnd vdd FILL
XFILL_28_5_1 gnd vdd FILL
XBUFX2_609 BUFX2_609/A gnd majID4_o[33] vdd BUFX2
XFILL_27_0_0 gnd vdd FILL
XFILL_0_CLKBUF1_73 gnd vdd FILL
XFILL_0_CLKBUF1_40 gnd vdd FILL
XFILL_2_0_0 gnd vdd FILL
XFILL_3_5_1 gnd vdd FILL
XFILL_0_CLKBUF1_51 gnd vdd FILL
XFILL_0_CLKBUF1_62 gnd vdd FILL
XFILL_0_CLKBUF1_95 gnd vdd FILL
XFILL_0_CLKBUF1_84 gnd vdd FILL
XFILL_1_NAND2X1_750 gnd vdd FILL
XFILL_0_OAI21X1_1350 gnd vdd FILL
XFILL_1_NAND2X1_761 gnd vdd FILL
XFILL_0_NAND2X1_590 gnd vdd FILL
XFILL_0_DFFPOSX1_951 gnd vdd FILL
XFILL_0_DFFPOSX1_940 gnd vdd FILL
XFILL_0_OAI21X1_1394 gnd vdd FILL
XFILL_0_OAI21X1_1383 gnd vdd FILL
XFILL_0_OAI21X1_1372 gnd vdd FILL
XFILL_0_OAI21X1_1361 gnd vdd FILL
XFILL_0_DFFPOSX1_962 gnd vdd FILL
XFILL_0_DFFPOSX1_984 gnd vdd FILL
XFILL_0_DFFPOSX1_995 gnd vdd FILL
XFILL_0_DFFPOSX1_973 gnd vdd FILL
XFILL_11_4_1 gnd vdd FILL
XINVX2_105 INVX2_105/A gnd INVX2_105/Y vdd INVX2
XFILL_0_BUFX2_305 gnd vdd FILL
XFILL_0_OR2X2_1 gnd vdd FILL
XFILL_0_BUFX2_338 gnd vdd FILL
XFILL_0_BUFX2_327 gnd vdd FILL
XINVX2_127 bundlePid_i[21] gnd INVX2_127/Y vdd INVX2
XINVX2_138 bundlePid_i[10] gnd INVX2_138/Y vdd INVX2
XFILL_20_15_0 gnd vdd FILL
XFILL_0_BUFX2_316 gnd vdd FILL
XINVX2_116 bundlePid_i[0] gnd INVX2_116/Y vdd INVX2
XFILL_0_BUFX2_349 gnd vdd FILL
XINVX2_149 bundleTid_i[60] gnd INVX2_149/Y vdd INVX2
XFILL_19_5_1 gnd vdd FILL
XFILL_2_NOR3X1_11 gnd vdd FILL
XFILL_18_0_0 gnd vdd FILL
XFILL_2_OAI21X1_1444 gnd vdd FILL
XFILL_0_INVX1_3 gnd vdd FILL
XFILL_25_14_0 gnd vdd FILL
XFILL_1_NAND3X1_12 gnd vdd FILL
XFILL_1_OAI21X1_1023 gnd vdd FILL
XFILL_1_NAND3X1_45 gnd vdd FILL
XFILL_1_NAND3X1_34 gnd vdd FILL
XFILL_1_NAND3X1_23 gnd vdd FILL
XDFFPOSX1_404 BUFX2_436/A CLKBUF1_79/Y OAI21X1_376/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1001 gnd vdd FILL
XFILL_1_OAI21X1_1012 gnd vdd FILL
XFILL_0_BUFX2_861 gnd vdd FILL
XFILL_0_BUFX2_850 gnd vdd FILL
XDFFPOSX1_415 BUFX2_448/A CLKBUF1_11/Y OAI21X1_387/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1045 gnd vdd FILL
XFILL_1_DFFPOSX1_624 gnd vdd FILL
XFILL_1_DFFPOSX1_613 gnd vdd FILL
XFILL_1_NAND3X1_56 gnd vdd FILL
XFILL_1_NAND3X1_67 gnd vdd FILL
XFILL_1_DFFPOSX1_602 gnd vdd FILL
XDFFPOSX1_426 BUFX2_513/A CLKBUF1_10/Y OAI21X1_407/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1034 gnd vdd FILL
XDFFPOSX1_437 BUFX2_466/A CLKBUF1_24/Y OAI21X1_425/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1056 gnd vdd FILL
XFILL_0_BUFX2_883 gnd vdd FILL
XFILL_0_BUFX2_872 gnd vdd FILL
XFILL_0_BUFX2_894 gnd vdd FILL
XFILL_1_OAI21X1_1067 gnd vdd FILL
XDFFPOSX1_459 BUFX2_490/A CLKBUF1_5/Y OAI21X1_457/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1078 gnd vdd FILL
XFILL_1_OAI21X1_1089 gnd vdd FILL
XFILL_1_DFFPOSX1_635 gnd vdd FILL
XFILL_1_DFFPOSX1_657 gnd vdd FILL
XFILL_1_DFFPOSX1_646 gnd vdd FILL
XINVX1_160 bundle_i[108] gnd INVX1_160/Y vdd INVX1
XDFFPOSX1_448 BUFX2_478/A CLKBUF1_33/Y OAI21X1_443/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_679 gnd vdd FILL
XINVX1_171 bundle_i[97] gnd INVX1_171/Y vdd INVX1
XFILL_1_DFFPOSX1_668 gnd vdd FILL
XINVX1_182 BUFX2_88/A gnd INVX1_182/Y vdd INVX1
XNAND2X1_518 bundleAddress_i[39] bundleAddress_i[38] gnd NOR2X1_142/B vdd NAND2X1
XINVX1_193 INVX1_193/A gnd INVX1_193/Y vdd INVX1
XNAND2X1_507 bundleAddress_i[43] NOR2X1_137/Y gnd NAND2X1_507/Y vdd NAND2X1
XNAND2X1_529 BUFX4_238/Y NOR2X1_148/B gnd NAND2X1_529/Y vdd NAND2X1
XFILL_6_DFFPOSX1_250 gnd vdd FILL
XFILL_0_INVX2_81 gnd vdd FILL
XFILL_0_INVX2_70 gnd vdd FILL
XFILL_0_INVX2_92 gnd vdd FILL
XFILL_1_NOR3X1_1 gnd vdd FILL
XFILL_0_AND2X2_19 gnd vdd FILL
XFILL_0_DFFPOSX1_214 gnd vdd FILL
XFILL_0_DFFPOSX1_203 gnd vdd FILL
XFILL_0_15_0 gnd vdd FILL
XFILL_0_DFFPOSX1_247 gnd vdd FILL
XFILL_0_DFFPOSX1_225 gnd vdd FILL
XFILL_0_DFFPOSX1_236 gnd vdd FILL
XFILL_0_DFFPOSX1_258 gnd vdd FILL
XFILL_0_DFFPOSX1_269 gnd vdd FILL
XFILL_3_DFFPOSX1_718 gnd vdd FILL
XFILL_3_DFFPOSX1_729 gnd vdd FILL
XFILL_3_DFFPOSX1_707 gnd vdd FILL
XFILL_3_CLKBUF1_39 gnd vdd FILL
XFILL_3_CLKBUF1_17 gnd vdd FILL
XFILL_3_CLKBUF1_28 gnd vdd FILL
XOAI21X1_1392 bundleAddress_i[61] bundleAddress_i[60] bundleAddress_i[59] gnd OAI21X1_1393/C
+ vdd OAI21X1
XOAI21X1_1381 AOI21X1_59/Y OAI21X1_1381/B OAI21X1_1381/C gnd OAI21X1_1381/Y vdd OAI21X1
XDFFPOSX1_960 BUFX2_210/A CLKBUF1_35/Y OAI21X1_1455/Y gnd vdd DFFPOSX1
XOAI21X1_1370 BUFX4_6/A BUFX4_364/Y BUFX2_183/A gnd OAI21X1_1371/C vdd OAI21X1
XFILL_1_OAI21X1_1590 gnd vdd FILL
XDFFPOSX1_982 BUFX2_234/A CLKBUF1_68/Y OAI21X1_1524/Y gnd vdd DFFPOSX1
XFILL_1_NOR2X1_113 gnd vdd FILL
XDFFPOSX1_993 INVX1_227/A CLKBUF1_20/Y OAI21X1_1557/Y gnd vdd DFFPOSX1
XDFFPOSX1_971 BUFX2_222/A CLKBUF1_81/Y OAI21X1_1488/Y gnd vdd DFFPOSX1
XFILL_1_NOR2X1_124 gnd vdd FILL
XFILL_1_NOR2X1_146 gnd vdd FILL
XFILL_0_OAI21X1_370 gnd vdd FILL
XFILL_0_OAI21X1_381 gnd vdd FILL
XFILL_2_OAI21X1_734 gnd vdd FILL
XFILL_1_OAI21X1_541 gnd vdd FILL
XFILL_1_OAI21X1_552 gnd vdd FILL
XFILL_1_NOR2X1_135 gnd vdd FILL
XFILL_1_OAI21X1_563 gnd vdd FILL
XFILL_1_OAI21X1_530 gnd vdd FILL
XFILL_1_NOR2X1_179 gnd vdd FILL
XFILL_2_OAI21X1_745 gnd vdd FILL
XFILL_2_OAI21X1_756 gnd vdd FILL
XFILL_1_OAI21X1_596 gnd vdd FILL
XFILL_0_OAI21X1_392 gnd vdd FILL
XFILL_1_NOR2X1_157 gnd vdd FILL
XFILL_1_OAI21X1_585 gnd vdd FILL
XFILL_1_OAI21X1_574 gnd vdd FILL
XFILL_5_14_0 gnd vdd FILL
XFILL_2_DFFPOSX1_319 gnd vdd FILL
XFILL_2_DFFPOSX1_308 gnd vdd FILL
XBUFX2_406 BUFX2_406/A gnd majID1_o[43] vdd BUFX2
XBUFX2_417 BUFX2_417/A gnd majID1_o[33] vdd BUFX2
XBUFX2_439 BUFX2_439/A gnd majID1_o[13] vdd BUFX2
XBUFX2_428 BUFX2_428/A gnd majID1_o[23] vdd BUFX2
XFILL_1_BUFX4_322 gnd vdd FILL
XFILL_1_BUFX4_311 gnd vdd FILL
XFILL_1_BUFX4_300 gnd vdd FILL
XFILL_1_NAND2X1_591 gnd vdd FILL
XFILL_1_BUFX4_344 gnd vdd FILL
XFILL_0_DFFPOSX1_770 gnd vdd FILL
XFILL_0_OAI21X1_1180 gnd vdd FILL
XFILL_1_BUFX4_333 gnd vdd FILL
XFILL_1_BUFX4_355 gnd vdd FILL
XFILL_0_OAI21X1_1191 gnd vdd FILL
XFILL_1_BUFX4_377 gnd vdd FILL
XFILL_1_BUFX4_366 gnd vdd FILL
XFILL_0_DFFPOSX1_792 gnd vdd FILL
XFILL_1_BUFX4_388 gnd vdd FILL
XFILL_0_DFFPOSX1_781 gnd vdd FILL
XFILL_0_BUFX2_102 gnd vdd FILL
XFILL_0_BUFX2_113 gnd vdd FILL
XFILL_0_BUFX2_135 gnd vdd FILL
XFILL_0_BUFX2_124 gnd vdd FILL
XFILL_0_BUFX2_146 gnd vdd FILL
XFILL_0_BUFX2_157 gnd vdd FILL
XFILL_0_BUFX2_168 gnd vdd FILL
XFILL_0_BUFX2_179 gnd vdd FILL
XFILL_2_OAI21X1_1241 gnd vdd FILL
XFILL_14_11_1 gnd vdd FILL
XFILL_2_DFFPOSX1_820 gnd vdd FILL
XFILL_2_DFFPOSX1_842 gnd vdd FILL
XBUFX2_940 BUFX2_940/A gnd tid3_o[23] vdd BUFX2
XFILL_2_DFFPOSX1_831 gnd vdd FILL
XBUFX2_973 BUFX2_973/A gnd tid4_o[51] vdd BUFX2
XBUFX2_951 BUFX2_951/A gnd tid3_o[13] vdd BUFX2
XFILL_2_DFFPOSX1_875 gnd vdd FILL
XFILL_34_3_1 gnd vdd FILL
XFILL_2_DFFPOSX1_853 gnd vdd FILL
XFILL_2_DFFPOSX1_864 gnd vdd FILL
XBUFX2_962 BUFX2_962/A gnd tid3_o[3] vdd BUFX2
XFILL_2_DFFPOSX1_886 gnd vdd FILL
XBUFX2_984 BUFX2_984/A gnd tid4_o[41] vdd BUFX2
XFILL_2_DFFPOSX1_897 gnd vdd FILL
XBUFX2_995 BUFX2_995/A gnd tid4_o[31] vdd BUFX2
XOAI21X1_309 INVX2_200/Y BUFX4_290/Y OAI21X1_309/C gnd OAI21X1_309/Y vdd OAI21X1
XDFFPOSX1_212 BUFX2_884/A CLKBUF1_14/Y OAI21X1_56/Y gnd vdd DFFPOSX1
XDFFPOSX1_201 BUFX2_872/A CLKBUF1_98/Y OAI21X1_45/Y gnd vdd DFFPOSX1
XBUFX4_7 BUFX4_7/A gnd BUFX4_7/Y vdd BUFX4
XDFFPOSX1_245 BUFX2_914/A CLKBUF1_74/Y OAI21X1_107/Y gnd vdd DFFPOSX1
XDFFPOSX1_234 BUFX2_961/A CLKBUF1_86/Y OAI21X1_85/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_421 gnd vdd FILL
XFILL_1_DFFPOSX1_410 gnd vdd FILL
XDFFPOSX1_223 BUFX2_896/A CLKBUF1_51/Y OAI21X1_67/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_432 gnd vdd FILL
XFILL_0_BUFX2_680 gnd vdd FILL
XDFFPOSX1_278 BUFX2_951/A CLKBUF1_59/Y OAI21X1_173/Y gnd vdd DFFPOSX1
XDFFPOSX1_289 BUFX2_963/A CLKBUF1_55/Y OAI21X1_195/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_691 gnd vdd FILL
XDFFPOSX1_267 BUFX2_938/A CLKBUF1_40/Y OAI21X1_151/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_443 gnd vdd FILL
XFILL_1_DFFPOSX1_465 gnd vdd FILL
XDFFPOSX1_256 BUFX2_926/A CLKBUF1_71/Y OAI21X1_129/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_454 gnd vdd FILL
XNAND2X1_304 OAI21X1_642/Y OAI21X1_645/A gnd OAI21X1_643/A vdd NAND2X1
XFILL_19_10_1 gnd vdd FILL
XFILL_1_DFFPOSX1_476 gnd vdd FILL
XNAND2X1_326 bundleStartMajId_i[29] NOR2X1_110/Y gnd INVX1_41/A vdd NAND2X1
XFILL_1_DFFPOSX1_498 gnd vdd FILL
XNAND2X1_315 bundleStartMajId_i[47] NOR2X1_105/Y gnd INVX1_36/A vdd NAND2X1
XFILL_1_DFFPOSX1_487 gnd vdd FILL
XFILL_4_DFFPOSX1_903 gnd vdd FILL
XNAND2X1_337 OAI21X1_839/A NAND2X1_337/B gnd OAI21X1_834/A vdd NAND2X1
XFILL_4_DFFPOSX1_914 gnd vdd FILL
XNAND2X1_348 BUFX4_268/Y bundle_i[21] gnd OAI21X1_854/C vdd NAND2X1
XNAND2X1_359 BUFX4_262/Y bundle_i[10] gnd OAI21X1_865/C vdd NAND2X1
XFILL_4_DFFPOSX1_936 gnd vdd FILL
XFILL_4_DFFPOSX1_947 gnd vdd FILL
XFILL_4_DFFPOSX1_925 gnd vdd FILL
XFILL_32_12_1 gnd vdd FILL
XFILL_4_DFFPOSX1_969 gnd vdd FILL
XNOR3X1_11 INVX2_38/Y INVX4_28/Y NOR3X1_11/C gnd NOR3X1_11/Y vdd NOR3X1
XFILL_4_DFFPOSX1_958 gnd vdd FILL
XFILL_25_3_1 gnd vdd FILL
XFILL_0_3_1 gnd vdd FILL
XFILL_1_BUFX2_804 gnd vdd FILL
XFILL_1_INVX2_26 gnd vdd FILL
XFILL_0_XNOR2X1_3 gnd vdd FILL
XINVX4_7 bundleStartMajId_i[46] gnd INVX4_7/Y vdd INVX4
XFILL_1_INVX2_48 gnd vdd FILL
XFILL_1_BUFX2_837 gnd vdd FILL
XFILL_1_BUFX2_848 gnd vdd FILL
XOAI21X1_832 NOR2X1_117/Y OAI21X1_832/B OAI21X1_832/C gnd OAI21X1_832/Y vdd OAI21X1
XOAI21X1_810 NOR3X1_8/C NOR3X1_8/B NOR3X1_8/A gnd OAI21X1_811/C vdd OAI21X1
XOAI21X1_821 OAI21X1_821/A BUFX4_295/Y OAI21X1_821/C gnd OAI21X1_821/Y vdd OAI21X1
XFILL_3_DFFPOSX1_504 gnd vdd FILL
XFILL_3_DFFPOSX1_515 gnd vdd FILL
XFILL_3_DFFPOSX1_537 gnd vdd FILL
XFILL_3_DFFPOSX1_526 gnd vdd FILL
XOAI21X1_843 OAI21X1_843/A NOR2X1_120/Y OAI21X1_843/C gnd OAI21X1_843/Y vdd OAI21X1
XOAI21X1_876 INVX1_77/Y BUFX4_180/Y OAI21X1_876/C gnd OAI21X1_876/Y vdd OAI21X1
XOAI21X1_854 INVX1_55/Y BUFX4_268/Y OAI21X1_854/C gnd OAI21X1_854/Y vdd OAI21X1
XOAI21X1_865 INVX1_66/Y BUFX4_262/Y OAI21X1_865/C gnd OAI21X1_865/Y vdd OAI21X1
XOAI21X1_898 INVX1_99/Y BUFX4_220/Y OAI21X1_898/C gnd OAI21X1_898/Y vdd OAI21X1
XFILL_3_DFFPOSX1_548 gnd vdd FILL
XFILL_3_DFFPOSX1_559 gnd vdd FILL
XOAI21X1_887 INVX1_88/Y BUFX4_232/Y OAI21X1_887/C gnd OAI21X1_887/Y vdd OAI21X1
XFILL_37_11_1 gnd vdd FILL
XDFFPOSX1_790 BUFX2_42/A CLKBUF1_30/Y OAI21X1_1082/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_371 gnd vdd FILL
XFILL_1_OAI21X1_360 gnd vdd FILL
XFILL_8_4_1 gnd vdd FILL
XFILL_1_CLKBUF1_3 gnd vdd FILL
XFILL_2_OAI21X1_553 gnd vdd FILL
XFILL_1_OAI21X1_382 gnd vdd FILL
XFILL_1_OAI21X1_393 gnd vdd FILL
XFILL_0_NAND3X1_20 gnd vdd FILL
XFILL_2_DFFPOSX1_127 gnd vdd FILL
XBUFX2_203 BUFX2_203/A gnd addr4_o[45] vdd BUFX2
XBUFX2_214 BUFX2_214/A gnd addr4_o[35] vdd BUFX2
XFILL_2_DFFPOSX1_116 gnd vdd FILL
XFILL_0_NAND3X1_42 gnd vdd FILL
XFILL_0_NAND3X1_31 gnd vdd FILL
XFILL_0_NAND3X1_53 gnd vdd FILL
XBUFX2_225 BUFX2_225/A gnd addr4_o[25] vdd BUFX2
XFILL_2_DFFPOSX1_105 gnd vdd FILL
XFILL_2_DFFPOSX1_138 gnd vdd FILL
XBUFX2_269 INVX1_61/A gnd instr1_o[15] vdd BUFX2
XFILL_2_DFFPOSX1_149 gnd vdd FILL
XBUFX2_258 BUFX2_258/A gnd enable2_o vdd BUFX2
XFILL_0_NAND3X1_64 gnd vdd FILL
XBUFX2_236 BUFX2_236/A gnd addr4_o[15] vdd BUFX2
XBUFX2_247 BUFX2_247/A gnd addr4_o[5] vdd BUFX2
XFILL_16_3_1 gnd vdd FILL
XFILL_5_DFFPOSX1_609 gnd vdd FILL
XFILL_1_BUFX4_130 gnd vdd FILL
XFILL_1_BUFX4_141 gnd vdd FILL
XFILL_1_BUFX4_152 gnd vdd FILL
XFILL_1_BUFX4_163 gnd vdd FILL
XFILL_1_BUFX4_174 gnd vdd FILL
XFILL_1_BUFX4_185 gnd vdd FILL
XFILL_1_BUFX4_196 gnd vdd FILL
XFILL_2_CLKBUF1_14 gnd vdd FILL
XFILL_2_CLKBUF1_25 gnd vdd FILL
XFILL_2_CLKBUF1_47 gnd vdd FILL
XFILL_2_CLKBUF1_36 gnd vdd FILL
XFILL_2_DFFPOSX1_650 gnd vdd FILL
XFILL_2_CLKBUF1_69 gnd vdd FILL
XFILL_2_CLKBUF1_58 gnd vdd FILL
XFILL_2_DFFPOSX1_672 gnd vdd FILL
XFILL_2_DFFPOSX1_683 gnd vdd FILL
XBUFX2_781 BUFX2_781/A gnd tid1_o[51] vdd BUFX2
XFILL_2_DFFPOSX1_661 gnd vdd FILL
XBUFX2_770 BUFX2_770/A gnd pid4_o[0] vdd BUFX2
XFILL_2_DFFPOSX1_694 gnd vdd FILL
XFILL_0_NOR2X1_121 gnd vdd FILL
XBUFX2_792 BUFX2_792/A gnd tid1_o[41] vdd BUFX2
XFILL_0_NOR2X1_110 gnd vdd FILL
XFILL_0_NOR2X1_132 gnd vdd FILL
XFILL_0_NOR2X1_143 gnd vdd FILL
XFILL_0_NOR2X1_154 gnd vdd FILL
XOAI21X1_106 BUFX4_101/Y BUFX4_312/Y BUFX2_914/A gnd OAI21X1_107/C vdd OAI21X1
XOAI21X1_117 BUFX4_162/Y INVX2_168/Y OAI21X1_117/C gnd OAI21X1_117/Y vdd OAI21X1
XFILL_0_NOR2X1_165 gnd vdd FILL
XFILL_0_NOR2X1_176 gnd vdd FILL
XFILL_0_NOR2X1_187 gnd vdd FILL
XFILL_0_NOR2X1_198 gnd vdd FILL
XOAI21X1_128 BUFX4_1/A BUFX4_343/Y BUFX2_926/A gnd OAI21X1_129/C vdd OAI21X1
XOAI21X1_139 BUFX4_143/Y INVX2_179/Y OAI21X1_139/C gnd OAI21X1_139/Y vdd OAI21X1
XFILL_0_DFFPOSX1_1017 gnd vdd FILL
XFILL_0_DFFPOSX1_1006 gnd vdd FILL
XFILL_0_DFFPOSX1_1028 gnd vdd FILL
XBUFX2_4 BUFX2_4/A gnd addr1_o[52] vdd BUFX2
XFILL_1_DFFPOSX1_240 gnd vdd FILL
XFILL_1_DFFPOSX1_273 gnd vdd FILL
XFILL_1_DFFPOSX1_262 gnd vdd FILL
XFILL_1_DFFPOSX1_251 gnd vdd FILL
XNAND2X1_101 BUFX2_415/A BUFX4_314/Y gnd OAI21X1_357/C vdd NAND2X1
XFILL_1_DFFPOSX1_284 gnd vdd FILL
XNAND2X1_134 BUFX2_452/A BUFX4_356/Y gnd OAI21X1_390/C vdd NAND2X1
XNAND2X1_123 BUFX2_440/A BUFX4_323/Y gnd OAI21X1_379/C vdd NAND2X1
XFILL_1_DFFPOSX1_295 gnd vdd FILL
XNAND2X1_112 BUFX2_428/A BUFX4_365/Y gnd OAI21X1_368/C vdd NAND2X1
XFILL_4_DFFPOSX1_700 gnd vdd FILL
XFILL_4_DFFPOSX1_711 gnd vdd FILL
XFILL_4_DFFPOSX1_722 gnd vdd FILL
XNAND2X1_178 bundleStartMajId_i[44] bundleStartMajId_i[43] gnd OR2X2_2/B vdd NAND2X1
XNAND2X1_156 BUFX2_459/A BUFX4_181/Y gnd OAI21X1_415/C vdd NAND2X1
XNAND2X1_145 bundleStartMajId_i[59] bundleStartMajId_i[58] gnd NOR2X1_4/A vdd NAND2X1
XNAND2X1_167 NOR2X1_7/Y AND2X2_2/B gnd NOR2X1_11/B vdd NAND2X1
XFILL_1_OAI21X1_32 gnd vdd FILL
XFILL_4_DFFPOSX1_755 gnd vdd FILL
XFILL_4_DFFPOSX1_744 gnd vdd FILL
XNAND2X1_189 BUFX2_475/A BUFX4_209/Y gnd OAI21X1_437/C vdd NAND2X1
XFILL_1_OAI21X1_43 gnd vdd FILL
XFILL_4_DFFPOSX1_733 gnd vdd FILL
XFILL_1_OAI21X1_10 gnd vdd FILL
XFILL_1_OAI21X1_21 gnd vdd FILL
XFILL_1_OAI21X1_65 gnd vdd FILL
XFILL_4_DFFPOSX1_788 gnd vdd FILL
XFILL_4_DFFPOSX1_777 gnd vdd FILL
XFILL_1_OAI21X1_54 gnd vdd FILL
XFILL_1_OAI21X1_76 gnd vdd FILL
XFILL_4_DFFPOSX1_766 gnd vdd FILL
XFILL_1_OAI21X1_87 gnd vdd FILL
XFILL_4_DFFPOSX1_799 gnd vdd FILL
XFILL_1_OAI21X1_98 gnd vdd FILL
XFILL_0_DFFPOSX1_8 gnd vdd FILL
XFILL_1_BUFX2_601 gnd vdd FILL
XFILL_1_BUFX2_634 gnd vdd FILL
XFILL_1_BUFX2_645 gnd vdd FILL
XINVX2_4 bundleTid_i[3] gnd INVX2_4/Y vdd INVX2
XFILL_1_BUFX2_656 gnd vdd FILL
XFILL_1_BUFX2_678 gnd vdd FILL
XFILL_0_BUFX4_208 gnd vdd FILL
XOAI21X1_651 AOI21X1_25/Y OAI21X1_651/B OAI21X1_651/C gnd OAI21X1_651/Y vdd OAI21X1
XFILL_3_DFFPOSX1_301 gnd vdd FILL
XFILL_3_DFFPOSX1_312 gnd vdd FILL
XFILL_0_BUFX4_219 gnd vdd FILL
XFILL_23_17_1 gnd vdd FILL
XOAI21X1_640 OAI21X1_640/A AOI21X1_21/Y OAI21X1_640/C gnd OAI21X1_640/Y vdd OAI21X1
XFILL_1_BUFX2_689 gnd vdd FILL
XFILL_3_DFFPOSX1_345 gnd vdd FILL
XFILL_3_DFFPOSX1_323 gnd vdd FILL
XAOI21X1_4 INVX1_43/A INVX1_22/Y bundleStartMajId_i[4] gnd AOI21X1_4/Y vdd AOI21X1
XOAI21X1_662 bundleStartMajId_i[63] bundleStartMajId_i[62] bundleStartMajId_i[61]
+ gnd OAI21X1_663/C vdd OAI21X1
XOAI21X1_684 BUFX4_167/Y BUFX4_30/Y BUFX2_648/A gnd OAI21X1_685/C vdd OAI21X1
XOAI21X1_673 NOR2X1_4/A INVX2_52/Y OAI21X1_673/C gnd OAI21X1_675/A vdd OAI21X1
XFILL_3_DFFPOSX1_334 gnd vdd FILL
XFILL_3_DFFPOSX1_356 gnd vdd FILL
XOAI21X1_695 AND2X2_20/A OAI21X1_695/B OAI21X1_695/C gnd OAI21X1_695/Y vdd OAI21X1
XFILL_3_DFFPOSX1_378 gnd vdd FILL
XFILL_3_DFFPOSX1_367 gnd vdd FILL
XFILL_3_DFFPOSX1_389 gnd vdd FILL
XFILL_0_INVX4_27 gnd vdd FILL
XFILL_0_INVX4_16 gnd vdd FILL
XFILL_0_INVX4_38 gnd vdd FILL
XXNOR2X1_23 XNOR2X1_23/A INVX4_26/Y gnd XNOR2X1_23/Y vdd XNOR2X1
XFILL_0_INVX4_49 gnd vdd FILL
XXNOR2X1_12 NOR3X1_1/Y bundleStartMajId_i[33] gnd XNOR2X1_12/Y vdd XNOR2X1
XFILL_1_INVX2_130 gnd vdd FILL
XXNOR2X1_56 INVX2_95/A bundleAddress_i[52] gnd XNOR2X1_56/Y vdd XNOR2X1
XXNOR2X1_45 XNOR2X1_45/A INVX4_9/Y gnd XNOR2X1_45/Y vdd XNOR2X1
XXNOR2X1_34 NOR2X1_75/Y bundleStartMajId_i[30] gnd XNOR2X1_34/Y vdd XNOR2X1
XNAND2X1_690 BUFX2_711/A BUFX4_193/Y gnd NAND2X1_690/Y vdd NAND2X1
XXNOR2X1_89 XNOR2X1_89/A INVX4_46/Y gnd XNOR2X1_89/Y vdd XNOR2X1
XXNOR2X1_78 NOR3X1_18/C INVX4_35/Y gnd XNOR2X1_78/Y vdd XNOR2X1
XFILL_1_OAI21X1_190 gnd vdd FILL
XXNOR2X1_67 XNOR2X1_67/A bundleAddress_i[28] gnd XNOR2X1_67/Y vdd XNOR2X1
XINVX1_91 bundle_i[49] gnd INVX1_91/Y vdd INVX1
XFILL_0_NAND2X1_408 gnd vdd FILL
XBUFX2_11 BUFX2_11/A gnd addr1_o[45] vdd BUFX2
XINVX1_80 bundle_i[60] gnd INVX1_80/Y vdd INVX1
XFILL_0_NAND2X1_419 gnd vdd FILL
XBUFX2_22 BUFX2_22/A gnd addr1_o[35] vdd BUFX2
XBUFX2_44 BUFX2_44/A gnd addr1_o[15] vdd BUFX2
XBUFX2_33 BUFX2_33/A gnd addr1_o[25] vdd BUFX2
XBUFX2_77 BUFX2_77/A gnd addr2_o[61] vdd BUFX2
XBUFX2_66 BUFX2_66/A gnd addr2_o[62] vdd BUFX2
XBUFX2_55 BUFX2_55/A gnd addr1_o[5] vdd BUFX2
XBUFX2_99 BUFX2_99/A gnd addr2_o[59] vdd BUFX2
XBUFX2_88 BUFX2_88/A gnd addr2_o[60] vdd BUFX2
XFILL_31_1_1 gnd vdd FILL
XFILL_28_16_1 gnd vdd FILL
XFILL_5_DFFPOSX1_406 gnd vdd FILL
XFILL_5_DFFPOSX1_417 gnd vdd FILL
XFILL_1_BUFX4_11 gnd vdd FILL
XFILL_5_DFFPOSX1_439 gnd vdd FILL
XFILL_5_DFFPOSX1_428 gnd vdd FILL
XFILL_1_BUFX4_44 gnd vdd FILL
XFILL_1_BUFX4_22 gnd vdd FILL
XFILL_1_BUFX4_33 gnd vdd FILL
XFILL_1_BUFX4_55 gnd vdd FILL
XFILL_1_BUFX4_77 gnd vdd FILL
XFILL_22_12_0 gnd vdd FILL
XFILL_1_BUFX4_88 gnd vdd FILL
XFILL_1_BUFX4_66 gnd vdd FILL
XFILL_1_BUFX4_99 gnd vdd FILL
XFILL_0_OAI21X1_914 gnd vdd FILL
XFILL_3_DFFPOSX1_890 gnd vdd FILL
XNOR2X1_2 NOR2X1_2/A INVX1_7/Y gnd NOR2X1_2/Y vdd NOR2X1
XFILL_0_OAI21X1_903 gnd vdd FILL
XFILL_0_OAI21X1_936 gnd vdd FILL
XFILL_0_OAI21X1_925 gnd vdd FILL
XFILL_0_OAI21X1_947 gnd vdd FILL
XFILL_0_OAI21X1_969 gnd vdd FILL
XFILL_0_OAI21X1_958 gnd vdd FILL
XFILL_1_OR2X2_14 gnd vdd FILL
XFILL_3_17_1 gnd vdd FILL
XFILL_0_OAI21X1_1713 gnd vdd FILL
XFILL_0_OAI21X1_1724 gnd vdd FILL
XFILL_0_OAI21X1_1702 gnd vdd FILL
XFILL_0_OAI21X1_1757 gnd vdd FILL
XFILL_0_OAI21X1_1746 gnd vdd FILL
XFILL_2_DFFPOSX1_480 gnd vdd FILL
XFILL_0_OAI21X1_1768 gnd vdd FILL
XFILL_0_OAI21X1_1735 gnd vdd FILL
XFILL_2_DFFPOSX1_491 gnd vdd FILL
XFILL_22_1_1 gnd vdd FILL
XFILL_0_OAI21X1_1779 gnd vdd FILL
XFILL_27_11_0 gnd vdd FILL
XFILL_5_DFFPOSX1_940 gnd vdd FILL
XFILL_5_DFFPOSX1_962 gnd vdd FILL
XFILL_5_DFFPOSX1_951 gnd vdd FILL
XFILL_5_DFFPOSX1_973 gnd vdd FILL
XFILL_5_DFFPOSX1_984 gnd vdd FILL
XAOI21X1_23 AOI21X1_23/A OR2X2_12/Y NOR2X1_96/Y gnd AOI21X1_23/Y vdd AOI21X1
XFILL_5_DFFPOSX1_995 gnd vdd FILL
XAOI21X1_34 bundleStartMajId_i[10] NOR3X1_8/Y bundleStartMajId_i[9] gnd AOI21X1_34/Y
+ vdd AOI21X1
XAOI21X1_12 AOI21X1_12/A NAND3X1_19/Y NOR2X1_81/Y gnd AOI21X1_12/Y vdd AOI21X1
XFILL_0_NOR2X1_19 gnd vdd FILL
XAOI21X1_45 INVX1_199/A NOR2X1_174/B bundleAddress_i[2] gnd AOI21X1_45/Y vdd AOI21X1
XAOI21X1_56 bundleAddress_i[10] XNOR2X1_87/A bundleAddress_i[9] gnd AOI21X1_56/Y vdd
+ AOI21X1
XOAI21X1_7 OAI21X1_7/A INVX2_7/Y OAI21X1_7/C gnd OAI21X1_7/Y vdd OAI21X1
XXNOR2X1_104 NAND3X1_69/Y INVX4_46/Y gnd XNOR2X1_104/Y vdd XNOR2X1
XFILL_8_16_1 gnd vdd FILL
XBUFX4_309 BUFX4_310/A gnd INVX8_6/A vdd BUFX4
XFILL_4_DFFPOSX1_530 gnd vdd FILL
XFILL_5_2_1 gnd vdd FILL
XFILL_4_DFFPOSX1_541 gnd vdd FILL
XFILL_4_DFFPOSX1_563 gnd vdd FILL
XFILL_4_DFFPOSX1_552 gnd vdd FILL
XFILL_4_DFFPOSX1_585 gnd vdd FILL
XFILL_4_DFFPOSX1_596 gnd vdd FILL
XFILL_4_DFFPOSX1_574 gnd vdd FILL
XFILL_2_12_0 gnd vdd FILL
XFILL_1_BUFX2_1032 gnd vdd FILL
XFILL_13_1_1 gnd vdd FILL
XFILL_1_BUFX2_431 gnd vdd FILL
XFILL_1_BUFX2_442 gnd vdd FILL
XFILL_1_BUFX2_453 gnd vdd FILL
XFILL_1_CLKBUF1_11 gnd vdd FILL
XFILL_1_CLKBUF1_22 gnd vdd FILL
XFILL_1_BUFX2_486 gnd vdd FILL
XFILL_1_BUFX2_497 gnd vdd FILL
XFILL_3_DFFPOSX1_120 gnd vdd FILL
XFILL_3_DFFPOSX1_153 gnd vdd FILL
XFILL_3_DFFPOSX1_164 gnd vdd FILL
XFILL_1_OAI21X1_1408 gnd vdd FILL
XFILL_1_OAI21X1_1419 gnd vdd FILL
XFILL_3_DFFPOSX1_131 gnd vdd FILL
XOAI21X1_492 AOI21X1_4/Y OAI21X1_492/B OAI21X1_492/C gnd OAI21X1_492/Y vdd OAI21X1
XFILL_1_CLKBUF1_55 gnd vdd FILL
XFILL_1_INVX8_6 gnd vdd FILL
XFILL_1_CLKBUF1_44 gnd vdd FILL
XFILL_1_CLKBUF1_33 gnd vdd FILL
XFILL_3_DFFPOSX1_142 gnd vdd FILL
XOAI21X1_481 XNOR2X1_22/Y BUFX4_182/Y OAI21X1_481/C gnd OAI21X1_481/Y vdd OAI21X1
XOAI21X1_470 INVX1_16/Y NOR3X1_9/B BUFX4_244/Y gnd OAI21X1_471/B vdd OAI21X1
XFILL_3_DFFPOSX1_175 gnd vdd FILL
XFILL_3_DFFPOSX1_197 gnd vdd FILL
XFILL_3_DFFPOSX1_186 gnd vdd FILL
XFILL_1_CLKBUF1_88 gnd vdd FILL
XFILL_1_CLKBUF1_77 gnd vdd FILL
XFILL_1_CLKBUF1_66 gnd vdd FILL
XFILL_1_CLKBUF1_99 gnd vdd FILL
XFILL_6_DFFPOSX1_624 gnd vdd FILL
XFILL_6_DFFPOSX1_635 gnd vdd FILL
XFILL_6_DFFPOSX1_679 gnd vdd FILL
XFILL_6_DFFPOSX1_668 gnd vdd FILL
XFILL_6_DFFPOSX1_657 gnd vdd FILL
XFILL_6_DFFPOSX1_646 gnd vdd FILL
XFILL_7_11_0 gnd vdd FILL
XFILL_0_NAND2X1_216 gnd vdd FILL
XFILL_0_NAND2X1_205 gnd vdd FILL
XFILL_0_NAND2X1_238 gnd vdd FILL
XFILL_0_NAND2X1_249 gnd vdd FILL
XFILL_0_NAND2X1_227 gnd vdd FILL
XFILL_0_OAI21X1_1009 gnd vdd FILL
XFILL_33_9_0 gnd vdd FILL
XFILL_5_DFFPOSX1_214 gnd vdd FILL
XFILL_5_DFFPOSX1_225 gnd vdd FILL
XFILL_5_DFFPOSX1_203 gnd vdd FILL
XFILL_5_DFFPOSX1_258 gnd vdd FILL
XFILL_5_DFFPOSX1_247 gnd vdd FILL
XFILL_5_DFFPOSX1_236 gnd vdd FILL
XFILL_5_DFFPOSX1_269 gnd vdd FILL
XFILL_0_OAI21X1_51 gnd vdd FILL
XFILL_0_OAI21X1_40 gnd vdd FILL
XOAI21X1_1711 INVX2_117/Y BUFX4_301/Y OAI21X1_1711/C gnd DFFPOSX1_68/D vdd OAI21X1
XFILL_0_OAI21X1_62 gnd vdd FILL
XFILL_0_OAI21X1_84 gnd vdd FILL
XFILL_0_OAI21X1_73 gnd vdd FILL
XOAI21X1_1700 BUFX4_97/Y OAI21X1_1/A BUFX2_733/A gnd OAI21X1_1701/C vdd OAI21X1
XOAI21X1_1733 INVX2_128/Y BUFX4_296/Y OAI21X1_1733/C gnd DFFPOSX1_79/D vdd OAI21X1
XOAI21X1_1722 BUFX4_173/Y BUFX4_69/Y BUFX2_773/A gnd OAI21X1_1723/C vdd OAI21X1
XFILL_0_OAI21X1_95 gnd vdd FILL
XOAI21X1_1755 INVX2_139/Y BUFX4_292/Y OAI21X1_1755/C gnd DFFPOSX1_90/D vdd OAI21X1
XOAI21X1_1744 OR2X2_20/B BUFX4_55/A BUFX2_754/A gnd OAI21X1_1745/C vdd OAI21X1
XOAI21X1_1766 BUFX4_179/Y BUFX4_42/Y BUFX2_766/A gnd OAI21X1_1767/C vdd OAI21X1
XOAI21X1_1788 BUFX4_380/Y INVX2_160/Y NAND2X1_729/Y gnd OAI21X1_1788/Y vdd OAI21X1
XOAI21X1_1799 BUFX4_363/Y INVX2_171/Y NAND2X1_740/Y gnd OAI21X1_1799/Y vdd OAI21X1
XFILL_0_OAI21X1_711 gnd vdd FILL
XFILL_0_OAI21X1_722 gnd vdd FILL
XOAI21X1_1777 BUFX4_365/Y INVX2_149/Y NAND2X1_718/Y gnd OAI21X1_1777/Y vdd OAI21X1
XFILL_0_OAI21X1_700 gnd vdd FILL
XFILL_1_OAI21X1_915 gnd vdd FILL
XFILL_1_OAI21X1_937 gnd vdd FILL
XFILL_0_OAI21X1_744 gnd vdd FILL
XFILL_0_OAI21X1_766 gnd vdd FILL
XFILL_0_OAI21X1_733 gnd vdd FILL
XFILL_0_OAI21X1_755 gnd vdd FILL
XFILL_1_OAI21X1_904 gnd vdd FILL
XFILL_1_OAI21X1_926 gnd vdd FILL
XFILL_1_OAI21X1_948 gnd vdd FILL
XFILL_0_OAI21X1_799 gnd vdd FILL
XFILL_0_OAI21X1_777 gnd vdd FILL
XFILL_0_OAI21X1_788 gnd vdd FILL
XFILL_1_OAI21X1_959 gnd vdd FILL
XFILL_13_17_0 gnd vdd FILL
XFILL_2_NAND3X1_27 gnd vdd FILL
XFILL_0_OAI21X1_1532 gnd vdd FILL
XFILL_0_OAI21X1_1521 gnd vdd FILL
XFILL_0_NAND2X1_750 gnd vdd FILL
XFILL_0_OAI21X1_1510 gnd vdd FILL
XFILL_0_OAI21X1_1543 gnd vdd FILL
XFILL_0_NAND2X1_761 gnd vdd FILL
XFILL_24_9_0 gnd vdd FILL
XFILL_0_OAI21X1_1576 gnd vdd FILL
XFILL_0_OAI21X1_1565 gnd vdd FILL
XFILL_0_OAI21X1_1554 gnd vdd FILL
XFILL_0_OAI21X1_1598 gnd vdd FILL
XFILL_0_OAI21X1_1587 gnd vdd FILL
XFILL_5_DFFPOSX1_770 gnd vdd FILL
XFILL_5_DFFPOSX1_781 gnd vdd FILL
XFILL_5_DFFPOSX1_792 gnd vdd FILL
XFILL_0_BUFX2_509 gnd vdd FILL
XFILL_18_16_0 gnd vdd FILL
XBUFX4_128 BUFX4_14/Y gnd BUFX4_128/Y vdd BUFX4
XBUFX4_106 BUFX4_4/A gnd BUFX4_106/Y vdd BUFX4
XBUFX4_117 INVX8_4/Y gnd BUFX4_381/A vdd BUFX4
XFILL_31_18_0 gnd vdd FILL
XFILL_4_DFFPOSX1_382 gnd vdd FILL
XFILL_0_INVX1_28 gnd vdd FILL
XFILL_0_INVX1_17 gnd vdd FILL
XFILL_0_INVX1_39 gnd vdd FILL
XFILL_4_DFFPOSX1_360 gnd vdd FILL
XFILL_4_DFFPOSX1_371 gnd vdd FILL
XBUFX4_139 BUFX4_16/Y gnd BUFX4_139/Y vdd BUFX4
XFILL_2_DFFPOSX1_1030 gnd vdd FILL
XFILL_4_DFFPOSX1_393 gnd vdd FILL
XFILL_1_AND2X2_9 gnd vdd FILL
XFILL_0_OAI22X1_1 gnd vdd FILL
XFILL_15_9_0 gnd vdd FILL
XFILL_1_BUFX2_250 gnd vdd FILL
XFILL_1_BUFX2_283 gnd vdd FILL
XFILL_1_BUFX2_294 gnd vdd FILL
XOAI21X1_1007 BUFX4_296/Y INVX1_158/Y OAI21X1_1007/C gnd OAI21X1_1007/Y vdd OAI21X1
XOAI21X1_1018 BUFX4_125/Y BUFX4_81/A BUFX2_373/A gnd OAI21X1_1019/C vdd OAI21X1
XFILL_1_OAI21X1_1205 gnd vdd FILL
XOAI21X1_1029 BUFX4_291/Y INVX1_169/Y OAI21X1_1029/C gnd OAI21X1_1029/Y vdd OAI21X1
XFILL_1_OAI21X1_1227 gnd vdd FILL
XFILL_1_OAI21X1_1216 gnd vdd FILL
XFILL_1_OAI21X1_1238 gnd vdd FILL
XFILL_1_DFFPOSX1_806 gnd vdd FILL
XDFFPOSX1_608 BUFX2_642/A CLKBUF1_24/Y OAI21X1_834/Y gnd vdd DFFPOSX1
XDFFPOSX1_619 INVX1_48/A CLKBUF1_6/Y OAI21X1_847/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1249 gnd vdd FILL
XFILL_1_DFFPOSX1_839 gnd vdd FILL
XFILL_1_DFFPOSX1_817 gnd vdd FILL
XFILL_1_DFFPOSX1_828 gnd vdd FILL
XFILL_6_DFFPOSX1_410 gnd vdd FILL
XFILL_6_DFFPOSX1_421 gnd vdd FILL
XFILL_6_DFFPOSX1_432 gnd vdd FILL
XFILL_36_17_0 gnd vdd FILL
XFILL_1_1 gnd vdd FILL
XFILL_36_0_1 gnd vdd FILL
XFILL_1_NAND2X1_239 gnd vdd FILL
XFILL_1_NAND3X1_2 gnd vdd FILL
XFILL_1_NAND2X1_206 gnd vdd FILL
XFILL_0_DFFPOSX1_418 gnd vdd FILL
XFILL_0_DFFPOSX1_407 gnd vdd FILL
XFILL_0_DFFPOSX1_429 gnd vdd FILL
XFILL_5_DFFPOSX1_1001 gnd vdd FILL
XFILL_5_DFFPOSX1_1012 gnd vdd FILL
XFILL_5_DFFPOSX1_1023 gnd vdd FILL
XDFFPOSX1_12 BUFX2_711/A CLKBUF1_42/Y DFFPOSX1_12/D gnd vdd DFFPOSX1
XDFFPOSX1_45 BUFX2_744/A CLKBUF1_42/Y DFFPOSX1_45/D gnd vdd DFFPOSX1
XOAI21X1_1530 AOI21X1_62/Y OAI21X1_1530/B OAI21X1_1530/C gnd OAI21X1_1530/Y vdd OAI21X1
XOAI21X1_1541 OR2X2_21/A INVX1_196/A BUFX4_286/Y gnd OAI21X1_1542/B vdd OAI21X1
XDFFPOSX1_23 BUFX2_692/A CLKBUF1_92/Y DFFPOSX1_23/D gnd vdd DFFPOSX1
XDFFPOSX1_34 BUFX2_705/A CLKBUF1_75/Y DFFPOSX1_34/D gnd vdd DFFPOSX1
XFILL_0_BUFX4_380 gnd vdd FILL
XDFFPOSX1_78 BUFX2_747/A CLKBUF1_8/Y DFFPOSX1_78/D gnd vdd DFFPOSX1
XDFFPOSX1_56 BUFX2_726/A CLKBUF1_67/Y DFFPOSX1_56/D gnd vdd DFFPOSX1
XOAI21X1_1574 XNOR2X1_104/Y BUFX4_297/Y OAI21X1_1574/C gnd OAI21X1_1574/Y vdd OAI21X1
XFILL_1_OAI21X1_1761 gnd vdd FILL
XOAI21X1_1563 NOR2X1_232/Y OAI21X1_1563/B OAI21X1_1563/C gnd OAI21X1_1563/Y vdd OAI21X1
XFILL_1_OAI21X1_1750 gnd vdd FILL
XDFFPOSX1_67 BUFX2_738/A CLKBUF1_66/Y DFFPOSX1_67/D gnd vdd DFFPOSX1
XOAI21X1_1552 NOR2X1_230/Y OAI21X1_1552/B OAI21X1_1552/C gnd OAI21X1_1552/Y vdd OAI21X1
XOAI21X1_1596 BUFX4_380/Y INVX2_132/Y NAND2X1_665/Y gnd OAI21X1_1596/Y vdd OAI21X1
XDFFPOSX1_89 BUFX2_759/A CLKBUF1_64/Y DFFPOSX1_89/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1783 gnd vdd FILL
XFILL_1_OAI21X1_712 gnd vdd FILL
XOAI21X1_1585 BUFX4_367/Y INVX2_121/Y NAND2X1_654/Y gnd OAI21X1_1585/Y vdd OAI21X1
XFILL_1_OAI21X1_701 gnd vdd FILL
XFILL_1_OAI21X1_1794 gnd vdd FILL
XFILL_1_OAI21X1_1772 gnd vdd FILL
XFILL_0_OAI21X1_530 gnd vdd FILL
XFILL_1_OAI21X1_745 gnd vdd FILL
XFILL_1_OAI21X1_734 gnd vdd FILL
XFILL_1_OAI21X1_723 gnd vdd FILL
XFILL_0_OAI21X1_541 gnd vdd FILL
XFILL_0_OAI21X1_552 gnd vdd FILL
XFILL_0_OAI21X1_563 gnd vdd FILL
XFILL_0_OAI21X1_574 gnd vdd FILL
XFILL_2_OAI21X1_949 gnd vdd FILL
XFILL_1_OAI21X1_756 gnd vdd FILL
XFILL_2_OAI21X1_938 gnd vdd FILL
XFILL_1_OAI21X1_767 gnd vdd FILL
XFILL_0_OAI21X1_596 gnd vdd FILL
XFILL_1_OAI21X1_778 gnd vdd FILL
XFILL_0_OAI21X1_585 gnd vdd FILL
XFILL_1_OAI21X1_789 gnd vdd FILL
XFILL_0_CLKBUF1_30 gnd vdd FILL
XFILL_27_0_1 gnd vdd FILL
XFILL_0_CLKBUF1_63 gnd vdd FILL
XFILL_0_CLKBUF1_41 gnd vdd FILL
XFILL_2_0_1 gnd vdd FILL
XFILL_0_CLKBUF1_52 gnd vdd FILL
XFILL_0_CLKBUF1_74 gnd vdd FILL
XFILL_0_CLKBUF1_96 gnd vdd FILL
XFILL_0_CLKBUF1_85 gnd vdd FILL
XFILL_0_OAI21X1_1340 gnd vdd FILL
XFILL_0_OAI21X1_1351 gnd vdd FILL
XFILL_0_NAND2X1_580 gnd vdd FILL
XFILL_0_OAI21X1_1384 gnd vdd FILL
XFILL_1_NAND2X1_762 gnd vdd FILL
XFILL_0_NAND2X1_591 gnd vdd FILL
XFILL_0_DFFPOSX1_952 gnd vdd FILL
XFILL_0_DFFPOSX1_941 gnd vdd FILL
XFILL_0_OAI21X1_1373 gnd vdd FILL
XFILL_0_DFFPOSX1_930 gnd vdd FILL
XFILL_0_OAI21X1_1362 gnd vdd FILL
XFILL_0_DFFPOSX1_985 gnd vdd FILL
XFILL_0_DFFPOSX1_963 gnd vdd FILL
XFILL_0_OAI21X1_1395 gnd vdd FILL
XFILL_0_DFFPOSX1_974 gnd vdd FILL
XFILL_0_DFFPOSX1_996 gnd vdd FILL
XFILL_0_OR2X2_2 gnd vdd FILL
XINVX2_117 bundlePid_i[31] gnd INVX2_117/Y vdd INVX2
XFILL_0_BUFX2_306 gnd vdd FILL
XFILL_0_BUFX2_339 gnd vdd FILL
XFILL_0_BUFX2_328 gnd vdd FILL
XINVX2_128 bundlePid_i[20] gnd INVX2_128/Y vdd INVX2
XINVX2_106 INVX2_106/A gnd INVX2_106/Y vdd INVX2
XFILL_0_BUFX2_317 gnd vdd FILL
XINVX2_139 bundlePid_i[9] gnd INVX2_139/Y vdd INVX2
XFILL_20_15_1 gnd vdd FILL
XFILL_4_DFFPOSX1_190 gnd vdd FILL
XFILL_18_0_1 gnd vdd FILL
XFILL_2_NOR3X1_12 gnd vdd FILL
XFILL_2_OAI21X1_1478 gnd vdd FILL
XFILL_0_INVX1_4 gnd vdd FILL
XFILL_30_7_0 gnd vdd FILL
XFILL_25_14_1 gnd vdd FILL
XFILL_1_NAND3X1_13 gnd vdd FILL
XFILL_1_NAND3X1_46 gnd vdd FILL
XFILL_1_NAND3X1_35 gnd vdd FILL
XFILL_1_NAND3X1_24 gnd vdd FILL
XFILL_1_OAI21X1_1002 gnd vdd FILL
XFILL_1_OAI21X1_1013 gnd vdd FILL
XFILL_1_OAI21X1_1046 gnd vdd FILL
XDFFPOSX1_416 BUFX2_450/A CLKBUF1_19/Y OAI21X1_388/Y gnd vdd DFFPOSX1
XDFFPOSX1_405 BUFX2_437/A CLKBUF1_100/Y OAI21X1_377/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_851 gnd vdd FILL
XFILL_0_BUFX2_840 gnd vdd FILL
XFILL_1_NAND3X1_57 gnd vdd FILL
XFILL_1_DFFPOSX1_603 gnd vdd FILL
XFILL_1_NAND3X1_68 gnd vdd FILL
XDFFPOSX1_427 BUFX2_518/A CLKBUF1_75/Y OAI21X1_409/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1024 gnd vdd FILL
XFILL_1_DFFPOSX1_614 gnd vdd FILL
XDFFPOSX1_438 BUFX2_467/A CLKBUF1_24/Y OAI21X1_427/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1035 gnd vdd FILL
XFILL_0_BUFX2_884 gnd vdd FILL
XFILL_1_DFFPOSX1_636 gnd vdd FILL
XFILL_0_BUFX2_873 gnd vdd FILL
XINVX1_150 bundle_i[118] gnd INVX1_150/Y vdd INVX1
XFILL_1_OAI21X1_1068 gnd vdd FILL
XFILL_1_OAI21X1_1079 gnd vdd FILL
XINVX1_161 bundle_i[107] gnd INVX1_161/Y vdd INVX1
XFILL_1_DFFPOSX1_647 gnd vdd FILL
XFILL_1_DFFPOSX1_625 gnd vdd FILL
XFILL_0_BUFX2_862 gnd vdd FILL
XDFFPOSX1_449 BUFX2_479/A CLKBUF1_33/Y OAI21X1_444/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1057 gnd vdd FILL
XINVX1_183 INVX1_183/A gnd INVX1_183/Y vdd INVX1
XINVX1_194 INVX1_194/A gnd INVX1_194/Y vdd INVX1
XFILL_0_BUFX2_895 gnd vdd FILL
XFILL_1_DFFPOSX1_658 gnd vdd FILL
XFILL_1_DFFPOSX1_669 gnd vdd FILL
XNAND2X1_508 BUFX2_79/A BUFX4_192/Y gnd NAND2X1_508/Y vdd NAND2X1
XINVX1_172 bundle_i[96] gnd INVX1_172/Y vdd INVX1
XNAND2X1_519 NOR2X1_140/Y NOR2X1_142/Y gnd INVX1_189/A vdd NAND2X1
XFILL_6_DFFPOSX1_273 gnd vdd FILL
XFILL_6_DFFPOSX1_284 gnd vdd FILL
XFILL_6_DFFPOSX1_295 gnd vdd FILL
XFILL_38_8_0 gnd vdd FILL
XFILL_0_INVX2_60 gnd vdd FILL
XFILL_0_INVX2_82 gnd vdd FILL
XFILL_0_INVX2_71 gnd vdd FILL
XFILL_0_INVX2_93 gnd vdd FILL
XFILL_1_NOR3X1_2 gnd vdd FILL
XFILL_0_15_1 gnd vdd FILL
XFILL_0_DFFPOSX1_204 gnd vdd FILL
XFILL_0_DFFPOSX1_237 gnd vdd FILL
XFILL_0_DFFPOSX1_248 gnd vdd FILL
XFILL_0_DFFPOSX1_215 gnd vdd FILL
XFILL_0_DFFPOSX1_226 gnd vdd FILL
XFILL_0_DFFPOSX1_259 gnd vdd FILL
XFILL_21_7_0 gnd vdd FILL
XFILL_3_DFFPOSX1_719 gnd vdd FILL
XFILL_3_DFFPOSX1_708 gnd vdd FILL
XFILL_3_CLKBUF1_29 gnd vdd FILL
XFILL_3_CLKBUF1_18 gnd vdd FILL
XDFFPOSX1_950 BUFX2_199/A CLKBUF1_70/Y OAI21X1_1427/Y gnd vdd DFFPOSX1
XOAI21X1_1382 BUFX4_99/Y BUFX4_360/Y BUFX2_189/A gnd OAI21X1_1383/C vdd OAI21X1
XOAI21X1_1360 NOR2X1_209/Y OAI21X1_1360/B OAI21X1_1360/C gnd OAI21X1_1360/Y vdd OAI21X1
XOAI21X1_1371 OAI21X1_1371/A BUFX4_160/Y OAI21X1_1371/C gnd OAI21X1_1371/Y vdd OAI21X1
XFILL_1_OAI21X1_1591 gnd vdd FILL
XOAI21X1_1393 NAND2X1_591/B bundleAddress_i[61] OAI21X1_1393/C gnd OAI21X1_1395/A
+ vdd OAI21X1
XDFFPOSX1_961 BUFX2_211/A CLKBUF1_55/Y OAI21X1_1457/Y gnd vdd DFFPOSX1
XDFFPOSX1_983 BUFX2_235/A CLKBUF1_30/Y OAI21X1_1527/Y gnd vdd DFFPOSX1
XDFFPOSX1_994 BUFX2_247/A CLKBUF1_36/Y OAI21X1_1560/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1580 gnd vdd FILL
XDFFPOSX1_972 BUFX2_223/A CLKBUF1_85/Y OAI21X1_1492/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_520 gnd vdd FILL
XFILL_1_NOR2X1_103 gnd vdd FILL
XFILL_1_NOR2X1_125 gnd vdd FILL
XFILL_1_NOR2X1_147 gnd vdd FILL
XFILL_0_OAI21X1_371 gnd vdd FILL
XFILL_1_NOR2X1_136 gnd vdd FILL
XFILL_1_OAI21X1_553 gnd vdd FILL
XFILL_0_OAI21X1_360 gnd vdd FILL
XFILL_0_OAI21X1_382 gnd vdd FILL
XFILL_1_OAI21X1_542 gnd vdd FILL
XFILL_1_OAI21X1_531 gnd vdd FILL
XFILL_2_OAI21X1_768 gnd vdd FILL
XFILL_1_OAI21X1_597 gnd vdd FILL
XFILL_1_OAI21X1_575 gnd vdd FILL
XFILL_0_OAI21X1_393 gnd vdd FILL
XFILL_1_NOR2X1_169 gnd vdd FILL
XFILL_1_OAI21X1_564 gnd vdd FILL
XFILL_1_OAI21X1_586 gnd vdd FILL
XFILL_29_8_0 gnd vdd FILL
XFILL_5_14_1 gnd vdd FILL
XFILL_2_DFFPOSX1_309 gnd vdd FILL
XBUFX2_418 BUFX2_418/A gnd majID1_o[32] vdd BUFX2
XBUFX2_407 BUFX2_407/A gnd majID1_o[42] vdd BUFX2
XFILL_4_8_0 gnd vdd FILL
XBUFX2_429 BUFX2_429/A gnd majID1_o[22] vdd BUFX2
XFILL_1_BUFX4_312 gnd vdd FILL
XFILL_1_BUFX4_301 gnd vdd FILL
XFILL_1_NAND2X1_592 gnd vdd FILL
XFILL_0_OAI21X1_1170 gnd vdd FILL
XFILL_1_BUFX4_356 gnd vdd FILL
XFILL_0_DFFPOSX1_760 gnd vdd FILL
XFILL_1_BUFX4_323 gnd vdd FILL
XFILL_1_BUFX4_334 gnd vdd FILL
XFILL_1_NAND2X1_581 gnd vdd FILL
XFILL_0_OAI21X1_1181 gnd vdd FILL
XFILL_1_BUFX4_345 gnd vdd FILL
XFILL_0_OAI21X1_1192 gnd vdd FILL
XFILL_1_NAND2X1_570 gnd vdd FILL
XFILL_0_DFFPOSX1_771 gnd vdd FILL
XFILL_0_DFFPOSX1_793 gnd vdd FILL
XFILL_1_BUFX4_378 gnd vdd FILL
XFILL_1_BUFX4_367 gnd vdd FILL
XFILL_12_7_0 gnd vdd FILL
XFILL_0_DFFPOSX1_782 gnd vdd FILL
XFILL_2_OAI21X1_58 gnd vdd FILL
XFILL_0_BUFX2_103 gnd vdd FILL
XFILL_0_BUFX2_136 gnd vdd FILL
XFILL_0_BUFX2_125 gnd vdd FILL
XFILL_0_BUFX2_114 gnd vdd FILL
XFILL_0_BUFX2_147 gnd vdd FILL
XFILL_0_BUFX2_169 gnd vdd FILL
XFILL_0_BUFX2_158 gnd vdd FILL
XFILL_1_NAND2X1_90 gnd vdd FILL
XFILL_2_DFFPOSX1_821 gnd vdd FILL
XFILL_2_DFFPOSX1_810 gnd vdd FILL
XFILL_2_DFFPOSX1_832 gnd vdd FILL
XBUFX2_930 BUFX2_930/A gnd tid3_o[32] vdd BUFX2
XBUFX2_963 BUFX2_963/A gnd tid3_o[2] vdd BUFX2
XFILL_2_DFFPOSX1_854 gnd vdd FILL
XBUFX2_952 BUFX2_952/A gnd tid3_o[12] vdd BUFX2
XFILL_2_DFFPOSX1_843 gnd vdd FILL
XBUFX2_974 BUFX2_974/A gnd tid4_o[50] vdd BUFX2
XBUFX2_941 BUFX2_941/A gnd tid3_o[22] vdd BUFX2
XFILL_2_DFFPOSX1_865 gnd vdd FILL
XBUFX2_996 BUFX2_996/A gnd tid4_o[30] vdd BUFX2
XFILL_2_DFFPOSX1_887 gnd vdd FILL
XFILL_2_DFFPOSX1_876 gnd vdd FILL
XBUFX2_985 BUFX2_985/A gnd tid4_o[40] vdd BUFX2
XFILL_2_DFFPOSX1_898 gnd vdd FILL
XDFFPOSX1_202 BUFX2_873/A CLKBUF1_99/Y OAI21X1_46/Y gnd vdd DFFPOSX1
XDFFPOSX1_213 BUFX2_885/A CLKBUF1_67/Y OAI21X1_57/Y gnd vdd DFFPOSX1
XBUFX4_8 BUFX4_8/A gnd BUFX4_8/Y vdd BUFX4
XDFFPOSX1_246 BUFX2_915/A CLKBUF1_27/Y OAI21X1_109/Y gnd vdd DFFPOSX1
XDFFPOSX1_235 BUFX2_966/A CLKBUF1_26/Y OAI21X1_87/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_422 gnd vdd FILL
XFILL_1_DFFPOSX1_400 gnd vdd FILL
XFILL_1_DFFPOSX1_411 gnd vdd FILL
XDFFPOSX1_224 BUFX2_898/A CLKBUF1_52/Y OAI21X1_68/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_670 gnd vdd FILL
XFILL_0_BUFX2_681 gnd vdd FILL
XDFFPOSX1_279 BUFX2_952/A CLKBUF1_38/Y OAI21X1_175/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_692 gnd vdd FILL
XFILL_1_DFFPOSX1_433 gnd vdd FILL
XDFFPOSX1_268 BUFX2_940/A CLKBUF1_2/Y OAI21X1_153/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_466 gnd vdd FILL
XDFFPOSX1_257 BUFX2_927/A CLKBUF1_62/Y OAI21X1_131/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_455 gnd vdd FILL
XFILL_1_DFFPOSX1_444 gnd vdd FILL
XNAND2X1_305 INVX1_43/A NOR2X1_97/Y gnd OAI21X1_648/A vdd NAND2X1
XFILL_1_DFFPOSX1_477 gnd vdd FILL
XNAND2X1_327 bundleStartMajId_i[25] AND2X2_21/A gnd XNOR2X1_51/A vdd NAND2X1
XFILL_1_DFFPOSX1_499 gnd vdd FILL
XNAND2X1_316 OAI21X1_704/Y INVX1_36/A gnd OAI21X1_706/A vdd NAND2X1
XFILL_1_DFFPOSX1_488 gnd vdd FILL
XNAND2X1_349 BUFX4_267/Y bundle_i[20] gnd OAI21X1_855/C vdd NAND2X1
XFILL_4_DFFPOSX1_904 gnd vdd FILL
XNAND2X1_338 BUFX4_264/Y bundle_i[31] gnd OAI21X1_844/C vdd NAND2X1
XFILL_4_DFFPOSX1_937 gnd vdd FILL
XFILL_4_DFFPOSX1_915 gnd vdd FILL
XFILL_4_DFFPOSX1_926 gnd vdd FILL
XFILL_4_DFFPOSX1_948 gnd vdd FILL
XNOR3X1_12 INVX4_44/Y NOR3X1_12/B NOR3X1_14/C gnd NOR3X1_12/Y vdd NOR3X1
XFILL_4_DFFPOSX1_959 gnd vdd FILL
XFILL_10_15_0 gnd vdd FILL
XFILL_0_XNOR2X1_4 gnd vdd FILL
XFILL_1_BUFX2_816 gnd vdd FILL
XFILL_1_BUFX2_827 gnd vdd FILL
XOAI21X1_800 BUFX4_155/Y BUFX4_57/Y BUFX2_629/A gnd OAI21X1_801/C vdd OAI21X1
XINVX4_8 bundleStartMajId_i[42] gnd INVX4_8/Y vdd INVX4
XOAI21X1_822 NOR3X1_8/C NOR3X1_4/A INVX2_37/Y gnd OAI21X1_822/Y vdd OAI21X1
XOAI21X1_811 INVX2_53/Y OR2X2_13/B OAI21X1_811/C gnd OAI21X1_813/A vdd OAI21X1
XFILL_1_BUFX2_838 gnd vdd FILL
XOAI21X1_833 BUFX4_177/Y BUFX4_74/Y BUFX2_642/A gnd OAI21X1_834/C vdd OAI21X1
XOAI21X1_855 INVX1_56/Y BUFX4_267/Y OAI21X1_855/C gnd OAI21X1_855/Y vdd OAI21X1
XFILL_3_DFFPOSX1_516 gnd vdd FILL
XFILL_3_DFFPOSX1_527 gnd vdd FILL
XFILL_3_DFFPOSX1_538 gnd vdd FILL
XOAI21X1_866 INVX1_67/Y BUFX4_261/Y OAI21X1_866/C gnd OAI21X1_866/Y vdd OAI21X1
XOAI21X1_844 INVX1_45/Y BUFX4_264/Y OAI21X1_844/C gnd OAI21X1_844/Y vdd OAI21X1
XFILL_3_DFFPOSX1_505 gnd vdd FILL
XOAI21X1_888 INVX1_89/Y BUFX4_193/Y OAI21X1_888/C gnd OAI21X1_888/Y vdd OAI21X1
XOAI21X1_877 INVX1_78/Y BUFX4_211/Y OAI21X1_877/C gnd OAI21X1_877/Y vdd OAI21X1
XOAI21X1_899 INVX1_100/Y BUFX4_232/Y OAI21X1_899/C gnd OAI21X1_899/Y vdd OAI21X1
XFILL_3_DFFPOSX1_549 gnd vdd FILL
XOAI21X1_1190 NAND3X1_48/Y INVX4_45/Y BUFX4_242/Y gnd OAI21X1_1191/A vdd OAI21X1
XDFFPOSX1_791 BUFX2_43/A CLKBUF1_30/Y OAI21X1_1083/Y gnd vdd DFFPOSX1
XDFFPOSX1_780 BUFX2_31/A CLKBUF1_28/Y OAI21X1_1072/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_350 gnd vdd FILL
XFILL_0_OAI21X1_190 gnd vdd FILL
XFILL_1_OAI21X1_361 gnd vdd FILL
XFILL_2_OAI21X1_576 gnd vdd FILL
XFILL_1_OAI21X1_372 gnd vdd FILL
XFILL_1_OAI21X1_394 gnd vdd FILL
XFILL_1_CLKBUF1_4 gnd vdd FILL
XFILL_1_OAI21X1_383 gnd vdd FILL
XFILL_0_NAND3X1_10 gnd vdd FILL
XFILL_15_14_0 gnd vdd FILL
XFILL_2_OAI21X1_598 gnd vdd FILL
XFILL_2_DFFPOSX1_117 gnd vdd FILL
XFILL_0_NAND3X1_54 gnd vdd FILL
XFILL_2_DFFPOSX1_106 gnd vdd FILL
XFILL_0_NAND3X1_32 gnd vdd FILL
XBUFX2_215 BUFX2_215/A gnd addr4_o[34] vdd BUFX2
XFILL_0_NAND3X1_21 gnd vdd FILL
XBUFX2_204 BUFX2_204/A gnd addr4_o[44] vdd BUFX2
XFILL_2_DFFPOSX1_128 gnd vdd FILL
XBUFX2_226 BUFX2_226/A gnd addr4_o[24] vdd BUFX2
XFILL_0_NAND3X1_43 gnd vdd FILL
XBUFX2_237 BUFX2_237/A gnd addr4_o[14] vdd BUFX2
XFILL_2_DFFPOSX1_139 gnd vdd FILL
XBUFX2_248 BUFX2_248/A gnd addr4_o[4] vdd BUFX2
XFILL_0_NAND3X1_65 gnd vdd FILL
XBUFX2_259 BUFX2_259/A gnd enable3_o vdd BUFX2
XFILL_1_BUFX4_120 gnd vdd FILL
XFILL_1_BUFX4_164 gnd vdd FILL
XFILL_1_BUFX4_142 gnd vdd FILL
XFILL_1_BUFX4_153 gnd vdd FILL
XFILL_1_BUFX4_131 gnd vdd FILL
XFILL_1_BUFX4_197 gnd vdd FILL
XFILL_1_BUFX4_175 gnd vdd FILL
XFILL_0_DFFPOSX1_590 gnd vdd FILL
XFILL_1_BUFX4_186 gnd vdd FILL
XFILL_33_15_0 gnd vdd FILL
XFILL_2_CLKBUF1_26 gnd vdd FILL
XFILL_2_CLKBUF1_48 gnd vdd FILL
XFILL_2_CLKBUF1_37 gnd vdd FILL
XFILL_2_CLKBUF1_15 gnd vdd FILL
XFILL_35_6_0 gnd vdd FILL
XFILL_2_DFFPOSX1_640 gnd vdd FILL
XFILL_2_CLKBUF1_59 gnd vdd FILL
XFILL_2_DFFPOSX1_662 gnd vdd FILL
XBUFX2_760 BUFX2_760/A gnd pid4_o[9] vdd BUFX2
XFILL_2_DFFPOSX1_651 gnd vdd FILL
XBUFX2_771 BUFX2_771/A gnd pid4_o[27] vdd BUFX2
XFILL_2_DFFPOSX1_673 gnd vdd FILL
XBUFX2_782 BUFX2_782/A gnd tid1_o[50] vdd BUFX2
XFILL_2_DFFPOSX1_684 gnd vdd FILL
XFILL_0_NOR2X1_100 gnd vdd FILL
XFILL_0_NOR2X1_122 gnd vdd FILL
XBUFX2_793 BUFX2_793/A gnd tid1_o[40] vdd BUFX2
XFILL_0_NOR2X1_111 gnd vdd FILL
XFILL_2_DFFPOSX1_695 gnd vdd FILL
XFILL_0_NOR2X1_133 gnd vdd FILL
XFILL_0_NOR2X1_144 gnd vdd FILL
XFILL_0_NOR2X1_155 gnd vdd FILL
XOAI21X1_107 BUFX4_132/Y INVX2_163/Y OAI21X1_107/C gnd OAI21X1_107/Y vdd OAI21X1
XOAI21X1_118 BUFX4_11/A BUFX4_322/Y BUFX2_921/A gnd OAI21X1_119/C vdd OAI21X1
XFILL_0_NOR2X1_177 gnd vdd FILL
XFILL_0_NOR2X1_166 gnd vdd FILL
XFILL_0_NOR2X1_188 gnd vdd FILL
XOAI21X1_129 BUFX4_158/Y INVX2_174/Y OAI21X1_129/C gnd OAI21X1_129/Y vdd OAI21X1
XFILL_0_DFFPOSX1_1018 gnd vdd FILL
XFILL_0_DFFPOSX1_1007 gnd vdd FILL
XFILL_0_NOR2X1_199 gnd vdd FILL
XFILL_0_DFFPOSX1_1029 gnd vdd FILL
XBUFX2_5 BUFX2_5/A gnd addr1_o[51] vdd BUFX2
XFILL_1_DFFPOSX1_230 gnd vdd FILL
XFILL_1_DFFPOSX1_241 gnd vdd FILL
XFILL_38_14_0 gnd vdd FILL
XFILL_1_DFFPOSX1_252 gnd vdd FILL
XFILL_1_DFFPOSX1_263 gnd vdd FILL
XFILL_1_DFFPOSX1_274 gnd vdd FILL
XFILL_1_DFFPOSX1_296 gnd vdd FILL
XFILL_1_DFFPOSX1_285 gnd vdd FILL
XNAND2X1_113 BUFX2_429/A BUFX4_362/Y gnd OAI21X1_369/C vdd NAND2X1
XNAND2X1_124 BUFX2_441/A BUFX4_358/Y gnd OAI21X1_380/C vdd NAND2X1
XNAND2X1_102 BUFX2_417/A BUFX4_319/Y gnd OAI21X1_358/C vdd NAND2X1
XNAND2X1_135 BUFX2_453/A BUFX4_373/Y gnd OAI21X1_391/C vdd NAND2X1
XFILL_4_DFFPOSX1_701 gnd vdd FILL
XNAND2X1_168 bundleStartMajId_i[47] NOR2X1_11/Y gnd INVX1_10/A vdd NAND2X1
XFILL_4_DFFPOSX1_712 gnd vdd FILL
XNAND2X1_157 INVX1_9/Y NOR2X1_5/Y gnd XNOR2X1_2/A vdd NAND2X1
XNAND2X1_146 BUFX2_502/A BUFX4_222/Y gnd OAI21X1_404/C vdd NAND2X1
XFILL_1_OAI21X1_22 gnd vdd FILL
XFILL_4_DFFPOSX1_756 gnd vdd FILL
XFILL_1_OAI21X1_33 gnd vdd FILL
XFILL_4_DFFPOSX1_745 gnd vdd FILL
XFILL_4_DFFPOSX1_734 gnd vdd FILL
XFILL_4_DFFPOSX1_723 gnd vdd FILL
XNAND2X1_179 BUFX2_470/A BUFX4_194/Y gnd OAI21X1_431/C vdd NAND2X1
XFILL_1_OAI21X1_11 gnd vdd FILL
XFILL_1_OAI21X1_55 gnd vdd FILL
XFILL_1_OAI21X1_44 gnd vdd FILL
XFILL_4_DFFPOSX1_789 gnd vdd FILL
XFILL_4_DFFPOSX1_778 gnd vdd FILL
XFILL_1_OAI21X1_66 gnd vdd FILL
XFILL_4_DFFPOSX1_767 gnd vdd FILL
XFILL_26_6_0 gnd vdd FILL
XFILL_1_OAI21X1_99 gnd vdd FILL
XFILL_1_OAI21X1_77 gnd vdd FILL
XFILL_1_OAI21X1_88 gnd vdd FILL
XFILL_1_6_0 gnd vdd FILL
XNOR2X1_190 OR2X2_17/Y NOR3X1_18/C gnd NOR2X1_190/Y vdd NOR2X1
XFILL_0_DFFPOSX1_9 gnd vdd FILL
XFILL_1_BUFX2_613 gnd vdd FILL
XFILL_1_BUFX2_624 gnd vdd FILL
XINVX2_5 bundleTid_i[2] gnd INVX2_5/Y vdd INVX2
XFILL_1_BUFX2_635 gnd vdd FILL
XFILL_1_BUFX2_679 gnd vdd FILL
XOAI21X1_641 BUFX4_251/Y BUFX4_328/Y BUFX2_574/A gnd OAI21X1_643/C vdd OAI21X1
XFILL_3_DFFPOSX1_313 gnd vdd FILL
XOAI21X1_630 XNOR2X1_38/Y BUFX4_145/Y OAI21X1_630/C gnd OAI21X1_630/Y vdd OAI21X1
XFILL_0_BUFX4_209 gnd vdd FILL
XFILL_1_BUFX2_668 gnd vdd FILL
XFILL_3_DFFPOSX1_302 gnd vdd FILL
XOAI21X1_652 BUFX4_3/A BUFX4_386/Y BUFX2_579/A gnd OAI21X1_654/C vdd OAI21X1
XFILL_3_DFFPOSX1_346 gnd vdd FILL
XFILL_3_DFFPOSX1_335 gnd vdd FILL
XAOI21X1_5 INVX1_44/A NOR2X1_52/Y bundleStartMajId_i[3] gnd AOI21X1_5/Y vdd AOI21X1
XOAI21X1_663 OAI21X1_663/A bundleStartMajId_i[63] OAI21X1_663/C gnd OAI21X1_665/A
+ vdd OAI21X1
XFILL_3_DFFPOSX1_324 gnd vdd FILL
XOAI21X1_674 BUFX4_173/Y BUFX4_46/Y BUFX2_630/A gnd OAI21X1_675/C vdd OAI21X1
XFILL_3_DFFPOSX1_357 gnd vdd FILL
XFILL_3_DFFPOSX1_368 gnd vdd FILL
XOAI21X1_696 BUFX4_167/Y BUFX4_72/Y BUFX2_590/A gnd OAI21X1_697/C vdd OAI21X1
XFILL_3_DFFPOSX1_379 gnd vdd FILL
XOAI21X1_685 XNOR2X1_41/Y BUFX4_299/Y OAI21X1_685/C gnd OAI21X1_685/Y vdd OAI21X1
XFILL_6_DFFPOSX1_806 gnd vdd FILL
XFILL_6_DFFPOSX1_817 gnd vdd FILL
XFILL_0_INVX4_17 gnd vdd FILL
XFILL_6_DFFPOSX1_828 gnd vdd FILL
XFILL_6_DFFPOSX1_839 gnd vdd FILL
XFILL_0_INVX4_28 gnd vdd FILL
XFILL_0_INVX4_39 gnd vdd FILL
XXNOR2X1_13 INVX1_15/A INVX4_15/Y gnd XNOR2X1_13/Y vdd XNOR2X1
XFILL_9_7_0 gnd vdd FILL
XFILL_1_OAI21X1_180 gnd vdd FILL
XXNOR2X1_57 XNOR2X1_57/A bundleAddress_i[48] gnd XNOR2X1_57/Y vdd XNOR2X1
XXNOR2X1_46 XNOR2X1_46/A INVX4_12/Y gnd XNOR2X1_46/Y vdd XNOR2X1
XXNOR2X1_35 NOR2X1_79/Y bundleStartMajId_i[25] gnd XNOR2X1_35/Y vdd XNOR2X1
XXNOR2X1_24 INVX4_29/Y INVX4_2/Y gnd XNOR2X1_24/Y vdd XNOR2X1
XNAND2X1_691 BUFX2_712/A BUFX4_218/Y gnd NAND2X1_691/Y vdd NAND2X1
XXNOR2X1_79 XNOR2X1_79/A INVX2_71/Y gnd XNOR2X1_79/Y vdd XNOR2X1
XNAND2X1_680 BUFX2_673/A BUFX4_373/Y gnd NAND2X1_680/Y vdd NAND2X1
XFILL_1_OAI21X1_191 gnd vdd FILL
XXNOR2X1_68 XNOR2X1_68/A bundleAddress_i[27] gnd XNOR2X1_68/Y vdd XNOR2X1
XFILL_1_INVX2_197 gnd vdd FILL
XINVX1_92 bundle_i[48] gnd INVX1_92/Y vdd INVX1
XINVX1_70 INVX1_70/A gnd INVX1_70/Y vdd INVX1
XINVX1_81 bundle_i[59] gnd INVX1_81/Y vdd INVX1
XFILL_0_NAND2X1_409 gnd vdd FILL
XBUFX2_23 BUFX2_23/A gnd addr1_o[34] vdd BUFX2
XBUFX2_45 BUFX2_45/A gnd addr1_o[14] vdd BUFX2
XBUFX2_12 BUFX2_12/A gnd addr1_o[44] vdd BUFX2
XBUFX2_34 BUFX2_34/A gnd addr1_o[24] vdd BUFX2
XBUFX2_67 BUFX2_67/A gnd addr2_o[53] vdd BUFX2
XBUFX2_56 BUFX2_56/A gnd addr1_o[4] vdd BUFX2
XFILL_17_6_0 gnd vdd FILL
XBUFX2_78 BUFX2_78/A gnd addr2_o[43] vdd BUFX2
XBUFX2_89 BUFX2_89/A gnd addr2_o[33] vdd BUFX2
XFILL_5_DFFPOSX1_418 gnd vdd FILL
XFILL_5_DFFPOSX1_407 gnd vdd FILL
XFILL_5_DFFPOSX1_429 gnd vdd FILL
XFILL_1_BUFX4_34 gnd vdd FILL
XFILL_1_BUFX4_23 gnd vdd FILL
XFILL_1_BUFX4_45 gnd vdd FILL
XFILL_1_BUFX4_12 gnd vdd FILL
XFILL_1_BUFX4_67 gnd vdd FILL
XFILL_22_12_1 gnd vdd FILL
XFILL_1_BUFX4_56 gnd vdd FILL
XFILL_1_BUFX4_78 gnd vdd FILL
XFILL_1_BUFX4_89 gnd vdd FILL
XFILL_0_OAI21X1_915 gnd vdd FILL
XFILL_3_DFFPOSX1_880 gnd vdd FILL
XFILL_3_DFFPOSX1_891 gnd vdd FILL
XNOR2X1_3 INVX1_7/A NOR2X1_3/B gnd NOR2X1_3/Y vdd NOR2X1
XFILL_0_OAI21X1_904 gnd vdd FILL
XFILL_0_OAI21X1_948 gnd vdd FILL
XFILL_0_OAI21X1_937 gnd vdd FILL
XFILL_0_OAI21X1_926 gnd vdd FILL
XFILL_0_OAI21X1_959 gnd vdd FILL
XFILL_2_BUFX4_118 gnd vdd FILL
XFILL_1_OR2X2_15 gnd vdd FILL
XFILL_0_OAI21X1_1725 gnd vdd FILL
XFILL_0_OAI21X1_1714 gnd vdd FILL
XFILL_0_OAI21X1_1703 gnd vdd FILL
XFILL_0_OAI21X1_1758 gnd vdd FILL
XFILL_0_OAI21X1_1736 gnd vdd FILL
XFILL_2_DFFPOSX1_470 gnd vdd FILL
XFILL_2_DFFPOSX1_481 gnd vdd FILL
XFILL_0_OAI21X1_1747 gnd vdd FILL
XBUFX2_590 BUFX2_590/A gnd majID4_o[50] vdd BUFX2
XFILL_2_DFFPOSX1_492 gnd vdd FILL
XFILL_0_OAI21X1_1769 gnd vdd FILL
XFILL_27_11_1 gnd vdd FILL
XFILL_5_DFFPOSX1_930 gnd vdd FILL
XFILL_5_DFFPOSX1_952 gnd vdd FILL
XFILL_5_DFFPOSX1_941 gnd vdd FILL
XFILL_5_DFFPOSX1_963 gnd vdd FILL
XFILL_5_DFFPOSX1_974 gnd vdd FILL
XAOI21X1_24 bundleStartMajId_i[6] NOR2X1_97/Y bundleStartMajId_i[5] gnd AOI21X1_24/Y
+ vdd AOI21X1
XFILL_5_DFFPOSX1_985 gnd vdd FILL
XAOI21X1_35 bundleStartMajId_i[2] NOR2X1_119/B bundleStartMajId_i[1] gnd AOI21X1_35/Y
+ vdd AOI21X1
XAOI21X1_13 bundleStartMajId_i[22] NOR2X1_84/Y bundleStartMajId_i[21] gnd AOI21X1_13/Y
+ vdd AOI21X1
XFILL_5_DFFPOSX1_996 gnd vdd FILL
XAOI21X1_46 bundleAddress_i[46] NOR2X1_184/Y bundleAddress_i[45] gnd AOI21X1_46/Y
+ vdd AOI21X1
XAOI21X1_57 INVX2_104/A INVX1_215/Y bundleAddress_i[6] gnd AOI21X1_57/Y vdd AOI21X1
XOAI21X1_8 OAI21X1_8/A OAI21X1_8/B OAI21X1_8/C gnd OAI21X1_8/Y vdd OAI21X1
XFILL_4_DFFPOSX1_520 gnd vdd FILL
XFILL_4_DFFPOSX1_531 gnd vdd FILL
XFILL_4_DFFPOSX1_542 gnd vdd FILL
XFILL_4_DFFPOSX1_564 gnd vdd FILL
XFILL_4_DFFPOSX1_553 gnd vdd FILL
XFILL_4_DFFPOSX1_575 gnd vdd FILL
XFILL_4_DFFPOSX1_586 gnd vdd FILL
XFILL_4_DFFPOSX1_597 gnd vdd FILL
XFILL_2_12_1 gnd vdd FILL
XFILL_1_BUFX2_1011 gnd vdd FILL
XFILL_1_BUFX2_1022 gnd vdd FILL
XFILL_1_BUFX2_421 gnd vdd FILL
XFILL_1_BUFX2_432 gnd vdd FILL
XFILL_3_DFFPOSX1_121 gnd vdd FILL
XFILL_1_CLKBUF1_12 gnd vdd FILL
XFILL_1_BUFX2_487 gnd vdd FILL
XFILL_1_BUFX2_476 gnd vdd FILL
XFILL_3_DFFPOSX1_110 gnd vdd FILL
XFILL_1_BUFX2_465 gnd vdd FILL
XFILL_3_DFFPOSX1_154 gnd vdd FILL
XFILL_3_DFFPOSX1_143 gnd vdd FILL
XFILL_1_OAI21X1_1409 gnd vdd FILL
XFILL_1_INVX8_7 gnd vdd FILL
XFILL_1_CLKBUF1_23 gnd vdd FILL
XOAI21X1_493 OAI21X1_493/A NOR3X1_4/B BUFX4_240/Y gnd OAI21X1_494/A vdd OAI21X1
XFILL_1_CLKBUF1_45 gnd vdd FILL
XOAI21X1_460 NOR3X1_2/C INVX4_19/Y INVX4_20/Y gnd OAI21X1_460/Y vdd OAI21X1
XFILL_1_CLKBUF1_34 gnd vdd FILL
XOAI21X1_482 AND2X2_10/Y bundleStartMajId_i[9] BUFX4_240/Y gnd OAI21X1_483/A vdd OAI21X1
XFILL_1_CLKBUF1_56 gnd vdd FILL
XFILL_3_DFFPOSX1_132 gnd vdd FILL
XOAI21X1_471 NOR2X1_40/Y OAI21X1_471/B OAI21X1_471/C gnd OAI21X1_471/Y vdd OAI21X1
XFILL_3_DFFPOSX1_176 gnd vdd FILL
XFILL_3_DFFPOSX1_187 gnd vdd FILL
XFILL_1_CLKBUF1_67 gnd vdd FILL
XFILL_1_CLKBUF1_89 gnd vdd FILL
XFILL_1_CLKBUF1_78 gnd vdd FILL
XFILL_3_DFFPOSX1_165 gnd vdd FILL
XFILL_3_DFFPOSX1_198 gnd vdd FILL
XFILL_6_DFFPOSX1_603 gnd vdd FILL
XFILL_6_DFFPOSX1_614 gnd vdd FILL
XFILL_7_11_1 gnd vdd FILL
XFILL_2_OAI21X1_181 gnd vdd FILL
XFILL_0_NAND2X1_206 gnd vdd FILL
XFILL_0_INVX1_220 gnd vdd FILL
XFILL_0_NAND2X1_239 gnd vdd FILL
XFILL_0_NAND2X1_217 gnd vdd FILL
XFILL_0_NAND2X1_228 gnd vdd FILL
XFILL_33_9_1 gnd vdd FILL
XFILL_32_4_0 gnd vdd FILL
XFILL_5_DFFPOSX1_215 gnd vdd FILL
XFILL_5_DFFPOSX1_226 gnd vdd FILL
XFILL_5_DFFPOSX1_204 gnd vdd FILL
XFILL_5_DFFPOSX1_237 gnd vdd FILL
XFILL_5_DFFPOSX1_248 gnd vdd FILL
XFILL_5_DFFPOSX1_259 gnd vdd FILL
XFILL_0_OAI21X1_41 gnd vdd FILL
XFILL_0_OAI21X1_30 gnd vdd FILL
XFILL_0_OAI21X1_52 gnd vdd FILL
XOAI21X1_1712 BUFX4_132/Y BUFX4_29/Y BUFX2_746/A gnd OAI21X1_1713/C vdd OAI21X1
XOAI21X1_1701 BUFX4_168/Y INVX2_144/Y OAI21X1_1701/C gnd DFFPOSX1_63/D vdd OAI21X1
XFILL_0_OAI21X1_74 gnd vdd FILL
XFILL_0_OAI21X1_63 gnd vdd FILL
XOAI21X1_1723 INVX2_123/Y BUFX4_302/Y OAI21X1_1723/C gnd DFFPOSX1_74/D vdd OAI21X1
XOAI21X1_1756 BUFX4_123/Y BUFX4_60/Y BUFX2_761/A gnd OAI21X1_1757/C vdd OAI21X1
XFILL_0_OAI21X1_96 gnd vdd FILL
XFILL_0_OAI21X1_85 gnd vdd FILL
XOAI21X1_1745 INVX2_134/Y BUFX4_301/Y OAI21X1_1745/C gnd DFFPOSX1_85/D vdd OAI21X1
XOAI21X1_1734 BUFX4_176/Y BUFX4_46/Y BUFX2_749/A gnd OAI21X1_1735/C vdd OAI21X1
XOAI21X1_1778 BUFX4_385/Y INVX2_150/Y NAND2X1_719/Y gnd OAI21X1_1778/Y vdd OAI21X1
XOAI21X1_1789 BUFX4_368/Y INVX2_161/Y NAND2X1_730/Y gnd OAI21X1_1789/Y vdd OAI21X1
XOAI21X1_1767 INVX2_145/Y BUFX4_290/Y OAI21X1_1767/C gnd DFFPOSX1_96/D vdd OAI21X1
XFILL_0_OAI21X1_712 gnd vdd FILL
XFILL_0_OAI21X1_723 gnd vdd FILL
XFILL_0_OAI21X1_701 gnd vdd FILL
XFILL_0_OAI21X1_745 gnd vdd FILL
XFILL_0_OAI21X1_756 gnd vdd FILL
XFILL_0_OAI21X1_734 gnd vdd FILL
XFILL_1_OAI21X1_905 gnd vdd FILL
XFILL_1_OAI21X1_927 gnd vdd FILL
XFILL_1_OAI21X1_916 gnd vdd FILL
XFILL_1_OAI21X1_949 gnd vdd FILL
XFILL_1_OAI21X1_938 gnd vdd FILL
XFILL_0_OAI21X1_767 gnd vdd FILL
XFILL_0_OAI21X1_778 gnd vdd FILL
XFILL_0_OAI21X1_789 gnd vdd FILL
XFILL_2_NAND3X1_28 gnd vdd FILL
XFILL_13_17_1 gnd vdd FILL
XFILL_0_OAI21X1_1500 gnd vdd FILL
XFILL_0_NAND2X1_740 gnd vdd FILL
XFILL_0_NAND2X1_762 gnd vdd FILL
XFILL_0_OAI21X1_1533 gnd vdd FILL
XFILL_0_NAND2X1_751 gnd vdd FILL
XFILL_0_OAI21X1_1522 gnd vdd FILL
XFILL_0_OAI21X1_1511 gnd vdd FILL
XFILL_24_9_1 gnd vdd FILL
XFILL_23_4_0 gnd vdd FILL
XFILL_0_OAI21X1_1566 gnd vdd FILL
XFILL_0_OAI21X1_1544 gnd vdd FILL
XFILL_0_OAI21X1_1555 gnd vdd FILL
XFILL_0_OAI21X1_1588 gnd vdd FILL
XFILL_0_OAI21X1_1599 gnd vdd FILL
XFILL_0_OAI21X1_1577 gnd vdd FILL
XFILL_5_DFFPOSX1_771 gnd vdd FILL
XFILL_5_DFFPOSX1_760 gnd vdd FILL
XFILL_5_DFFPOSX1_782 gnd vdd FILL
XFILL_5_DFFPOSX1_793 gnd vdd FILL
XFILL_18_16_1 gnd vdd FILL
XBUFX4_118 INVX8_4/Y gnd BUFX4_380/A vdd BUFX4
XBUFX4_107 BUFX4_2/A gnd BUFX4_107/Y vdd BUFX4
XFILL_6_5_0 gnd vdd FILL
XFILL_31_18_1 gnd vdd FILL
XBUFX4_129 BUFX4_15/Y gnd BUFX4_129/Y vdd BUFX4
XFILL_0_INVX1_18 gnd vdd FILL
XFILL_0_INVX1_29 gnd vdd FILL
XFILL_4_DFFPOSX1_350 gnd vdd FILL
XFILL_2_OAI21X1_1638 gnd vdd FILL
XFILL_4_DFFPOSX1_361 gnd vdd FILL
XFILL_4_DFFPOSX1_372 gnd vdd FILL
XFILL_2_DFFPOSX1_1020 gnd vdd FILL
XFILL_2_DFFPOSX1_1031 gnd vdd FILL
XFILL_4_DFFPOSX1_394 gnd vdd FILL
XFILL_12_12_0 gnd vdd FILL
XFILL_4_DFFPOSX1_383 gnd vdd FILL
XFILL_0_OAI22X1_2 gnd vdd FILL
XFILL_15_9_1 gnd vdd FILL
XFILL_14_4_0 gnd vdd FILL
XFILL_1_BUFX2_262 gnd vdd FILL
XFILL_1_BUFX2_240 gnd vdd FILL
XOAI21X1_1019 BUFX4_296/Y INVX1_164/Y OAI21X1_1019/C gnd OAI21X1_1019/Y vdd OAI21X1
XFILL_1_BUFX2_273 gnd vdd FILL
XFILL_1_BUFX2_284 gnd vdd FILL
XOAI21X1_1008 BUFX4_173/Y BUFX4_46/Y BUFX2_367/A gnd OAI21X1_1009/C vdd OAI21X1
XOAI21X1_290 BUFX4_164/Y BUFX4_79/Y BUFX2_1009/A gnd OAI21X1_291/C vdd OAI21X1
XFILL_1_OAI21X1_1228 gnd vdd FILL
XFILL_1_OAI21X1_1217 gnd vdd FILL
XFILL_1_OAI21X1_1239 gnd vdd FILL
XDFFPOSX1_609 BUFX2_643/A CLKBUF1_29/Y OAI21X1_837/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1206 gnd vdd FILL
XFILL_1_DFFPOSX1_818 gnd vdd FILL
XFILL_1_DFFPOSX1_807 gnd vdd FILL
XFILL_1_DFFPOSX1_829 gnd vdd FILL
XFILL_36_17_1 gnd vdd FILL
XFILL_6_DFFPOSX1_477 gnd vdd FILL
XFILL_17_11_0 gnd vdd FILL
XFILL_6_DFFPOSX1_466 gnd vdd FILL
XFILL_6_DFFPOSX1_455 gnd vdd FILL
XFILL_6_DFFPOSX1_499 gnd vdd FILL
XFILL_6_DFFPOSX1_488 gnd vdd FILL
XFILL_30_13_0 gnd vdd FILL
XFILL_1_NAND2X1_218 gnd vdd FILL
XFILL_1_NAND3X1_3 gnd vdd FILL
XFILL_1_NAND2X1_229 gnd vdd FILL
XFILL_1_NAND2X1_207 gnd vdd FILL
XFILL_36_1 gnd vdd FILL
XFILL_0_DFFPOSX1_408 gnd vdd FILL
XFILL_0_DFFPOSX1_419 gnd vdd FILL
XFILL_5_DFFPOSX1_1013 gnd vdd FILL
XFILL_5_DFFPOSX1_1024 gnd vdd FILL
XFILL_5_DFFPOSX1_1002 gnd vdd FILL
XDFFPOSX1_13 BUFX2_712/A CLKBUF1_57/Y DFFPOSX1_13/D gnd vdd DFFPOSX1
XDFFPOSX1_24 BUFX2_694/A CLKBUF1_67/Y DFFPOSX1_24/D gnd vdd DFFPOSX1
XOAI21X1_1520 BUFX4_128/Y BUFX4_47/Y BUFX2_233/A gnd OAI21X1_1521/C vdd OAI21X1
XOAI21X1_1531 INVX1_225/A INVX1_195/A INVX2_83/Y gnd NAND2X1_642/B vdd OAI21X1
XFILL_0_BUFX4_370 gnd vdd FILL
XDFFPOSX1_35 BUFX2_706/A CLKBUF1_41/Y DFFPOSX1_35/D gnd vdd DFFPOSX1
XDFFPOSX1_68 BUFX2_745/A CLKBUF1_25/Y DFFPOSX1_68/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1740 gnd vdd FILL
XDFFPOSX1_57 BUFX2_727/A CLKBUF1_61/Y DFFPOSX1_57/D gnd vdd DFFPOSX1
XDFFPOSX1_46 BUFX2_715/A CLKBUF1_8/Y DFFPOSX1_46/D gnd vdd DFFPOSX1
XOAI21X1_1575 BUFX4_328/Y INVX2_113/Y NAND2X1_648/Y gnd OAI21X1_1575/Y vdd OAI21X1
XFILL_0_BUFX4_381 gnd vdd FILL
XOAI21X1_1564 BUFX4_141/Y BUFX4_51/Y BUFX2_250/A gnd OAI21X1_1566/C vdd OAI21X1
XFILL_1_OAI21X1_1751 gnd vdd FILL
XOAI21X1_1542 AOI21X1_63/Y OAI21X1_1542/B OAI21X1_1542/C gnd OAI21X1_1542/Y vdd OAI21X1
XOAI21X1_1553 BUFX4_121/Y BUFX4_66/Y BUFX2_245/A gnd OAI21X1_1555/C vdd OAI21X1
XOAI21X1_1597 BUFX4_312/Y INVX2_133/Y NAND2X1_666/Y gnd OAI21X1_1597/Y vdd OAI21X1
XFILL_1_OAI21X1_1762 gnd vdd FILL
XDFFPOSX1_79 BUFX2_748/A CLKBUF1_22/Y DFFPOSX1_79/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_702 gnd vdd FILL
XFILL_0_OAI21X1_520 gnd vdd FILL
XFILL_1_OAI21X1_1784 gnd vdd FILL
XFILL_1_OAI21X1_1773 gnd vdd FILL
XOAI21X1_1586 OAI21X1_7/A INVX2_122/Y NAND2X1_655/Y gnd OAI21X1_1586/Y vdd OAI21X1
XFILL_0_OAI21X1_531 gnd vdd FILL
XFILL_1_OAI21X1_1795 gnd vdd FILL
XFILL_0_BUFX2_1030 gnd vdd FILL
XFILL_0_OAI21X1_553 gnd vdd FILL
XFILL_1_OAI21X1_713 gnd vdd FILL
XFILL_1_OAI21X1_735 gnd vdd FILL
XFILL_1_OAI21X1_724 gnd vdd FILL
XFILL_0_OAI21X1_542 gnd vdd FILL
XFILL_0_OAI21X1_564 gnd vdd FILL
XFILL_2_OAI21X1_928 gnd vdd FILL
XFILL_1_OAI21X1_768 gnd vdd FILL
XFILL_1_OAI21X1_757 gnd vdd FILL
XFILL_1_OAI21X1_779 gnd vdd FILL
XFILL_1_OAI21X1_746 gnd vdd FILL
XFILL_0_OAI21X1_597 gnd vdd FILL
XFILL_0_OAI21X1_575 gnd vdd FILL
XFILL_0_OAI21X1_586 gnd vdd FILL
XFILL_35_12_0 gnd vdd FILL
XFILL_0_CLKBUF1_20 gnd vdd FILL
XFILL_0_CLKBUF1_42 gnd vdd FILL
XFILL_0_CLKBUF1_31 gnd vdd FILL
XFILL_0_CLKBUF1_53 gnd vdd FILL
XFILL_0_CLKBUF1_86 gnd vdd FILL
XFILL_0_CLKBUF1_64 gnd vdd FILL
XFILL_0_CLKBUF1_97 gnd vdd FILL
XFILL_0_CLKBUF1_75 gnd vdd FILL
XFILL_1_NAND2X1_741 gnd vdd FILL
XFILL_1_NAND2X1_730 gnd vdd FILL
XFILL_0_OAI21X1_1341 gnd vdd FILL
XFILL_0_OAI21X1_1330 gnd vdd FILL
XFILL_0_NAND2X1_570 gnd vdd FILL
XFILL_0_OAI21X1_1385 gnd vdd FILL
XFILL_1_NAND2X1_763 gnd vdd FILL
XFILL_0_NAND2X1_592 gnd vdd FILL
XFILL_0_DFFPOSX1_942 gnd vdd FILL
XFILL_0_DFFPOSX1_920 gnd vdd FILL
XFILL_0_OAI21X1_1374 gnd vdd FILL
XFILL_0_DFFPOSX1_931 gnd vdd FILL
XFILL_0_NAND2X1_581 gnd vdd FILL
XFILL_0_OAI21X1_1352 gnd vdd FILL
XFILL_0_OAI21X1_1363 gnd vdd FILL
XFILL_0_OAI21X1_1396 gnd vdd FILL
XFILL_0_DFFPOSX1_953 gnd vdd FILL
XFILL_0_DFFPOSX1_964 gnd vdd FILL
XFILL_0_DFFPOSX1_986 gnd vdd FILL
XFILL_0_DFFPOSX1_975 gnd vdd FILL
XFILL_0_DFFPOSX1_997 gnd vdd FILL
XFILL_5_DFFPOSX1_590 gnd vdd FILL
XFILL_0_OR2X2_3 gnd vdd FILL
XINVX2_118 bundlePid_i[30] gnd INVX2_118/Y vdd INVX2
XFILL_0_BUFX2_318 gnd vdd FILL
XFILL_0_BUFX2_329 gnd vdd FILL
XINVX2_129 bundlePid_i[19] gnd INVX2_129/Y vdd INVX2
XINVX2_107 NOR3X1_17/B gnd INVX2_107/Y vdd INVX2
XFILL_0_BUFX2_307 gnd vdd FILL
XFILL_1_BUFX4_1 gnd vdd FILL
XFILL_4_DFFPOSX1_180 gnd vdd FILL
XFILL_2_OAI21X1_1424 gnd vdd FILL
XFILL_2_NOR3X1_13 gnd vdd FILL
XFILL_2_OAI21X1_1446 gnd vdd FILL
XFILL_4_DFFPOSX1_191 gnd vdd FILL
XFILL_0_INVX1_5 gnd vdd FILL
XFILL_30_7_1 gnd vdd FILL
XFILL_1_NAND3X1_36 gnd vdd FILL
XFILL_1_NAND3X1_25 gnd vdd FILL
XFILL_1_OAI21X1_1014 gnd vdd FILL
XFILL_1_OAI21X1_1003 gnd vdd FILL
XFILL_1_NAND3X1_14 gnd vdd FILL
XFILL_0_BUFX2_830 gnd vdd FILL
XFILL_0_BUFX2_841 gnd vdd FILL
XFILL_1_OAI21X1_1036 gnd vdd FILL
XFILL_1_OAI21X1_1047 gnd vdd FILL
XFILL_0_BUFX2_852 gnd vdd FILL
XDFFPOSX1_406 BUFX2_439/A CLKBUF1_91/Y OAI21X1_378/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_615 gnd vdd FILL
XFILL_1_DFFPOSX1_604 gnd vdd FILL
XFILL_1_NAND3X1_69 gnd vdd FILL
XFILL_1_NAND3X1_58 gnd vdd FILL
XFILL_1_INVX4_1 gnd vdd FILL
XFILL_1_NAND3X1_47 gnd vdd FILL
XDFFPOSX1_428 BUFX2_519/A CLKBUF1_13/Y OAI21X1_411/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1025 gnd vdd FILL
XDFFPOSX1_417 BUFX2_451/A CLKBUF1_24/Y OAI21X1_389/Y gnd vdd DFFPOSX1
XINVX1_140 bundle_i[64] gnd INVX1_140/Y vdd INVX1
XINVX1_151 bundle_i[117] gnd INVX1_151/Y vdd INVX1
XFILL_0_BUFX2_885 gnd vdd FILL
XFILL_1_OAI21X1_1069 gnd vdd FILL
XDFFPOSX1_439 BUFX2_468/A CLKBUF1_1/Y OAI21X1_429/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_874 gnd vdd FILL
XFILL_1_DFFPOSX1_648 gnd vdd FILL
XFILL_1_DFFPOSX1_626 gnd vdd FILL
XFILL_1_DFFPOSX1_637 gnd vdd FILL
XFILL_0_BUFX2_863 gnd vdd FILL
XFILL_1_OAI21X1_1058 gnd vdd FILL
XINVX1_184 INVX1_184/A gnd INVX1_184/Y vdd INVX1
XINVX1_195 INVX1_195/A gnd INVX1_195/Y vdd INVX1
XNAND2X1_509 bundleAddress_i[42] bundleAddress_i[41] gnd OR2X2_17/B vdd NAND2X1
XINVX1_173 bundleAddress_i[43] gnd INVX1_173/Y vdd INVX1
XFILL_0_BUFX2_896 gnd vdd FILL
XFILL_1_DFFPOSX1_659 gnd vdd FILL
XINVX1_162 bundle_i[106] gnd INVX1_162/Y vdd INVX1
XFILL_6_DFFPOSX1_252 gnd vdd FILL
XFILL_6_DFFPOSX1_230 gnd vdd FILL
XFILL_6_DFFPOSX1_241 gnd vdd FILL
XFILL_6_DFFPOSX1_263 gnd vdd FILL
XFILL_38_8_1 gnd vdd FILL
XFILL_37_3_0 gnd vdd FILL
XFILL_0_INVX2_61 gnd vdd FILL
XFILL_0_INVX2_72 gnd vdd FILL
XFILL_0_INVX2_50 gnd vdd FILL
XFILL_0_INVX2_94 gnd vdd FILL
XFILL_0_INVX2_83 gnd vdd FILL
XFILL_1_NOR3X1_3 gnd vdd FILL
XFILL_0_DFFPOSX1_205 gnd vdd FILL
XFILL_0_DFFPOSX1_238 gnd vdd FILL
XFILL_0_DFFPOSX1_216 gnd vdd FILL
XFILL_0_DFFPOSX1_227 gnd vdd FILL
XFILL_0_DFFPOSX1_249 gnd vdd FILL
XFILL_21_7_1 gnd vdd FILL
XFILL_20_2_0 gnd vdd FILL
XFILL_3_DFFPOSX1_709 gnd vdd FILL
XFILL_3_CLKBUF1_19 gnd vdd FILL
XFILL_21_18_0 gnd vdd FILL
XOAI21X1_1350 BUFX4_1/Y BUFX4_357/Y BUFX2_177/A gnd OAI21X1_1352/C vdd OAI21X1
XDFFPOSX1_951 BUFX2_200/A CLKBUF1_1/Y OAI21X1_1429/Y gnd vdd DFFPOSX1
XDFFPOSX1_940 BUFX2_227/A CLKBUF1_84/Y OAI21X1_1395/Y gnd vdd DFFPOSX1
XOAI21X1_1383 XNOR2X1_89/Y BUFX4_162/Y OAI21X1_1383/C gnd OAI21X1_1383/Y vdd OAI21X1
XOAI21X1_1372 BUFX4_1/A BUFX4_330/Y BUFX2_184/A gnd OAI21X1_1373/C vdd OAI21X1
XOAI21X1_1361 BUFX4_1/A BUFX4_374/Y BUFX2_181/A gnd OAI21X1_1364/C vdd OAI21X1
XFILL_1_OAI21X1_1581 gnd vdd FILL
XFILL_1_OAI21X1_1592 gnd vdd FILL
XDFFPOSX1_962 BUFX2_212/A CLKBUF1_55/Y OAI21X1_1460/Y gnd vdd DFFPOSX1
XDFFPOSX1_984 BUFX2_236/A CLKBUF1_30/Y OAI21X1_1530/Y gnd vdd DFFPOSX1
XOAI21X1_1394 BUFX4_145/Y BUFX4_33/Y BUFX2_227/A gnd OAI21X1_1395/C vdd OAI21X1
XFILL_1_OAI21X1_1570 gnd vdd FILL
XDFFPOSX1_973 BUFX2_224/A CLKBUF1_85/Y OAI21X1_1496/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_510 gnd vdd FILL
XFILL_1_NOR2X1_104 gnd vdd FILL
XFILL_2_OAI21X1_714 gnd vdd FILL
XFILL_1_NOR2X1_115 gnd vdd FILL
XFILL_1_OAI21X1_554 gnd vdd FILL
XDFFPOSX1_995 BUFX2_248/A CLKBUF1_69/Y OAI21X1_1563/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_372 gnd vdd FILL
XFILL_1_OAI21X1_543 gnd vdd FILL
XFILL_0_OAI21X1_350 gnd vdd FILL
XFILL_1_OAI21X1_532 gnd vdd FILL
XFILL_1_OAI21X1_521 gnd vdd FILL
XFILL_0_OAI21X1_361 gnd vdd FILL
XFILL_2_OAI21X1_758 gnd vdd FILL
XFILL_1_OAI21X1_576 gnd vdd FILL
XFILL_0_OAI21X1_394 gnd vdd FILL
XFILL_1_NOR2X1_159 gnd vdd FILL
XFILL_0_OAI21X1_383 gnd vdd FILL
XFILL_1_OAI21X1_565 gnd vdd FILL
XFILL_1_OAI21X1_587 gnd vdd FILL
XFILL_1_OAI21X1_598 gnd vdd FILL
XFILL_29_8_1 gnd vdd FILL
XFILL_28_3_0 gnd vdd FILL
XBUFX2_408 BUFX2_408/A gnd majID1_o[41] vdd BUFX2
XFILL_4_8_1 gnd vdd FILL
XFILL_3_3_0 gnd vdd FILL
XBUFX2_419 BUFX2_419/A gnd majID1_o[31] vdd BUFX2
XFILL_1_BUFX4_313 gnd vdd FILL
XFILL_1_NAND2X1_560 gnd vdd FILL
XFILL_1_BUFX4_302 gnd vdd FILL
XFILL_0_OAI21X1_1160 gnd vdd FILL
XFILL_0_DFFPOSX1_761 gnd vdd FILL
XFILL_1_NAND2X1_593 gnd vdd FILL
XFILL_0_DFFPOSX1_750 gnd vdd FILL
XFILL_0_OAI21X1_1171 gnd vdd FILL
XFILL_1_NAND2X1_582 gnd vdd FILL
XFILL_1_BUFX4_346 gnd vdd FILL
XFILL_1_BUFX4_324 gnd vdd FILL
XFILL_0_OAI21X1_1182 gnd vdd FILL
XFILL_0_OAI21X1_1193 gnd vdd FILL
XFILL_1_BUFX4_335 gnd vdd FILL
XFILL_1_BUFX4_368 gnd vdd FILL
XFILL_1_BUFX4_379 gnd vdd FILL
XFILL_26_17_0 gnd vdd FILL
XFILL_0_DFFPOSX1_772 gnd vdd FILL
XFILL_1_BUFX4_357 gnd vdd FILL
XFILL_12_7_1 gnd vdd FILL
XFILL_11_2_0 gnd vdd FILL
XFILL_0_DFFPOSX1_783 gnd vdd FILL
XFILL_0_DFFPOSX1_794 gnd vdd FILL
XFILL_2_OAI21X1_15 gnd vdd FILL
XFILL_0_BUFX2_104 gnd vdd FILL
XFILL_0_BUFX2_126 gnd vdd FILL
XFILL_0_BUFX2_137 gnd vdd FILL
XFILL_0_BUFX2_115 gnd vdd FILL
XFILL_0_BUFX2_148 gnd vdd FILL
XFILL_0_BUFX2_159 gnd vdd FILL
XFILL_1_NAND2X1_91 gnd vdd FILL
XFILL_1_NAND2X1_80 gnd vdd FILL
XFILL_2_OAI21X1_1210 gnd vdd FILL
XFILL_19_3_0 gnd vdd FILL
XFILL_2_DFFPOSX1_822 gnd vdd FILL
XFILL_2_OAI21X1_1254 gnd vdd FILL
XFILL_2_DFFPOSX1_811 gnd vdd FILL
XFILL_2_DFFPOSX1_833 gnd vdd FILL
XBUFX2_920 BUFX2_920/A gnd tid3_o[41] vdd BUFX2
XFILL_2_DFFPOSX1_800 gnd vdd FILL
XBUFX2_931 BUFX2_931/A gnd tid3_o[31] vdd BUFX2
XFILL_2_DFFPOSX1_855 gnd vdd FILL
XFILL_2_DFFPOSX1_866 gnd vdd FILL
XBUFX2_964 BUFX2_964/A gnd tid3_o[1] vdd BUFX2
XFILL_1_18_0 gnd vdd FILL
XFILL_2_DFFPOSX1_844 gnd vdd FILL
XBUFX2_942 BUFX2_942/A gnd tid3_o[21] vdd BUFX2
XBUFX2_953 BUFX2_953/A gnd tid3_o[11] vdd BUFX2
XBUFX2_975 BUFX2_975/A gnd tid4_o[49] vdd BUFX2
XBUFX2_986 BUFX2_986/A gnd tid4_o[39] vdd BUFX2
XBUFX2_997 BUFX2_997/A gnd tid4_o[29] vdd BUFX2
XFILL_2_DFFPOSX1_888 gnd vdd FILL
XFILL_2_DFFPOSX1_877 gnd vdd FILL
XFILL_2_DFFPOSX1_899 gnd vdd FILL
XDFFPOSX1_203 BUFX2_874/A CLKBUF1_40/Y OAI21X1_47/Y gnd vdd DFFPOSX1
XDFFPOSX1_214 BUFX2_887/A CLKBUF1_57/Y OAI21X1_58/Y gnd vdd DFFPOSX1
XDFFPOSX1_225 BUFX2_899/A CLKBUF1_78/Y OAI21X1_69/Y gnd vdd DFFPOSX1
XBUFX4_9 BUFX4_9/A gnd BUFX4_9/Y vdd BUFX4
XFILL_1_DFFPOSX1_412 gnd vdd FILL
XFILL_0_BUFX2_660 gnd vdd FILL
XFILL_1_DFFPOSX1_423 gnd vdd FILL
XFILL_1_DFFPOSX1_401 gnd vdd FILL
XDFFPOSX1_236 BUFX2_967/A CLKBUF1_56/Y OAI21X1_89/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_682 gnd vdd FILL
XDFFPOSX1_258 BUFX2_929/A CLKBUF1_102/Y OAI21X1_133/Y gnd vdd DFFPOSX1
XDFFPOSX1_247 BUFX2_916/A CLKBUF1_23/Y OAI21X1_111/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_456 gnd vdd FILL
XFILL_1_DFFPOSX1_445 gnd vdd FILL
XFILL_0_BUFX2_693 gnd vdd FILL
XFILL_0_BUFX2_671 gnd vdd FILL
XFILL_1_DFFPOSX1_434 gnd vdd FILL
XDFFPOSX1_269 BUFX2_941/A CLKBUF1_37/Y OAI21X1_155/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_478 gnd vdd FILL
XNAND2X1_306 NOR2X1_99/Y NOR2X1_97/Y gnd OAI21X1_656/A vdd NAND2X1
XNAND2X1_317 bundleStartMajId_i[43] NOR2X1_106/Y gnd INVX1_37/A vdd NAND2X1
XFILL_1_DFFPOSX1_489 gnd vdd FILL
XFILL_1_DFFPOSX1_467 gnd vdd FILL
XFILL_4_DFFPOSX1_905 gnd vdd FILL
XNAND2X1_328 OAI21X1_770/Y INVX4_31/Y gnd OAI21X1_772/A vdd NAND2X1
XNAND2X1_339 BUFX4_268/Y bundle_i[30] gnd OAI21X1_845/C vdd NAND2X1
XFILL_4_DFFPOSX1_938 gnd vdd FILL
XFILL_4_DFFPOSX1_916 gnd vdd FILL
XFILL_4_DFFPOSX1_927 gnd vdd FILL
XFILL_6_17_0 gnd vdd FILL
XFILL_4_DFFPOSX1_949 gnd vdd FILL
XNOR3X1_13 INVX2_85/Y INVX2_86/Y NOR3X1_13/C gnd NOR3X1_13/Y vdd NOR3X1
XBUFX4_290 BUFX4_303/A gnd BUFX4_290/Y vdd BUFX4
XFILL_10_15_1 gnd vdd FILL
XFILL_0_XNOR2X1_5 gnd vdd FILL
XFILL_1_BUFX2_817 gnd vdd FILL
XFILL_1_BUFX2_806 gnd vdd FILL
XOAI21X1_812 BUFX4_161/Y BUFX4_43/Y BUFX2_633/A gnd OAI21X1_813/C vdd OAI21X1
XOAI21X1_823 BUFX4_127/Y BUFX4_27/Y BUFX2_637/A gnd OAI21X1_824/C vdd OAI21X1
XOAI21X1_801 XNOR2X1_53/Y BUFX4_299/Y OAI21X1_801/C gnd OAI21X1_801/Y vdd OAI21X1
XINVX4_9 bundleStartMajId_i[40] gnd INVX4_9/Y vdd INVX4
XOAI21X1_867 INVX1_68/Y BUFX4_263/Y OAI21X1_867/C gnd OAI21X1_867/Y vdd OAI21X1
XFILL_3_DFFPOSX1_528 gnd vdd FILL
XOAI21X1_845 INVX1_46/Y BUFX4_265/Y OAI21X1_845/C gnd OAI21X1_845/Y vdd OAI21X1
XOAI21X1_834 OAI21X1_834/A BUFX4_299/Y OAI21X1_834/C gnd OAI21X1_834/Y vdd OAI21X1
XOAI21X1_856 INVX1_57/Y BUFX4_264/Y OAI21X1_856/C gnd OAI21X1_856/Y vdd OAI21X1
XFILL_3_DFFPOSX1_506 gnd vdd FILL
XFILL_3_DFFPOSX1_517 gnd vdd FILL
XOAI21X1_889 INVX1_90/Y BUFX4_205/Y OAI21X1_889/C gnd OAI21X1_889/Y vdd OAI21X1
XOAI21X1_878 INVX1_79/Y BUFX4_211/Y OAI21X1_878/C gnd OAI21X1_878/Y vdd OAI21X1
XFILL_3_DFFPOSX1_539 gnd vdd FILL
XOAI21X1_1180 NOR3X1_14/C INVX4_44/Y BUFX4_239/Y gnd OAI21X1_1181/B vdd OAI21X1
XOAI21X1_1191 OAI21X1_1191/A NOR2X1_170/Y NAND2X1_577/Y gnd OAI21X1_1191/Y vdd OAI21X1
XDFFPOSX1_792 BUFX2_44/A CLKBUF1_67/Y OAI21X1_1084/Y gnd vdd DFFPOSX1
XDFFPOSX1_770 BUFX2_20/A CLKBUF1_35/Y OAI21X1_1062/Y gnd vdd DFFPOSX1
XDFFPOSX1_781 BUFX2_32/A CLKBUF1_77/Y OAI21X1_1073/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_180 gnd vdd FILL
XFILL_1_OAI21X1_340 gnd vdd FILL
XFILL_1_OAI21X1_351 gnd vdd FILL
XFILL_1_OAI21X1_362 gnd vdd FILL
XFILL_0_OAI21X1_191 gnd vdd FILL
XFILL_1_DFFPOSX1_990 gnd vdd FILL
XFILL_1_CLKBUF1_5 gnd vdd FILL
XFILL_1_OAI21X1_384 gnd vdd FILL
XFILL_1_OAI21X1_395 gnd vdd FILL
XFILL_1_OAI21X1_373 gnd vdd FILL
XFILL_0_NAND3X1_11 gnd vdd FILL
XFILL_15_14_1 gnd vdd FILL
XBUFX2_216 BUFX2_216/A gnd addr4_o[60] vdd BUFX2
XFILL_2_DFFPOSX1_118 gnd vdd FILL
XBUFX2_205 BUFX2_205/A gnd addr4_o[61] vdd BUFX2
XFILL_2_DFFPOSX1_107 gnd vdd FILL
XFILL_0_NAND3X1_33 gnd vdd FILL
XFILL_0_NAND3X1_22 gnd vdd FILL
XFILL_0_NAND3X1_44 gnd vdd FILL
XBUFX2_238 BUFX2_238/A gnd addr4_o[58] vdd BUFX2
XBUFX2_249 BUFX2_249/A gnd addr4_o[57] vdd BUFX2
XFILL_0_NAND3X1_55 gnd vdd FILL
XBUFX2_227 BUFX2_227/A gnd addr4_o[59] vdd BUFX2
XFILL_0_NAND3X1_66 gnd vdd FILL
XFILL_2_DFFPOSX1_129 gnd vdd FILL
XFILL_0_BUFX4_90 gnd vdd FILL
XFILL_1_BUFX4_110 gnd vdd FILL
XFILL_1_BUFX4_121 gnd vdd FILL
XFILL_1_NAND2X1_390 gnd vdd FILL
XFILL_1_BUFX4_143 gnd vdd FILL
XFILL_1_BUFX4_132 gnd vdd FILL
XFILL_1_BUFX4_154 gnd vdd FILL
XFILL_1_BUFX4_165 gnd vdd FILL
XFILL_1_BUFX4_198 gnd vdd FILL
XFILL_0_DFFPOSX1_591 gnd vdd FILL
XFILL_0_DFFPOSX1_580 gnd vdd FILL
XFILL_1_BUFX4_187 gnd vdd FILL
XFILL_1_BUFX4_176 gnd vdd FILL
XFILL_1_MUX2X1_1 gnd vdd FILL
XFILL_33_15_1 gnd vdd FILL
XFILL_2_CLKBUF1_16 gnd vdd FILL
XFILL_2_CLKBUF1_27 gnd vdd FILL
XFILL_2_CLKBUF1_38 gnd vdd FILL
XFILL_2_DFFPOSX1_630 gnd vdd FILL
XFILL_2_CLKBUF1_49 gnd vdd FILL
XFILL_2_DFFPOSX1_641 gnd vdd FILL
XBUFX2_761 BUFX2_761/A gnd pid4_o[8] vdd BUFX2
XFILL_35_6_1 gnd vdd FILL
XFILL_34_1_0 gnd vdd FILL
XBUFX2_750 BUFX2_750/A gnd pid4_o[18] vdd BUFX2
XNOR2X1_90 INVX2_32/Y INVX4_22/Y gnd NOR2X1_90/Y vdd NOR2X1
XFILL_2_DFFPOSX1_652 gnd vdd FILL
XFILL_2_DFFPOSX1_663 gnd vdd FILL
XFILL_2_DFFPOSX1_674 gnd vdd FILL
XBUFX2_772 BUFX2_772/A gnd pid4_o[26] vdd BUFX2
XBUFX2_783 BUFX2_783/A gnd tid1_o[49] vdd BUFX2
XBUFX2_794 BUFX2_794/A gnd tid1_o[39] vdd BUFX2
XFILL_0_NOR2X1_101 gnd vdd FILL
XFILL_0_NOR2X1_112 gnd vdd FILL
XFILL_2_DFFPOSX1_696 gnd vdd FILL
XFILL_2_DFFPOSX1_685 gnd vdd FILL
XFILL_0_NOR2X1_123 gnd vdd FILL
XFILL_0_NOR2X1_134 gnd vdd FILL
XFILL_0_NOR2X1_145 gnd vdd FILL
XOAI21X1_119 BUFX4_172/Y INVX2_169/Y OAI21X1_119/C gnd OAI21X1_119/Y vdd OAI21X1
XFILL_0_NOR2X1_178 gnd vdd FILL
XOAI21X1_108 BUFX4_97/Y BUFX4_377/Y BUFX2_915/A gnd OAI21X1_109/C vdd OAI21X1
XFILL_0_NOR2X1_167 gnd vdd FILL
XFILL_0_NOR2X1_189 gnd vdd FILL
XFILL_0_NOR2X1_156 gnd vdd FILL
XFILL_0_DFFPOSX1_1019 gnd vdd FILL
XFILL_0_DFFPOSX1_1008 gnd vdd FILL
XBUFX2_6 BUFX2_6/A gnd addr1_o[50] vdd BUFX2
XFILL_1_DFFPOSX1_220 gnd vdd FILL
XFILL_1_DFFPOSX1_231 gnd vdd FILL
XFILL_0_BUFX2_490 gnd vdd FILL
XFILL_1_DFFPOSX1_242 gnd vdd FILL
XFILL_1_DFFPOSX1_253 gnd vdd FILL
XFILL_1_DFFPOSX1_264 gnd vdd FILL
XFILL_38_14_1 gnd vdd FILL
XFILL_1_DFFPOSX1_275 gnd vdd FILL
XNAND2X1_125 BUFX2_442/A BUFX4_325/Y gnd OAI21X1_381/C vdd NAND2X1
XNAND2X1_114 BUFX2_430/A BUFX4_372/Y gnd OAI21X1_370/C vdd NAND2X1
XFILL_1_DFFPOSX1_297 gnd vdd FILL
XFILL_1_DFFPOSX1_286 gnd vdd FILL
XNAND2X1_103 BUFX2_418/A BUFX4_314/Y gnd OAI21X1_359/C vdd NAND2X1
XFILL_4_DFFPOSX1_713 gnd vdd FILL
XFILL_4_DFFPOSX1_702 gnd vdd FILL
XNAND2X1_158 BUFX2_460/A BUFX4_225/Y gnd OAI21X1_416/C vdd NAND2X1
XNAND2X1_136 BUFX2_457/A BUFX4_237/Y gnd OAI21X1_392/C vdd NAND2X1
XNAND2X1_147 bundleStartMajId_i[58] bundleStartMajId_i[57] gnd NOR2X1_60/A vdd NAND2X1
XNAND2X1_169 BUFX2_465/A BUFX4_236/Y gnd OAI21X1_424/C vdd NAND2X1
XFILL_1_OAI21X1_34 gnd vdd FILL
XFILL_1_OAI21X1_23 gnd vdd FILL
XFILL_1_OAI21X1_12 gnd vdd FILL
XNAND2X1_1 NAND2X1_1/A OAI21X1_1/A gnd OAI21X1_1/C vdd NAND2X1
XFILL_4_DFFPOSX1_746 gnd vdd FILL
XFILL_4_DFFPOSX1_735 gnd vdd FILL
XFILL_4_DFFPOSX1_724 gnd vdd FILL
XFILL_1_OAI21X1_56 gnd vdd FILL
XFILL_32_10_0 gnd vdd FILL
XFILL_4_DFFPOSX1_757 gnd vdd FILL
XFILL_1_OAI21X1_45 gnd vdd FILL
XFILL_1_OAI21X1_67 gnd vdd FILL
XFILL_4_DFFPOSX1_779 gnd vdd FILL
XFILL_4_DFFPOSX1_768 gnd vdd FILL
XFILL_1_OAI21X1_78 gnd vdd FILL
XFILL_1_OAI21X1_89 gnd vdd FILL
XFILL_26_6_1 gnd vdd FILL
XFILL_25_1_0 gnd vdd FILL
XFILL_1_6_1 gnd vdd FILL
XFILL_0_1_0 gnd vdd FILL
XNOR2X1_180 NOR2X1_180/A NOR2X1_180/B gnd NOR2X1_180/Y vdd NOR2X1
XNOR2X1_191 OR2X2_17/Y OR2X2_19/Y gnd INVX1_205/A vdd NOR2X1
XFILL_1_BUFX2_603 gnd vdd FILL
XFILL_1_BUFX2_614 gnd vdd FILL
XINVX2_6 bundleTid_i[1] gnd INVX2_6/Y vdd INVX2
XFILL_1_BUFX2_658 gnd vdd FILL
XFILL_1_BUFX2_669 gnd vdd FILL
XFILL_3_DFFPOSX1_303 gnd vdd FILL
XOAI21X1_642 NOR2X1_97/B OR2X2_13/Y INVX4_25/Y gnd OAI21X1_642/Y vdd OAI21X1
XOAI21X1_631 BUFX4_9/Y BUFX4_325/Y BUFX2_569/A gnd OAI21X1_633/C vdd OAI21X1
XOAI21X1_620 OAI21X1_620/A AOI21X1_15/Y OAI21X1_620/C gnd OAI21X1_620/Y vdd OAI21X1
XFILL_1_BUFX2_647 gnd vdd FILL
XFILL_3_DFFPOSX1_336 gnd vdd FILL
XFILL_3_DFFPOSX1_325 gnd vdd FILL
XOAI21X1_653 OAI21X1_656/A INVX4_27/Y BUFX4_305/Y gnd OAI21X1_654/B vdd OAI21X1
XAOI21X1_6 bundleStartMajId_i[2] NOR3X1_4/Y bundleStartMajId_i[1] gnd AOI21X1_6/Y
+ vdd AOI21X1
XFILL_3_DFFPOSX1_314 gnd vdd FILL
XOAI21X1_664 BUFX4_176/Y BUFX4_57/Y BUFX2_597/A gnd OAI21X1_665/C vdd OAI21X1
XOAI21X1_675 OAI21X1_675/A BUFX4_302/Y OAI21X1_675/C gnd OAI21X1_675/Y vdd OAI21X1
XFILL_3_DFFPOSX1_358 gnd vdd FILL
XFILL_3_DFFPOSX1_347 gnd vdd FILL
XOAI21X1_697 XNOR2X1_42/Y BUFX4_299/Y OAI21X1_697/C gnd OAI21X1_697/Y vdd OAI21X1
XOAI21X1_686 INVX1_35/A OR2X2_1/A BUFX4_285/Y gnd OAI21X1_688/B vdd OAI21X1
XFILL_3_DFFPOSX1_369 gnd vdd FILL
XFILL_0_INVX4_18 gnd vdd FILL
XFILL_0_INVX4_29 gnd vdd FILL
XXNOR2X1_14 NOR2X1_24/Y bundleStartMajId_i[28] gnd XNOR2X1_14/Y vdd XNOR2X1
XFILL_8_2_0 gnd vdd FILL
XFILL_9_7_1 gnd vdd FILL
XXNOR2X1_36 NOR2X1_87/B INVX4_20/Y gnd XNOR2X1_36/Y vdd XNOR2X1
XFILL_1_OAI21X1_170 gnd vdd FILL
XXNOR2X1_25 INVX4_30/A bundleStartMajId_i[54] gnd XNOR2X1_25/Y vdd XNOR2X1
XXNOR2X1_47 XNOR2X1_47/A INVX4_14/Y gnd XNOR2X1_47/Y vdd XNOR2X1
XFILL_2_OAI21X1_341 gnd vdd FILL
XFILL_1_INVX2_143 gnd vdd FILL
XFILL_1_OAI21X1_181 gnd vdd FILL
XNAND2X1_670 BUFX2_662/A BUFX4_339/Y gnd NAND2X1_670/Y vdd NAND2X1
XXNOR2X1_58 OR2X2_16/Y INVX4_34/Y gnd XNOR2X1_58/Y vdd XNOR2X1
XFILL_2_OAI21X1_385 gnd vdd FILL
XXNOR2X1_69 XNOR2X1_69/A INVX4_41/Y gnd XNOR2X1_69/Y vdd XNOR2X1
XINVX1_60 INVX1_60/A gnd INVX1_60/Y vdd INVX1
XNAND2X1_681 BUFX2_674/A BUFX4_320/Y gnd NAND2X1_681/Y vdd NAND2X1
XFILL_2_OAI21X1_352 gnd vdd FILL
XFILL_1_OAI21X1_192 gnd vdd FILL
XINVX1_93 bundle_i[47] gnd INVX1_93/Y vdd INVX1
XNAND2X1_692 BUFX2_683/A BUFX4_193/Y gnd NAND2X1_692/Y vdd NAND2X1
XINVX1_82 bundle_i[58] gnd INVX1_82/Y vdd INVX1
XINVX1_71 INVX1_71/A gnd INVX1_71/Y vdd INVX1
XFILL_2_OAI21X1_396 gnd vdd FILL
XBUFX2_24 BUFX2_24/A gnd addr1_o[60] vdd BUFX2
XBUFX2_13 BUFX2_13/A gnd addr1_o[61] vdd BUFX2
XBUFX2_35 BUFX2_35/A gnd addr1_o[59] vdd BUFX2
XBUFX2_68 BUFX2_68/A gnd addr2_o[52] vdd BUFX2
XBUFX2_57 BUFX2_57/A gnd addr1_o[57] vdd BUFX2
XBUFX2_46 BUFX2_46/A gnd addr1_o[58] vdd BUFX2
XFILL_17_6_1 gnd vdd FILL
XFILL_16_1_0 gnd vdd FILL
XDFFPOSX1_1 BUFX2_671/A CLKBUF1_38/Y DFFPOSX1_1/D gnd vdd DFFPOSX1
XBUFX2_79 BUFX2_79/A gnd addr2_o[42] vdd BUFX2
XFILL_5_DFFPOSX1_408 gnd vdd FILL
XFILL_5_DFFPOSX1_419 gnd vdd FILL
XFILL_1_BUFX4_35 gnd vdd FILL
XFILL_1_BUFX4_24 gnd vdd FILL
XFILL_1_BUFX4_13 gnd vdd FILL
XFILL_1_BUFX4_57 gnd vdd FILL
XFILL_1_BUFX4_46 gnd vdd FILL
XFILL_1_BUFX4_79 gnd vdd FILL
XFILL_1_BUFX4_68 gnd vdd FILL
XFILL_3_DFFPOSX1_881 gnd vdd FILL
XFILL_3_DFFPOSX1_870 gnd vdd FILL
XFILL_3_DFFPOSX1_892 gnd vdd FILL
XFILL_0_OAI21X1_905 gnd vdd FILL
XNOR2X1_4 NOR2X1_4/A NOR2X1_4/B gnd NOR2X1_4/Y vdd NOR2X1
XFILL_0_OAI21X1_938 gnd vdd FILL
XFILL_0_OAI21X1_927 gnd vdd FILL
XFILL_0_OAI21X1_916 gnd vdd FILL
XFILL_0_OAI21X1_949 gnd vdd FILL
XFILL_1_OR2X2_16 gnd vdd FILL
XFILL_0_OAI21X1_1715 gnd vdd FILL
XFILL_0_OAI21X1_1704 gnd vdd FILL
XFILL_0_OAI21X1_1726 gnd vdd FILL
XBUFX2_580 BUFX2_580/A gnd majID3_o[1] vdd BUFX2
XFILL_0_OAI21X1_1759 gnd vdd FILL
XFILL_0_OAI21X1_1737 gnd vdd FILL
XFILL_2_DFFPOSX1_471 gnd vdd FILL
XFILL_2_DFFPOSX1_482 gnd vdd FILL
XFILL_0_OAI21X1_1748 gnd vdd FILL
XFILL_2_DFFPOSX1_460 gnd vdd FILL
XFILL_2_DFFPOSX1_493 gnd vdd FILL
XBUFX2_591 BUFX2_591/A gnd majID4_o[49] vdd BUFX2
XFILL_5_DFFPOSX1_920 gnd vdd FILL
XFILL_5_DFFPOSX1_931 gnd vdd FILL
XFILL_5_DFFPOSX1_942 gnd vdd FILL
XFILL_5_DFFPOSX1_953 gnd vdd FILL
XFILL_5_DFFPOSX1_964 gnd vdd FILL
XAOI21X1_25 bundleStartMajId_i[4] NOR2X1_98/B bundleStartMajId_i[3] gnd AOI21X1_25/Y
+ vdd AOI21X1
XFILL_5_DFFPOSX1_997 gnd vdd FILL
XAOI21X1_14 bundleStartMajId_i[20] NOR2X1_85/B bundleStartMajId_i[19] gnd AOI21X1_14/Y
+ vdd AOI21X1
XFILL_5_DFFPOSX1_986 gnd vdd FILL
XFILL_5_DFFPOSX1_975 gnd vdd FILL
XAOI21X1_36 bundleAddress_i[61] INVX1_183/Y bundleAddress_i[58] gnd AOI21X1_36/Y vdd
+ AOI21X1
XAOI21X1_47 bundleAddress_i[36] NOR2X1_193/Y bundleAddress_i[35] gnd AOI21X1_47/Y
+ vdd AOI21X1
XAOI21X1_58 bundleAddress_i[4] XNOR2X1_88/A bundleAddress_i[3] gnd AOI21X1_58/Y vdd
+ AOI21X1
XOAI21X1_9 OAI21X1_9/A OAI21X1_9/B OAI21X1_9/C gnd OAI21X1_9/Y vdd OAI21X1
XFILL_4_DFFPOSX1_510 gnd vdd FILL
XFILL_4_DFFPOSX1_521 gnd vdd FILL
XFILL_4_DFFPOSX1_543 gnd vdd FILL
XFILL_4_DFFPOSX1_532 gnd vdd FILL
XFILL_4_DFFPOSX1_554 gnd vdd FILL
XFILL_4_DFFPOSX1_598 gnd vdd FILL
XFILL_4_DFFPOSX1_587 gnd vdd FILL
XFILL_4_DFFPOSX1_576 gnd vdd FILL
XFILL_4_DFFPOSX1_565 gnd vdd FILL
XFILL_1_BUFX2_1001 gnd vdd FILL
XFILL_1_BUFX2_1012 gnd vdd FILL
XFILL_1_BUFX2_411 gnd vdd FILL
XFILL_1_BUFX2_400 gnd vdd FILL
XFILL_1_BUFX2_422 gnd vdd FILL
XFILL_1_BUFX2_444 gnd vdd FILL
XFILL_3_DFFPOSX1_111 gnd vdd FILL
XFILL_3_DFFPOSX1_100 gnd vdd FILL
XFILL_23_15_0 gnd vdd FILL
XFILL_1_BUFX2_466 gnd vdd FILL
XFILL_1_BUFX2_455 gnd vdd FILL
XFILL_1_CLKBUF1_13 gnd vdd FILL
XOAI21X1_450 XNOR2X1_13/Y BUFX4_194/Y OAI21X1_450/C gnd OAI21X1_450/Y vdd OAI21X1
XFILL_3_DFFPOSX1_133 gnd vdd FILL
XFILL_3_DFFPOSX1_144 gnd vdd FILL
XFILL_3_DFFPOSX1_122 gnd vdd FILL
XFILL_1_CLKBUF1_35 gnd vdd FILL
XOAI21X1_472 INVX1_19/Y bundleStartMajId_i[15] BUFX4_241/Y gnd OAI21X1_473/A vdd OAI21X1
XFILL_3_DFFPOSX1_155 gnd vdd FILL
XOAI21X1_461 OAI21X1_461/A BUFX4_204/Y OAI21X1_461/C gnd OAI21X1_461/Y vdd OAI21X1
XFILL_1_CLKBUF1_24 gnd vdd FILL
XOAI21X1_483 OAI21X1_483/A NOR2X1_49/Y OAI21X1_483/C gnd OAI21X1_483/Y vdd OAI21X1
XFILL_1_BUFX2_499 gnd vdd FILL
XFILL_1_CLKBUF1_46 gnd vdd FILL
XFILL_3_DFFPOSX1_188 gnd vdd FILL
XFILL_1_CLKBUF1_57 gnd vdd FILL
XFILL_1_CLKBUF1_68 gnd vdd FILL
XOAI21X1_494 OAI21X1_494/A AOI21X1_5/Y OAI21X1_494/C gnd OAI21X1_494/Y vdd OAI21X1
XFILL_1_CLKBUF1_79 gnd vdd FILL
XFILL_3_DFFPOSX1_166 gnd vdd FILL
XFILL_3_DFFPOSX1_177 gnd vdd FILL
XFILL_3_DFFPOSX1_199 gnd vdd FILL
XFILL_6_DFFPOSX1_648 gnd vdd FILL
XFILL_6_DFFPOSX1_659 gnd vdd FILL
XFILL_6_DFFPOSX1_637 gnd vdd FILL
XFILL_0_NAND2X1_207 gnd vdd FILL
XFILL_0_INVX1_221 gnd vdd FILL
XFILL_0_INVX1_210 gnd vdd FILL
XFILL_0_NAND2X1_218 gnd vdd FILL
XFILL_0_NAND2X1_229 gnd vdd FILL
XFILL_32_4_1 gnd vdd FILL
XFILL_28_14_0 gnd vdd FILL
XFILL_5_DFFPOSX1_205 gnd vdd FILL
XFILL_5_DFFPOSX1_216 gnd vdd FILL
XFILL_5_DFFPOSX1_249 gnd vdd FILL
XFILL_5_DFFPOSX1_238 gnd vdd FILL
XFILL_5_DFFPOSX1_227 gnd vdd FILL
XFILL_0_OAI21X1_42 gnd vdd FILL
XFILL_0_OAI21X1_20 gnd vdd FILL
XFILL_0_OAI21X1_31 gnd vdd FILL
XFILL_0_OAI21X1_64 gnd vdd FILL
XFILL_0_OAI21X1_53 gnd vdd FILL
XOAI21X1_1713 INVX2_118/Y BUFX4_289/Y OAI21X1_1713/C gnd DFFPOSX1_69/D vdd OAI21X1
XOAI21X1_1724 BUFX4_148/Y BUFX4_65/Y BUFX2_774/A gnd OAI21X1_1725/C vdd OAI21X1
XFILL_0_OAI21X1_75 gnd vdd FILL
XOAI21X1_1702 BUFX4_93/Y BUFX4_362/Y BUFX2_734/A gnd OAI21X1_1703/C vdd OAI21X1
XOAI21X1_1757 INVX2_140/Y BUFX4_293/Y OAI21X1_1757/C gnd DFFPOSX1_91/D vdd OAI21X1
XFILL_0_OAI21X1_97 gnd vdd FILL
XOAI21X1_1746 BUFX4_125/Y BUFX4_81/Y BUFX2_755/A gnd OAI21X1_1747/C vdd OAI21X1
XFILL_0_OAI21X1_86 gnd vdd FILL
XOAI21X1_1735 INVX2_129/Y BUFX4_296/Y OAI21X1_1735/C gnd DFFPOSX1_80/D vdd OAI21X1
XFILL_0_OAI21X1_702 gnd vdd FILL
XOAI21X1_1768 BUFX4_162/Y BUFX4_38/Y BUFX2_767/A gnd OAI21X1_1769/C vdd OAI21X1
XFILL_0_OAI21X1_713 gnd vdd FILL
XOAI21X1_1779 BUFX4_374/Y INVX2_151/Y NAND2X1_720/Y gnd OAI21X1_1779/Y vdd OAI21X1
XFILL_1_OAI21X1_928 gnd vdd FILL
XFILL_0_OAI21X1_757 gnd vdd FILL
XFILL_0_OAI21X1_746 gnd vdd FILL
XFILL_0_OAI21X1_735 gnd vdd FILL
XFILL_0_OAI21X1_724 gnd vdd FILL
XFILL_1_OAI21X1_906 gnd vdd FILL
XFILL_1_OAI21X1_917 gnd vdd FILL
XFILL_0_OAI21X1_768 gnd vdd FILL
XFILL_0_OAI21X1_779 gnd vdd FILL
XFILL_1_OAI21X1_939 gnd vdd FILL
XFILL_2_NAND3X1_29 gnd vdd FILL
XFILL_3_15_0 gnd vdd FILL
XFILL_0_NAND2X1_741 gnd vdd FILL
XFILL_0_NAND2X1_730 gnd vdd FILL
XFILL_0_NAND2X1_752 gnd vdd FILL
XFILL_0_NAND2X1_763 gnd vdd FILL
XFILL_0_OAI21X1_1523 gnd vdd FILL
XFILL_0_OAI21X1_1512 gnd vdd FILL
XFILL_0_OAI21X1_1534 gnd vdd FILL
XFILL_0_OAI21X1_1501 gnd vdd FILL
XFILL_0_OAI21X1_1567 gnd vdd FILL
XFILL_2_DFFPOSX1_290 gnd vdd FILL
XFILL_0_OAI21X1_1556 gnd vdd FILL
XFILL_0_OAI21X1_1545 gnd vdd FILL
XFILL_0_OAI21X1_1589 gnd vdd FILL
XFILL_5_DFFPOSX1_90 gnd vdd FILL
XFILL_23_4_1 gnd vdd FILL
XFILL_0_OAI21X1_1578 gnd vdd FILL
XFILL_5_DFFPOSX1_761 gnd vdd FILL
XFILL_5_DFFPOSX1_750 gnd vdd FILL
XFILL_5_DFFPOSX1_772 gnd vdd FILL
XFILL_5_DFFPOSX1_783 gnd vdd FILL
XFILL_5_DFFPOSX1_794 gnd vdd FILL
XFILL_8_14_0 gnd vdd FILL
XBUFX4_108 BUFX4_10/A gnd BUFX4_108/Y vdd BUFX4
XBUFX4_119 INVX8_4/Y gnd BUFX4_385/A vdd BUFX4
XFILL_5_0_0 gnd vdd FILL
XFILL_6_5_1 gnd vdd FILL
XFILL_4_DFFPOSX1_340 gnd vdd FILL
XFILL_0_INVX1_19 gnd vdd FILL
XFILL_4_DFFPOSX1_373 gnd vdd FILL
XFILL_4_DFFPOSX1_362 gnd vdd FILL
XFILL_4_DFFPOSX1_351 gnd vdd FILL
XFILL_2_DFFPOSX1_1032 gnd vdd FILL
XFILL_2_DFFPOSX1_1021 gnd vdd FILL
XFILL_4_DFFPOSX1_395 gnd vdd FILL
XFILL_12_12_1 gnd vdd FILL
XFILL_4_DFFPOSX1_384 gnd vdd FILL
XFILL_2_DFFPOSX1_1010 gnd vdd FILL
XFILL_14_4_1 gnd vdd FILL
XFILL_1_BUFX2_252 gnd vdd FILL
XFILL_1_BUFX2_263 gnd vdd FILL
XFILL_1_BUFX2_296 gnd vdd FILL
XOAI21X1_1009 BUFX4_302/Y INVX1_159/Y OAI21X1_1009/C gnd OAI21X1_1009/Y vdd OAI21X1
XOAI21X1_291 INVX2_191/Y BUFX4_291/Y OAI21X1_291/C gnd OAI21X1_291/Y vdd OAI21X1
XFILL_1_OAI21X1_1229 gnd vdd FILL
XFILL_1_OAI21X1_1218 gnd vdd FILL
XFILL_1_OAI21X1_1207 gnd vdd FILL
XOAI21X1_280 BUFX4_124/Y BUFX4_40/Y BUFX2_1004/A gnd OAI21X1_281/C vdd OAI21X1
XFILL_1_DFFPOSX1_808 gnd vdd FILL
XFILL_1_DFFPOSX1_819 gnd vdd FILL
XFILL_6_DFFPOSX1_401 gnd vdd FILL
XFILL_6_DFFPOSX1_412 gnd vdd FILL
XFILL_6_DFFPOSX1_423 gnd vdd FILL
XFILL_6_DFFPOSX1_434 gnd vdd FILL
XFILL_6_DFFPOSX1_445 gnd vdd FILL
XFILL_17_11_1 gnd vdd FILL
XFILL_30_13_1 gnd vdd FILL
XFILL_1_NAND2X1_219 gnd vdd FILL
XFILL_1_NAND3X1_4 gnd vdd FILL
XFILL_36_2 gnd vdd FILL
XFILL_0_DFFPOSX1_409 gnd vdd FILL
XFILL_29_1 gnd vdd FILL
XFILL_5_DFFPOSX1_1014 gnd vdd FILL
XFILL_5_DFFPOSX1_1025 gnd vdd FILL
XFILL_5_DFFPOSX1_1003 gnd vdd FILL
XDFFPOSX1_36 BUFX2_713/A CLKBUF1_86/Y DFFPOSX1_36/D gnd vdd DFFPOSX1
XOAI21X1_1532 BUFX4_170/Y BUFX4_32/Y BUFX2_237/A gnd OAI21X1_1533/C vdd OAI21X1
XDFFPOSX1_25 BUFX2_695/A CLKBUF1_64/Y DFFPOSX1_25/D gnd vdd DFFPOSX1
XDFFPOSX1_14 BUFX2_683/A CLKBUF1_42/Y DFFPOSX1_14/D gnd vdd DFFPOSX1
XOAI21X1_1521 OAI21X1_1521/A BUFX4_297/Y OAI21X1_1521/C gnd OAI21X1_1521/Y vdd OAI21X1
XFILL_0_BUFX4_360 gnd vdd FILL
XOAI21X1_1510 INVX1_223/A INVX1_224/A INVX2_80/Y gnd NAND2X1_639/A vdd OAI21X1
XDFFPOSX1_69 BUFX2_746/A CLKBUF1_74/Y DFFPOSX1_69/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1730 gnd vdd FILL
XDFFPOSX1_58 BUFX2_728/A CLKBUF1_16/Y DFFPOSX1_58/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1741 gnd vdd FILL
XFILL_0_BUFX4_382 gnd vdd FILL
XFILL_1_OAI21X1_1752 gnd vdd FILL
XDFFPOSX1_47 BUFX2_716/A CLKBUF1_64/Y DFFPOSX1_47/D gnd vdd DFFPOSX1
XOAI21X1_1565 OR2X2_21/Y NOR2X1_176/B BUFX4_284/Y gnd OAI21X1_1566/B vdd OAI21X1
XFILL_0_BUFX4_371 gnd vdd FILL
XOAI21X1_1543 OR2X2_21/A INVX1_196/A INVX2_86/Y gnd OAI21X1_1544/C vdd OAI21X1
XOAI21X1_1554 INVX1_226/A INVX2_104/Y BUFX4_286/Y gnd OAI21X1_1555/B vdd OAI21X1
XFILL_1_OAI21X1_1785 gnd vdd FILL
XFILL_1_OAI21X1_1763 gnd vdd FILL
XOAI21X1_1598 BUFX4_318/Y INVX2_134/Y NAND2X1_667/Y gnd OAI21X1_1598/Y vdd OAI21X1
XFILL_1_OAI21X1_1774 gnd vdd FILL
XOAI21X1_1576 INVX2_113/Y BUFX4_213/Y NAND2X1_649/Y gnd OAI21X1_1576/Y vdd OAI21X1
XFILL_1_OAI21X1_703 gnd vdd FILL
XFILL_0_OAI21X1_510 gnd vdd FILL
XOAI21X1_1587 OAI21X1_6/A INVX2_123/Y NAND2X1_656/Y gnd OAI21X1_1587/Y vdd OAI21X1
XFILL_0_OAI21X1_521 gnd vdd FILL
XFILL_2_OAI21X1_907 gnd vdd FILL
XFILL_1_OAI21X1_1796 gnd vdd FILL
XFILL_1_OAI21X1_714 gnd vdd FILL
XFILL_0_OAI21X1_554 gnd vdd FILL
XFILL_1_OAI21X1_736 gnd vdd FILL
XFILL_0_BUFX2_1020 gnd vdd FILL
XFILL_0_OAI21X1_543 gnd vdd FILL
XFILL_0_BUFX2_1031 gnd vdd FILL
XFILL_1_OAI21X1_725 gnd vdd FILL
XFILL_0_OAI21X1_565 gnd vdd FILL
XFILL_0_OAI21X1_532 gnd vdd FILL
XFILL_1_OAI21X1_758 gnd vdd FILL
XFILL_1_OAI21X1_769 gnd vdd FILL
XFILL_0_OAI21X1_576 gnd vdd FILL
XFILL_1_OAI21X1_747 gnd vdd FILL
XFILL_0_OAI21X1_598 gnd vdd FILL
XFILL_0_OAI21X1_587 gnd vdd FILL
XFILL_35_12_1 gnd vdd FILL
XFILL_0_CLKBUF1_21 gnd vdd FILL
XFILL_0_CLKBUF1_10 gnd vdd FILL
XFILL_0_CLKBUF1_32 gnd vdd FILL
XFILL_0_CLKBUF1_43 gnd vdd FILL
XFILL_0_CLKBUF1_54 gnd vdd FILL
XFILL_0_CLKBUF1_65 gnd vdd FILL
XFILL_0_CLKBUF1_87 gnd vdd FILL
XFILL_0_CLKBUF1_76 gnd vdd FILL
XFILL_1_NAND2X1_742 gnd vdd FILL
XFILL_0_CLKBUF1_98 gnd vdd FILL
XFILL_1_NAND2X1_731 gnd vdd FILL
XFILL_0_NAND2X1_560 gnd vdd FILL
XFILL_0_OAI21X1_1342 gnd vdd FILL
XFILL_0_OAI21X1_1331 gnd vdd FILL
XFILL_0_NAND2X1_571 gnd vdd FILL
XFILL_0_OAI21X1_1320 gnd vdd FILL
XFILL_0_DFFPOSX1_910 gnd vdd FILL
XFILL_0_NAND2X1_593 gnd vdd FILL
XFILL_0_DFFPOSX1_943 gnd vdd FILL
XFILL_0_OAI21X1_1375 gnd vdd FILL
XFILL_0_DFFPOSX1_932 gnd vdd FILL
XFILL_0_NAND2X1_582 gnd vdd FILL
XFILL_0_DFFPOSX1_921 gnd vdd FILL
XFILL_0_OAI21X1_1353 gnd vdd FILL
XFILL_0_OAI21X1_1364 gnd vdd FILL
XFILL_0_OAI21X1_1397 gnd vdd FILL
XFILL_0_DFFPOSX1_954 gnd vdd FILL
XFILL_0_OAI21X1_1386 gnd vdd FILL
XFILL_0_DFFPOSX1_965 gnd vdd FILL
XFILL_0_DFFPOSX1_976 gnd vdd FILL
XFILL_6_DFFPOSX1_91 gnd vdd FILL
XFILL_0_DFFPOSX1_998 gnd vdd FILL
XFILL_0_DFFPOSX1_987 gnd vdd FILL
XFILL_5_DFFPOSX1_591 gnd vdd FILL
XFILL_5_DFFPOSX1_580 gnd vdd FILL
XFILL_0_OR2X2_4 gnd vdd FILL
XFILL_0_BUFX2_308 gnd vdd FILL
XINVX2_119 bundlePid_i[29] gnd INVX2_119/Y vdd INVX2
XINVX2_108 INVX2_108/A gnd INVX2_108/Y vdd INVX2
XFILL_0_BUFX2_319 gnd vdd FILL
XFILL_1_BUFX4_2 gnd vdd FILL
XFILL_4_DFFPOSX1_181 gnd vdd FILL
XFILL_2_OAI21X1_1425 gnd vdd FILL
XFILL_4_DFFPOSX1_170 gnd vdd FILL
XFILL_2_NOR3X1_14 gnd vdd FILL
XFILL_2_OAI21X1_1469 gnd vdd FILL
XFILL_4_DFFPOSX1_192 gnd vdd FILL
XFILL_2_BUFX4_280 gnd vdd FILL
XFILL_0_INVX1_6 gnd vdd FILL
XFILL_2_BUFX4_291 gnd vdd FILL
XFILL_1_NAND3X1_26 gnd vdd FILL
XFILL_1_NAND3X1_37 gnd vdd FILL
XFILL_1_OAI21X1_1004 gnd vdd FILL
XFILL_1_NAND3X1_15 gnd vdd FILL
XFILL_0_BUFX2_820 gnd vdd FILL
XDFFPOSX1_418 BUFX2_452/A CLKBUF1_70/Y OAI21X1_390/Y gnd vdd DFFPOSX1
XDFFPOSX1_407 BUFX2_440/A CLKBUF1_91/Y OAI21X1_379/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_605 gnd vdd FILL
XFILL_1_OAI21X1_1037 gnd vdd FILL
XFILL_1_NAND3X1_59 gnd vdd FILL
XFILL_1_NAND3X1_48 gnd vdd FILL
XFILL_1_OAI21X1_1015 gnd vdd FILL
XFILL_0_BUFX2_842 gnd vdd FILL
XFILL_0_BUFX2_831 gnd vdd FILL
XDFFPOSX1_429 BUFX2_520/A CLKBUF1_13/Y OAI21X1_412/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1026 gnd vdd FILL
XFILL_0_BUFX2_875 gnd vdd FILL
XFILL_1_OAI21X1_1048 gnd vdd FILL
XINVX1_130 bundle_i[74] gnd INVX1_130/Y vdd INVX1
XFILL_1_DFFPOSX1_627 gnd vdd FILL
XFILL_1_DFFPOSX1_616 gnd vdd FILL
XFILL_1_DFFPOSX1_638 gnd vdd FILL
XFILL_0_BUFX2_853 gnd vdd FILL
XINVX1_152 bundle_i[116] gnd INVX1_152/Y vdd INVX1
XINVX1_141 bundle_i[127] gnd INVX1_141/Y vdd INVX1
XFILL_1_OAI21X1_1059 gnd vdd FILL
XFILL_0_BUFX2_864 gnd vdd FILL
XINVX1_185 INVX1_185/A gnd INVX1_185/Y vdd INVX1
XFILL_1_DFFPOSX1_649 gnd vdd FILL
XFILL_0_BUFX2_897 gnd vdd FILL
XFILL_0_BUFX2_886 gnd vdd FILL
XINVX1_163 bundle_i[105] gnd INVX1_163/Y vdd INVX1
XINVX1_174 bundleAddress_i[40] gnd INVX1_174/Y vdd INVX1
XINVX1_196 INVX1_196/A gnd INVX1_196/Y vdd INVX1
XFILL_6_DFFPOSX1_286 gnd vdd FILL
XCLKBUF1_100 BUFX4_85/Y gnd CLKBUF1_100/Y vdd CLKBUF1
XFILL_6_DFFPOSX1_297 gnd vdd FILL
XFILL_37_3_1 gnd vdd FILL
XFILL_0_INVX2_62 gnd vdd FILL
XFILL_0_INVX2_73 gnd vdd FILL
XFILL_0_INVX2_51 gnd vdd FILL
XFILL_0_INVX2_40 gnd vdd FILL
XFILL_0_INVX2_95 gnd vdd FILL
XFILL_0_INVX2_84 gnd vdd FILL
XFILL_1_NOR3X1_4 gnd vdd FILL
XFILL_0_DFFPOSX1_217 gnd vdd FILL
XFILL_0_DFFPOSX1_239 gnd vdd FILL
XFILL_0_DFFPOSX1_228 gnd vdd FILL
XFILL_0_DFFPOSX1_206 gnd vdd FILL
XFILL_20_2_1 gnd vdd FILL
XOAI21X1_1340 INVX1_212/A INVX1_195/A BUFX4_310/Y gnd OAI21X1_1341/B vdd OAI21X1
XFILL_21_18_1 gnd vdd FILL
XDFFPOSX1_941 BUFX2_238/A CLKBUF1_31/Y OAI21X1_1399/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1560 gnd vdd FILL
XOAI21X1_1373 XNOR2X1_88/Y BUFX4_141/Y OAI21X1_1373/C gnd OAI21X1_1373/Y vdd OAI21X1
XOAI21X1_1351 NOR2X1_211/B NOR3X1_12/B BUFX4_308/Y gnd OAI21X1_1352/A vdd OAI21X1
XDFFPOSX1_930 BUFX2_183/A CLKBUF1_28/Y OAI21X1_1371/Y gnd vdd DFFPOSX1
XFILL_0_BUFX4_190 gnd vdd FILL
XOAI21X1_1362 INVX1_215/A INVX4_45/Y INVX2_88/Y gnd OAI21X1_1363/C vdd OAI21X1
XFILL_1_OAI21X1_1582 gnd vdd FILL
XOAI21X1_1384 BUFX4_178/Y BUFX4_50/Y BUFX2_193/A gnd OAI21X1_1385/C vdd OAI21X1
XDFFPOSX1_952 BUFX2_201/A CLKBUF1_23/Y OAI21X1_1433/Y gnd vdd DFFPOSX1
XDFFPOSX1_985 BUFX2_237/A CLKBUF1_86/Y OAI21X1_1533/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1571 gnd vdd FILL
XDFFPOSX1_963 BUFX2_213/A CLKBUF1_49/Y OAI21X1_1462/Y gnd vdd DFFPOSX1
XOAI21X1_1395 OAI21X1_1395/A BUFX4_299/Y OAI21X1_1395/C gnd OAI21X1_1395/Y vdd OAI21X1
XFILL_1_OAI21X1_1593 gnd vdd FILL
XFILL_1_OAI21X1_500 gnd vdd FILL
XFILL_1_NOR2X1_105 gnd vdd FILL
XFILL_0_OAI21X1_340 gnd vdd FILL
XFILL_1_OAI21X1_511 gnd vdd FILL
XDFFPOSX1_974 BUFX2_225/A CLKBUF1_28/Y OAI21X1_1499/Y gnd vdd DFFPOSX1
XFILL_1_NOR2X1_127 gnd vdd FILL
XDFFPOSX1_996 BUFX2_250/A CLKBUF1_40/Y OAI21X1_1566/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_373 gnd vdd FILL
XFILL_1_OAI21X1_533 gnd vdd FILL
XFILL_1_OAI21X1_544 gnd vdd FILL
XFILL_0_OAI21X1_351 gnd vdd FILL
XFILL_0_OAI21X1_362 gnd vdd FILL
XFILL_1_OAI21X1_522 gnd vdd FILL
XFILL_1_NOR2X1_138 gnd vdd FILL
XFILL_1_NOR2X1_149 gnd vdd FILL
XFILL_0_OAI21X1_384 gnd vdd FILL
XFILL_1_OAI21X1_566 gnd vdd FILL
XFILL_1_OAI21X1_555 gnd vdd FILL
XFILL_1_OAI21X1_577 gnd vdd FILL
XFILL_0_OAI21X1_395 gnd vdd FILL
XFILL_2_OAI21X1_726 gnd vdd FILL
XFILL_1_OAI21X1_599 gnd vdd FILL
XFILL_1_OAI21X1_588 gnd vdd FILL
XFILL_1_OAI21X1_1 gnd vdd FILL
XFILL_28_3_1 gnd vdd FILL
XBUFX2_409 BUFX2_409/A gnd majID1_o[40] vdd BUFX2
XFILL_3_3_1 gnd vdd FILL
XFILL_0_OAI21X1_1150 gnd vdd FILL
XFILL_1_BUFX4_303 gnd vdd FILL
XFILL_0_DFFPOSX1_751 gnd vdd FILL
XFILL_1_BUFX4_336 gnd vdd FILL
XFILL_0_DFFPOSX1_740 gnd vdd FILL
XFILL_0_NAND2X1_390 gnd vdd FILL
XFILL_1_BUFX4_347 gnd vdd FILL
XFILL_1_NAND2X1_561 gnd vdd FILL
XFILL_0_OAI21X1_1172 gnd vdd FILL
XFILL_1_BUFX4_325 gnd vdd FILL
XFILL_0_OAI21X1_1161 gnd vdd FILL
XFILL_1_BUFX4_314 gnd vdd FILL
XFILL_0_OAI21X1_1183 gnd vdd FILL
XFILL_0_DFFPOSX1_773 gnd vdd FILL
XFILL_26_17_1 gnd vdd FILL
XFILL_0_DFFPOSX1_762 gnd vdd FILL
XFILL_1_BUFX4_358 gnd vdd FILL
XFILL_0_OAI21X1_1194 gnd vdd FILL
XFILL_1_BUFX4_369 gnd vdd FILL
XFILL_0_DFFPOSX1_784 gnd vdd FILL
XFILL_11_2_1 gnd vdd FILL
XFILL_0_DFFPOSX1_795 gnd vdd FILL
XFILL_0_BUFX2_138 gnd vdd FILL
XFILL_0_BUFX2_127 gnd vdd FILL
XFILL_0_BUFX2_105 gnd vdd FILL
XFILL_0_BUFX2_116 gnd vdd FILL
XFILL_0_BUFX2_149 gnd vdd FILL
XFILL_20_13_0 gnd vdd FILL
XFILL_1_NAND2X1_70 gnd vdd FILL
XFILL_1_NAND2X1_81 gnd vdd FILL
XBUFX2_921 BUFX2_921/A gnd tid3_o[40] vdd BUFX2
XFILL_2_DFFPOSX1_812 gnd vdd FILL
XFILL_2_DFFPOSX1_823 gnd vdd FILL
XFILL_2_OAI21X1_1244 gnd vdd FILL
XFILL_19_3_1 gnd vdd FILL
XBUFX2_910 BUFX2_910/A gnd tid3_o[50] vdd BUFX2
XFILL_2_DFFPOSX1_801 gnd vdd FILL
XBUFX2_943 BUFX2_943/A gnd tid3_o[20] vdd BUFX2
XBUFX2_932 BUFX2_932/A gnd tid3_o[30] vdd BUFX2
XBUFX2_954 BUFX2_954/A gnd tid3_o[10] vdd BUFX2
XFILL_2_DFFPOSX1_856 gnd vdd FILL
XFILL_2_DFFPOSX1_834 gnd vdd FILL
XFILL_2_OAI21X1_1299 gnd vdd FILL
XBUFX2_965 BUFX2_965/A gnd tid3_o[0] vdd BUFX2
XFILL_2_DFFPOSX1_845 gnd vdd FILL
XFILL_2_OAI21X1_1266 gnd vdd FILL
XFILL_1_18_1 gnd vdd FILL
XBUFX2_987 BUFX2_987/A gnd tid4_o[38] vdd BUFX2
XBUFX2_976 BUFX2_976/A gnd tid4_o[48] vdd BUFX2
XFILL_2_DFFPOSX1_889 gnd vdd FILL
XFILL_2_DFFPOSX1_878 gnd vdd FILL
XBUFX2_998 BUFX2_998/A gnd tid4_o[28] vdd BUFX2
XFILL_2_DFFPOSX1_867 gnd vdd FILL
XFILL_25_12_0 gnd vdd FILL
XDFFPOSX1_204 BUFX2_876/A CLKBUF1_2/Y OAI21X1_48/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_650 gnd vdd FILL
XDFFPOSX1_237 BUFX2_968/A CLKBUF1_65/Y OAI21X1_91/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_413 gnd vdd FILL
XDFFPOSX1_215 BUFX2_888/A CLKBUF1_26/Y OAI21X1_59/Y gnd vdd DFFPOSX1
XFILL_2_AOI21X1_7 gnd vdd FILL
XFILL_1_DFFPOSX1_402 gnd vdd FILL
XDFFPOSX1_226 BUFX2_900/A CLKBUF1_41/Y OAI21X1_70/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_661 gnd vdd FILL
XFILL_0_BUFX2_672 gnd vdd FILL
XDFFPOSX1_248 BUFX2_918/A CLKBUF1_70/Y OAI21X1_113/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_694 gnd vdd FILL
XDFFPOSX1_259 BUFX2_930/A CLKBUF1_78/Y OAI21X1_135/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_457 gnd vdd FILL
XFILL_0_BUFX2_683 gnd vdd FILL
XFILL_1_DFFPOSX1_424 gnd vdd FILL
XFILL_1_DFFPOSX1_435 gnd vdd FILL
XFILL_1_DFFPOSX1_446 gnd vdd FILL
XNAND2X1_307 BUFX4_305/Y OAI21X1_656/A gnd OAI21X1_651/B vdd NAND2X1
XFILL_1_DFFPOSX1_479 gnd vdd FILL
XFILL_1_DFFPOSX1_468 gnd vdd FILL
XNAND2X1_318 AND2X2_18/Y AND2X2_2/Y gnd NOR3X1_9/A vdd NAND2X1
XNAND2X1_329 AND2X2_22/A OAI21X1_787/Y gnd OAI21X1_789/A vdd NAND2X1
XFILL_4_DFFPOSX1_906 gnd vdd FILL
XFILL_4_DFFPOSX1_917 gnd vdd FILL
XFILL_6_17_1 gnd vdd FILL
XFILL_4_DFFPOSX1_928 gnd vdd FILL
XFILL_4_DFFPOSX1_939 gnd vdd FILL
XNOR3X1_14 INVX2_87/Y INVX4_48/Y NOR3X1_14/C gnd NOR3X1_14/Y vdd NOR3X1
XBUFX4_291 BUFX4_303/A gnd BUFX4_291/Y vdd BUFX4
XBUFX4_280 INVX8_7/Y gnd BUFX4_80/A vdd BUFX4
XFILL_0_13_0 gnd vdd FILL
XFILL_0_INVX2_190 gnd vdd FILL
XFILL_0_XNOR2X1_6 gnd vdd FILL
XFILL_1_BUFX2_829 gnd vdd FILL
XOAI21X1_813 OAI21X1_813/A BUFX4_289/Y OAI21X1_813/C gnd OAI21X1_813/Y vdd OAI21X1
XOAI21X1_824 OAI21X1_824/A BUFX4_295/Y OAI21X1_824/C gnd OAI21X1_824/Y vdd OAI21X1
XOAI21X1_802 INVX2_53/Y INVX4_23/Y INVX2_33/Y gnd OAI21X1_803/C vdd OAI21X1
XOAI21X1_835 BUFX4_156/Y BUFX4_70/Y BUFX2_643/A gnd OAI21X1_837/C vdd OAI21X1
XFILL_3_DFFPOSX1_529 gnd vdd FILL
XOAI21X1_857 INVX1_58/Y BUFX4_261/Y OAI21X1_857/C gnd OAI21X1_857/Y vdd OAI21X1
XOAI21X1_846 INVX1_47/Y BUFX4_267/Y OAI21X1_846/C gnd OAI21X1_846/Y vdd OAI21X1
XFILL_3_DFFPOSX1_507 gnd vdd FILL
XFILL_3_DFFPOSX1_518 gnd vdd FILL
XOAI21X1_879 INVX1_80/Y BUFX4_205/Y OAI21X1_879/C gnd OAI21X1_879/Y vdd OAI21X1
XOAI21X1_868 INVX1_69/Y BUFX4_267/Y OAI21X1_868/C gnd OAI21X1_868/Y vdd OAI21X1
XOAI21X1_1170 XNOR2X1_72/Y BUFX4_202/Y NAND2X1_551/Y gnd OAI21X1_1170/Y vdd OAI21X1
XOAI21X1_1181 NOR2X1_167/Y OAI21X1_1181/B NAND2X1_567/Y gnd OAI21X1_1181/Y vdd OAI21X1
XOAI21X1_1192 NAND3X1_48/Y INVX2_104/Y BUFX4_242/Y gnd OAI21X1_1193/A vdd OAI21X1
XFILL_1_OAI21X1_1390 gnd vdd FILL
XDFFPOSX1_771 BUFX2_21/A CLKBUF1_55/Y OAI21X1_1063/Y gnd vdd DFFPOSX1
XDFFPOSX1_760 BUFX2_9/A CLKBUF1_23/Y OAI21X1_1052/Y gnd vdd DFFPOSX1
XDFFPOSX1_793 BUFX2_45/A CLKBUF1_68/Y OAI21X1_1085/Y gnd vdd DFFPOSX1
XDFFPOSX1_782 BUFX2_33/A CLKBUF1_53/Y OAI21X1_1074/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_181 gnd vdd FILL
XFILL_1_DFFPOSX1_980 gnd vdd FILL
XFILL_0_OAI21X1_170 gnd vdd FILL
XFILL_1_OAI21X1_330 gnd vdd FILL
XFILL_1_OAI21X1_341 gnd vdd FILL
XFILL_1_OAI21X1_352 gnd vdd FILL
XFILL_1_DFFPOSX1_991 gnd vdd FILL
XFILL_1_OAI21X1_385 gnd vdd FILL
XFILL_1_OAI21X1_396 gnd vdd FILL
XFILL_1_OAI21X1_374 gnd vdd FILL
XFILL_1_OAI21X1_363 gnd vdd FILL
XFILL_0_OAI21X1_192 gnd vdd FILL
XFILL_1_CLKBUF1_6 gnd vdd FILL
XFILL_5_12_0 gnd vdd FILL
XBUFX2_217 BUFX2_217/A gnd addr4_o[33] vdd BUFX2
XFILL_2_DFFPOSX1_119 gnd vdd FILL
XFILL_0_NAND3X1_12 gnd vdd FILL
XFILL_0_NAND3X1_45 gnd vdd FILL
XFILL_0_NAND3X1_34 gnd vdd FILL
XFILL_0_NAND3X1_23 gnd vdd FILL
XBUFX2_206 BUFX2_206/A gnd addr4_o[43] vdd BUFX2
XFILL_2_DFFPOSX1_108 gnd vdd FILL
XFILL_0_NAND3X1_56 gnd vdd FILL
XFILL_0_NAND3X1_67 gnd vdd FILL
XBUFX2_239 BUFX2_239/A gnd addr4_o[13] vdd BUFX2
XBUFX2_228 BUFX2_228/A gnd addr4_o[23] vdd BUFX2
XFILL_0_BUFX4_80 gnd vdd FILL
XFILL_1_BUFX4_100 gnd vdd FILL
XFILL_0_BUFX4_91 gnd vdd FILL
XFILL_1_BUFX4_111 gnd vdd FILL
XFILL_1_BUFX4_155 gnd vdd FILL
XFILL_1_BUFX4_133 gnd vdd FILL
XFILL_1_BUFX4_122 gnd vdd FILL
XFILL_1_BUFX4_144 gnd vdd FILL
XFILL_1_NAND2X1_391 gnd vdd FILL
XFILL_1_NAND2X1_380 gnd vdd FILL
XFILL_1_BUFX4_166 gnd vdd FILL
XFILL_0_DFFPOSX1_592 gnd vdd FILL
XFILL_1_BUFX4_177 gnd vdd FILL
XFILL_1_BUFX4_188 gnd vdd FILL
XFILL_0_DFFPOSX1_570 gnd vdd FILL
XFILL_0_DFFPOSX1_581 gnd vdd FILL
XFILL_1_BUFX4_199 gnd vdd FILL
XFILL_1_MUX2X1_2 gnd vdd FILL
XFILL_2_CLKBUF1_39 gnd vdd FILL
XFILL_2_CLKBUF1_17 gnd vdd FILL
XFILL_2_CLKBUF1_28 gnd vdd FILL
XFILL_11_18_0 gnd vdd FILL
XFILL_2_DFFPOSX1_620 gnd vdd FILL
XFILL_2_DFFPOSX1_631 gnd vdd FILL
XFILL_2_OAI21X1_1074 gnd vdd FILL
XFILL_2_DFFPOSX1_664 gnd vdd FILL
XFILL_34_1_1 gnd vdd FILL
XBUFX2_762 BUFX2_762/A gnd pid4_o[7] vdd BUFX2
XBUFX2_751 BUFX2_751/A gnd pid4_o[17] vdd BUFX2
XFILL_2_DFFPOSX1_642 gnd vdd FILL
XFILL_2_OAI21X1_1085 gnd vdd FILL
XNOR2X1_80 INVX2_48/Y OR2X2_10/Y gnd NOR2X1_80/Y vdd NOR2X1
XNOR2X1_91 INVX1_31/A NOR2X1_91/B gnd NOR2X1_91/Y vdd NOR2X1
XFILL_2_DFFPOSX1_675 gnd vdd FILL
XFILL_2_DFFPOSX1_653 gnd vdd FILL
XBUFX2_740 BUFX2_740/A gnd pid3_o[26] vdd BUFX2
XBUFX2_773 BUFX2_773/A gnd pid4_o[25] vdd BUFX2
XBUFX2_795 BUFX2_795/A gnd tid1_o[38] vdd BUFX2
XBUFX2_784 BUFX2_784/A gnd tid1_o[48] vdd BUFX2
XFILL_0_NOR2X1_113 gnd vdd FILL
XFILL_2_DFFPOSX1_697 gnd vdd FILL
XFILL_2_DFFPOSX1_686 gnd vdd FILL
XFILL_0_NOR2X1_102 gnd vdd FILL
XFILL_0_NOR2X1_124 gnd vdd FILL
XFILL_0_NOR2X1_146 gnd vdd FILL
XFILL_0_NOR2X1_135 gnd vdd FILL
XFILL_0_NOR2X1_179 gnd vdd FILL
XOAI21X1_109 BUFX4_138/Y INVX2_164/Y OAI21X1_109/C gnd OAI21X1_109/Y vdd OAI21X1
XFILL_0_NOR2X1_168 gnd vdd FILL
XFILL_11_1 gnd vdd FILL
XFILL_0_NOR2X1_157 gnd vdd FILL
XFILL_0_DFFPOSX1_1009 gnd vdd FILL
XBUFX2_7 BUFX2_7/A gnd addr1_o[49] vdd BUFX2
XFILL_1_DFFPOSX1_232 gnd vdd FILL
XFILL_1_DFFPOSX1_221 gnd vdd FILL
XFILL_1_DFFPOSX1_210 gnd vdd FILL
XFILL_1_DFFPOSX1_254 gnd vdd FILL
XFILL_1_DFFPOSX1_243 gnd vdd FILL
XFILL_1_DFFPOSX1_265 gnd vdd FILL
XFILL_0_BUFX2_480 gnd vdd FILL
XFILL_0_BUFX2_491 gnd vdd FILL
XFILL_1_DFFPOSX1_276 gnd vdd FILL
XNAND2X1_115 BUFX2_431/A BUFX4_325/Y gnd OAI21X1_371/C vdd NAND2X1
XFILL_1_DFFPOSX1_298 gnd vdd FILL
XNAND2X1_104 BUFX2_419/A BUFX4_346/Y gnd OAI21X1_360/C vdd NAND2X1
XNAND2X1_126 BUFX2_443/A BUFX4_346/Y gnd OAI21X1_382/C vdd NAND2X1
XFILL_1_DFFPOSX1_287 gnd vdd FILL
XNAND2X1_137 bundleStartMajId_i[63] bundleStartMajId_i[62] gnd INVX1_7/A vdd NAND2X1
XNAND2X1_148 BUFX2_513/A BUFX4_199/Y gnd OAI21X1_407/C vdd NAND2X1
XFILL_4_DFFPOSX1_703 gnd vdd FILL
XNAND2X1_159 bundleStartMajId_i[52] bundleStartMajId_i[51] gnd OR2X2_1/B vdd NAND2X1
XFILL_4_DFFPOSX1_747 gnd vdd FILL
XFILL_4_DFFPOSX1_725 gnd vdd FILL
XFILL_1_OAI21X1_24 gnd vdd FILL
XFILL_4_DFFPOSX1_736 gnd vdd FILL
XFILL_4_DFFPOSX1_714 gnd vdd FILL
XFILL_16_17_0 gnd vdd FILL
XNAND2X1_2 NAND2X1_2/A OAI21X1_2/A gnd OAI21X1_2/C vdd NAND2X1
XFILL_1_OAI21X1_13 gnd vdd FILL
XFILL_1_OAI21X1_35 gnd vdd FILL
XFILL_1_OAI21X1_46 gnd vdd FILL
XFILL_32_10_1 gnd vdd FILL
XFILL_4_DFFPOSX1_758 gnd vdd FILL
XFILL_1_OAI21X1_57 gnd vdd FILL
XFILL_4_DFFPOSX1_769 gnd vdd FILL
XFILL_1_OAI21X1_79 gnd vdd FILL
XFILL_1_OAI21X1_68 gnd vdd FILL
XFILL_25_1_1 gnd vdd FILL
XFILL_0_1_1 gnd vdd FILL
XNOR2X1_170 bundleAddress_i[8] NOR3X1_14/Y gnd NOR2X1_170/Y vdd NOR2X1
XNOR2X1_181 NOR2X1_185/A INVX1_201/A gnd INVX1_200/A vdd NOR2X1
XNOR2X1_192 INVX1_205/Y NOR3X1_18/C gnd AND2X2_29/A vdd NOR2X1
XFILL_1_BUFX2_637 gnd vdd FILL
XFILL_1_BUFX2_604 gnd vdd FILL
XINVX2_7 bundleTid_i[0] gnd INVX2_7/Y vdd INVX2
XFILL_1_BUFX2_626 gnd vdd FILL
XFILL_3_DFFPOSX1_304 gnd vdd FILL
XOAI21X1_632 NOR2X1_97/B OR2X2_13/B NOR2X1_96/B gnd OAI21X1_633/B vdd OAI21X1
XOAI21X1_610 OAI21X1_610/A INVX4_21/Y NOR2X1_96/B gnd OAI21X1_611/B vdd OAI21X1
XOAI21X1_621 BUFX4_107/Y BUFX4_372/Y BUFX2_563/A gnd OAI21X1_623/C vdd OAI21X1
XFILL_1_BUFX2_648 gnd vdd FILL
XFILL_3_DFFPOSX1_337 gnd vdd FILL
XFILL_3_DFFPOSX1_326 gnd vdd FILL
XFILL_3_DFFPOSX1_315 gnd vdd FILL
XOAI21X1_654 NOR2X1_100/Y OAI21X1_654/B OAI21X1_654/C gnd OAI21X1_654/Y vdd OAI21X1
XOAI21X1_643 OAI21X1_643/A BUFX4_146/Y OAI21X1_643/C gnd OAI21X1_643/Y vdd OAI21X1
XAOI21X1_7 bundleStartMajId_i[34] NOR2X1_72/Y bundleStartMajId_i[33] gnd AOI21X1_7/Y
+ vdd AOI21X1
XOAI21X1_665 OAI21X1_665/A BUFX4_302/Y OAI21X1_665/C gnd OAI21X1_665/Y vdd OAI21X1
XFILL_3_DFFPOSX1_348 gnd vdd FILL
XFILL_3_DFFPOSX1_359 gnd vdd FILL
XOAI21X1_687 BUFX4_167/Y BUFX4_82/A BUFX2_587/A gnd OAI21X1_688/C vdd OAI21X1
XOAI21X1_676 INVX1_34/A bundleStartMajId_i[57] BUFX4_285/Y gnd OAI21X1_678/B vdd OAI21X1
XOAI21X1_698 AND2X2_20/Y bundleStartMajId_i[49] OAI21X1_698/C gnd OAI21X1_700/A vdd
+ OAI21X1
XFILL_6_DFFPOSX1_819 gnd vdd FILL
XFILL_0_INVX4_19 gnd vdd FILL
XDFFPOSX1_590 BUFX2_622/A CLKBUF1_80/Y OAI21X1_778/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_160 gnd vdd FILL
XXNOR2X1_15 NOR2X1_33/B INVX4_17/Y gnd XNOR2X1_15/Y vdd XNOR2X1
XXNOR2X1_37 NOR2X1_97/B INVX4_23/Y gnd XNOR2X1_37/Y vdd XNOR2X1
XFILL_1_OAI21X1_171 gnd vdd FILL
XXNOR2X1_48 NOR3X1_7/C NOR3X1_7/A gnd XNOR2X1_48/Y vdd XNOR2X1
XXNOR2X1_26 OAI22X1_1/B INVX4_5/Y gnd XNOR2X1_26/Y vdd XNOR2X1
XFILL_8_2_1 gnd vdd FILL
XFILL_34_18_0 gnd vdd FILL
XNAND2X1_682 BUFX2_681/A BUFX4_234/Y gnd NAND2X1_682/Y vdd NAND2X1
XNAND2X1_660 BUFX2_651/A BUFX4_349/Y gnd NAND2X1_660/Y vdd NAND2X1
XXNOR2X1_59 XNOR2X1_59/A bundleAddress_i[46] gnd XNOR2X1_59/Y vdd XNOR2X1
XNAND2X1_671 BUFX2_663/A BUFX4_366/Y gnd NAND2X1_671/Y vdd NAND2X1
XINVX1_50 INVX1_50/A gnd INVX1_50/Y vdd INVX1
XFILL_1_OAI21X1_182 gnd vdd FILL
XFILL_1_OAI21X1_193 gnd vdd FILL
XINVX1_61 INVX1_61/A gnd INVX1_61/Y vdd INVX1
XNAND2X1_693 BUFX2_684/A BUFX4_211/Y gnd NAND2X1_693/Y vdd NAND2X1
XINVX1_83 bundle_i[57] gnd INVX1_83/Y vdd INVX1
XINVX1_72 INVX1_72/A gnd INVX1_72/Y vdd INVX1
XINVX1_94 bundle_i[46] gnd INVX1_94/Y vdd INVX1
XBUFX2_25 BUFX2_25/A gnd addr1_o[33] vdd BUFX2
XBUFX2_36 BUFX2_36/A gnd addr1_o[23] vdd BUFX2
XBUFX2_14 BUFX2_14/A gnd addr1_o[43] vdd BUFX2
XBUFX2_69 BUFX2_69/A gnd addr2_o[51] vdd BUFX2
XBUFX2_58 BUFX2_58/A gnd addr1_o[3] vdd BUFX2
XDFFPOSX1_2 BUFX2_673/A CLKBUF1_92/Y DFFPOSX1_2/D gnd vdd DFFPOSX1
XBUFX2_47 BUFX2_47/A gnd addr1_o[13] vdd BUFX2
XFILL_16_1_1 gnd vdd FILL
XFILL_5_DFFPOSX1_409 gnd vdd FILL
XFILL_1_BUFX4_36 gnd vdd FILL
XFILL_1_BUFX4_14 gnd vdd FILL
XFILL_1_BUFX4_25 gnd vdd FILL
XFILL_1_BUFX4_47 gnd vdd FILL
XFILL_1_BUFX4_69 gnd vdd FILL
XFILL_1_BUFX4_58 gnd vdd FILL
XFILL_3_DFFPOSX1_882 gnd vdd FILL
XFILL_3_DFFPOSX1_871 gnd vdd FILL
XFILL_3_DFFPOSX1_893 gnd vdd FILL
XFILL_0_OAI21X1_906 gnd vdd FILL
XNOR2X1_5 NOR2X1_5/A NOR2X1_5/B gnd NOR2X1_5/Y vdd NOR2X1
XFILL_3_DFFPOSX1_860 gnd vdd FILL
XFILL_0_OAI21X1_928 gnd vdd FILL
XFILL_0_OAI21X1_939 gnd vdd FILL
XFILL_0_OAI21X1_917 gnd vdd FILL
XFILL_36_9_0 gnd vdd FILL
XFILL_2_DFFPOSX1_450 gnd vdd FILL
XFILL_0_OAI21X1_1716 gnd vdd FILL
XFILL_0_OAI21X1_1705 gnd vdd FILL
XFILL_1_OR2X2_17 gnd vdd FILL
XFILL_0_OAI21X1_1727 gnd vdd FILL
XFILL_2_DFFPOSX1_483 gnd vdd FILL
XBUFX2_581 BUFX2_581/A gnd majID3_o[0] vdd BUFX2
XFILL_0_OAI21X1_1738 gnd vdd FILL
XBUFX2_570 BUFX2_570/A gnd majID3_o[10] vdd BUFX2
XFILL_0_OAI21X1_1749 gnd vdd FILL
XFILL_2_DFFPOSX1_461 gnd vdd FILL
XFILL_2_DFFPOSX1_472 gnd vdd FILL
XFILL_4_DFFPOSX1_90 gnd vdd FILL
XBUFX2_592 BUFX2_592/A gnd majID4_o[48] vdd BUFX2
XFILL_2_DFFPOSX1_494 gnd vdd FILL
XFILL_5_DFFPOSX1_921 gnd vdd FILL
XFILL_5_DFFPOSX1_910 gnd vdd FILL
XFILL_5_DFFPOSX1_954 gnd vdd FILL
XFILL_5_DFFPOSX1_943 gnd vdd FILL
XFILL_5_DFFPOSX1_932 gnd vdd FILL
XFILL_5_DFFPOSX1_965 gnd vdd FILL
XAOI21X1_26 bundleStartMajId_i[2] AND2X2_17/Y bundleStartMajId_i[1] gnd AOI21X1_26/Y
+ vdd AOI21X1
XFILL_5_DFFPOSX1_998 gnd vdd FILL
XAOI21X1_15 bundleStartMajId_i[18] INVX2_50/A bundleStartMajId_i[17] gnd AOI21X1_15/Y
+ vdd AOI21X1
XFILL_5_DFFPOSX1_987 gnd vdd FILL
XFILL_5_DFFPOSX1_976 gnd vdd FILL
XAOI21X1_37 bundleAddress_i[33] NOR2X1_146/B INVX4_39/Y gnd AOI21X1_37/Y vdd AOI21X1
XAOI21X1_48 bundleAddress_i[34] NOR2X1_195/B bundleAddress_i[33] gnd AOI21X1_48/Y
+ vdd AOI21X1
XAOI21X1_59 bundleAddress_i[2] INVX1_217/Y bundleAddress_i[1] gnd AOI21X1_59/Y vdd
+ AOI21X1
XFILL_0_AND2X2_1 gnd vdd FILL
XFILL_4_DFFPOSX1_500 gnd vdd FILL
XFILL_4_DFFPOSX1_522 gnd vdd FILL
XFILL_4_DFFPOSX1_511 gnd vdd FILL
XFILL_4_DFFPOSX1_544 gnd vdd FILL
XFILL_4_DFFPOSX1_555 gnd vdd FILL
XFILL_4_DFFPOSX1_533 gnd vdd FILL
XFILL_4_DFFPOSX1_588 gnd vdd FILL
XFILL_4_DFFPOSX1_566 gnd vdd FILL
XFILL_4_DFFPOSX1_577 gnd vdd FILL
XFILL_27_9_0 gnd vdd FILL
XFILL_4_DFFPOSX1_599 gnd vdd FILL
XFILL_2_9_0 gnd vdd FILL
XFILL_1_BUFX2_1024 gnd vdd FILL
XFILL_1_BUFX2_401 gnd vdd FILL
XFILL_1_BUFX2_445 gnd vdd FILL
XFILL_1_BUFX2_434 gnd vdd FILL
XFILL_3_DFFPOSX1_112 gnd vdd FILL
XFILL_10_8_0 gnd vdd FILL
XFILL_1_BUFX2_478 gnd vdd FILL
XFILL_3_DFFPOSX1_101 gnd vdd FILL
XOAI21X1_440 NAND3X1_2/Y INVX4_12/Y BUFX4_245/Y gnd OAI21X1_441/A vdd OAI21X1
XFILL_3_DFFPOSX1_134 gnd vdd FILL
XFILL_1_BUFX2_489 gnd vdd FILL
XFILL_3_DFFPOSX1_145 gnd vdd FILL
XFILL_1_CLKBUF1_25 gnd vdd FILL
XFILL_1_CLKBUF1_14 gnd vdd FILL
XFILL_3_DFFPOSX1_123 gnd vdd FILL
XFILL_1_CLKBUF1_47 gnd vdd FILL
XFILL_23_15_1 gnd vdd FILL
XFILL_1_CLKBUF1_36 gnd vdd FILL
XOAI21X1_473 OAI21X1_473/A NOR2X1_43/Y OAI21X1_473/C gnd OAI21X1_473/Y vdd OAI21X1
XOAI21X1_462 OAI21X1_462/A INVX2_28/Y BUFX4_241/Y gnd OAI21X1_463/A vdd OAI21X1
XOAI21X1_484 INVX1_20/A INVX1_21/A BUFX4_244/Y gnd OAI21X1_485/B vdd OAI21X1
XOAI21X1_451 NOR2X1_26/Y bundleStartMajId_i[29] BUFX4_245/Y gnd OAI21X1_452/A vdd
+ OAI21X1
XFILL_3_DFFPOSX1_178 gnd vdd FILL
XFILL_3_DFFPOSX1_156 gnd vdd FILL
XOAI21X1_495 OAI21X1_499/A INVX4_27/Y BUFX4_240/Y gnd OAI21X1_496/A vdd OAI21X1
XFILL_1_CLKBUF1_69 gnd vdd FILL
XFILL_1_CLKBUF1_58 gnd vdd FILL
XFILL_3_DFFPOSX1_167 gnd vdd FILL
XFILL_3_DFFPOSX1_189 gnd vdd FILL
XFILL_6_DFFPOSX1_627 gnd vdd FILL
XFILL_6_DFFPOSX1_605 gnd vdd FILL
XFILL_6_DFFPOSX1_616 gnd vdd FILL
XNAND2X1_490 NAND2X1_490/A NAND2X1_492/B gnd NAND2X1_490/Y vdd NAND2X1
XFILL_2_OAI21X1_194 gnd vdd FILL
XFILL_0_INVX1_200 gnd vdd FILL
XFILL_0_INVX1_211 gnd vdd FILL
XFILL_18_9_0 gnd vdd FILL
XFILL_0_NAND2X1_219 gnd vdd FILL
XFILL_0_INVX1_222 gnd vdd FILL
XFILL_0_NAND2X1_208 gnd vdd FILL
XFILL_5_DFFPOSX1_217 gnd vdd FILL
XFILL_28_14_1 gnd vdd FILL
XFILL_5_DFFPOSX1_206 gnd vdd FILL
XFILL_5_DFFPOSX1_239 gnd vdd FILL
XFILL_5_DFFPOSX1_228 gnd vdd FILL
XFILL_0_OAI21X1_32 gnd vdd FILL
XFILL_0_OAI21X1_10 gnd vdd FILL
XFILL_0_OAI21X1_21 gnd vdd FILL
XOAI21X1_1714 BUFX4_137/Y BUFX4_60/A BUFX2_757/A gnd OAI21X1_1715/C vdd OAI21X1
XFILL_0_OAI21X1_65 gnd vdd FILL
XOAI21X1_1703 BUFX4_179/Y INVX2_145/Y OAI21X1_1703/C gnd DFFPOSX1_64/D vdd OAI21X1
XFILL_22_10_0 gnd vdd FILL
XFILL_0_OAI21X1_43 gnd vdd FILL
XFILL_0_OAI21X1_54 gnd vdd FILL
XFILL_1_BUFX2_990 gnd vdd FILL
XOAI21X1_1725 INVX2_124/Y BUFX4_292/Y OAI21X1_1725/C gnd DFFPOSX1_75/D vdd OAI21X1
XOAI21X1_1736 BUFX4_138/Y BUFX4_40/Y BUFX2_750/A gnd OAI21X1_1737/C vdd OAI21X1
XOAI21X1_1747 INVX2_135/Y BUFX4_296/Y OAI21X1_1747/C gnd DFFPOSX1_86/D vdd OAI21X1
XFILL_0_OAI21X1_87 gnd vdd FILL
XFILL_0_OAI21X1_98 gnd vdd FILL
XFILL_0_OAI21X1_76 gnd vdd FILL
XFILL_3_DFFPOSX1_690 gnd vdd FILL
XOAI21X1_1758 BUFX4_138/Y BUFX4_55/Y BUFX2_762/A gnd OAI21X1_1759/C vdd OAI21X1
XFILL_0_OAI21X1_714 gnd vdd FILL
XFILL_0_OAI21X1_703 gnd vdd FILL
XOAI21X1_1769 INVX2_114/Y BUFX4_297/Y OAI21X1_1769/C gnd DFFPOSX1_97/D vdd OAI21X1
XFILL_1_OAI21X1_907 gnd vdd FILL
XFILL_0_OAI21X1_747 gnd vdd FILL
XFILL_0_OAI21X1_736 gnd vdd FILL
XFILL_0_OAI21X1_725 gnd vdd FILL
XFILL_1_OAI21X1_918 gnd vdd FILL
XFILL_1_OAI21X1_929 gnd vdd FILL
XFILL_0_OAI21X1_758 gnd vdd FILL
XFILL_0_OAI21X1_769 gnd vdd FILL
XFILL_2_NAND3X1_19 gnd vdd FILL
XFILL_3_15_1 gnd vdd FILL
XFILL_0_NAND2X1_720 gnd vdd FILL
XFILL_0_NAND2X1_742 gnd vdd FILL
XFILL_0_NAND2X1_753 gnd vdd FILL
XFILL_0_NAND2X1_731 gnd vdd FILL
XFILL_0_OAI21X1_1524 gnd vdd FILL
XFILL_0_OAI21X1_1513 gnd vdd FILL
XFILL_0_OAI21X1_1502 gnd vdd FILL
XFILL_0_NAND2X1_764 gnd vdd FILL
XFILL_2_DFFPOSX1_291 gnd vdd FILL
XFILL_4_NOR3X1_1 gnd vdd FILL
XFILL_0_OAI21X1_1557 gnd vdd FILL
XFILL_0_OAI21X1_1546 gnd vdd FILL
XFILL_0_OAI21X1_1535 gnd vdd FILL
XFILL_2_DFFPOSX1_280 gnd vdd FILL
XFILL_5_DFFPOSX1_91 gnd vdd FILL
XFILL_0_OAI21X1_1568 gnd vdd FILL
XFILL_5_DFFPOSX1_80 gnd vdd FILL
XFILL_0_OAI21X1_1579 gnd vdd FILL
XFILL_5_DFFPOSX1_740 gnd vdd FILL
XFILL_5_DFFPOSX1_751 gnd vdd FILL
XFILL_5_DFFPOSX1_773 gnd vdd FILL
XFILL_5_DFFPOSX1_762 gnd vdd FILL
XFILL_5_DFFPOSX1_784 gnd vdd FILL
XFILL_5_DFFPOSX1_795 gnd vdd FILL
XFILL_8_14_1 gnd vdd FILL
XFILL_4_DFFPOSX1_330 gnd vdd FILL
XBUFX4_109 BUFX4_95/A gnd BUFX4_109/Y vdd BUFX4
XFILL_2_OAI21X1_1607 gnd vdd FILL
XFILL_4_DFFPOSX1_341 gnd vdd FILL
XFILL_4_DFFPOSX1_352 gnd vdd FILL
XFILL_5_0_1 gnd vdd FILL
XFILL_4_DFFPOSX1_363 gnd vdd FILL
XFILL_2_DFFPOSX1_1011 gnd vdd FILL
XFILL_2_DFFPOSX1_1000 gnd vdd FILL
XFILL_4_DFFPOSX1_374 gnd vdd FILL
XFILL_2_DFFPOSX1_1022 gnd vdd FILL
XFILL_4_DFFPOSX1_396 gnd vdd FILL
XFILL_4_DFFPOSX1_385 gnd vdd FILL
XFILL_2_10_0 gnd vdd FILL
XFILL_1_BUFX2_253 gnd vdd FILL
XFILL_1_BUFX2_231 gnd vdd FILL
XFILL_1_BUFX2_242 gnd vdd FILL
XFILL_1_BUFX2_286 gnd vdd FILL
XFILL_1_BUFX2_275 gnd vdd FILL
XFILL_1_OAI21X1_1208 gnd vdd FILL
XFILL_1_OAI21X1_1219 gnd vdd FILL
XOAI21X1_270 BUFX4_145/Y BUFX4_62/Y BUFX2_998/A gnd OAI21X1_271/C vdd OAI21X1
XFILL_1_BUFX2_297 gnd vdd FILL
XOAI21X1_292 BUFX4_134/Y BUFX4_76/Y BUFX2_1010/A gnd OAI21X1_293/C vdd OAI21X1
XOAI21X1_281 INVX2_186/Y INVX8_2/A OAI21X1_281/C gnd OAI21X1_281/Y vdd OAI21X1
XFILL_1_DFFPOSX1_809 gnd vdd FILL
XFILL_6_DFFPOSX1_468 gnd vdd FILL
XFILL_6_DFFPOSX1_479 gnd vdd FILL
XFILL_1_NAND3X1_5 gnd vdd FILL
XFILL_1_NAND2X1_209 gnd vdd FILL
XFILL_36_3 gnd vdd FILL
XFILL_33_7_0 gnd vdd FILL
XFILL_29_2 gnd vdd FILL
XFILL_5_DFFPOSX1_1004 gnd vdd FILL
XFILL_5_DFFPOSX1_1015 gnd vdd FILL
XFILL_5_DFFPOSX1_1026 gnd vdd FILL
XFILL_0_BUFX4_361 gnd vdd FILL
XDFFPOSX1_26 BUFX2_696/A CLKBUF1_16/Y DFFPOSX1_26/D gnd vdd DFFPOSX1
XDFFPOSX1_15 BUFX2_684/A CLKBUF1_61/Y DFFPOSX1_15/D gnd vdd DFFPOSX1
XOAI21X1_1522 NOR2X1_226/B INVX2_111/Y INVX1_178/Y gnd NAND2X1_641/A vdd OAI21X1
XOAI21X1_1511 BUFX4_160/Y OAI21X1_1511/B BUFX2_230/A gnd OAI21X1_1512/C vdd OAI21X1
XOAI21X1_1500 BUFX4_169/Y BUFX4_71/Y BUFX2_226/A gnd OAI21X1_1501/C vdd OAI21X1
XFILL_0_BUFX4_350 gnd vdd FILL
XDFFPOSX1_59 BUFX2_729/A CLKBUF1_32/Y DFFPOSX1_59/D gnd vdd DFFPOSX1
XDFFPOSX1_37 BUFX2_714/A CLKBUF1_65/Y DFFPOSX1_37/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1742 gnd vdd FILL
XFILL_1_OAI21X1_1731 gnd vdd FILL
XOAI21X1_1533 NAND2X1_642/Y BUFX4_301/Y OAI21X1_1533/C gnd OAI21X1_1533/Y vdd OAI21X1
XDFFPOSX1_48 BUFX2_717/A CLKBUF1_87/Y DFFPOSX1_48/D gnd vdd DFFPOSX1
XOAI21X1_1566 AOI21X1_65/Y OAI21X1_1566/B OAI21X1_1566/C gnd OAI21X1_1566/Y vdd OAI21X1
XFILL_0_BUFX4_372 gnd vdd FILL
XOAI21X1_1544 INVX4_48/Y OR2X2_21/A OAI21X1_1544/C gnd OAI21X1_1546/A vdd OAI21X1
XOAI21X1_1555 AOI21X1_64/Y OAI21X1_1555/B OAI21X1_1555/C gnd OAI21X1_1555/Y vdd OAI21X1
XFILL_1_OAI21X1_1720 gnd vdd FILL
XFILL_0_BUFX4_383 gnd vdd FILL
XOAI21X1_1588 BUFX4_336/Y INVX2_124/Y NAND2X1_657/Y gnd OAI21X1_1588/Y vdd OAI21X1
XFILL_1_OAI21X1_1764 gnd vdd FILL
XFILL_1_OAI21X1_1753 gnd vdd FILL
XOAI21X1_1599 BUFX4_376/Y INVX2_135/Y NAND2X1_668/Y gnd OAI21X1_1599/Y vdd OAI21X1
XOAI21X1_1577 BUFX4_95/Y BUFX4_324/Y BUFX2_391/A gnd OAI21X1_1578/C vdd OAI21X1
XFILL_0_OAI21X1_500 gnd vdd FILL
XFILL_0_BUFX2_1010 gnd vdd FILL
XFILL_1_OAI21X1_1775 gnd vdd FILL
XFILL_0_OAI21X1_511 gnd vdd FILL
XFILL_0_OAI21X1_522 gnd vdd FILL
XFILL_0_BUFX2_1021 gnd vdd FILL
XFILL_1_OAI21X1_1786 gnd vdd FILL
XFILL_0_BUFX2_1032 gnd vdd FILL
XFILL_1_OAI21X1_1797 gnd vdd FILL
XFILL_1_OAI21X1_715 gnd vdd FILL
XFILL_0_OAI21X1_555 gnd vdd FILL
XFILL_0_OAI21X1_533 gnd vdd FILL
XFILL_0_OAI21X1_544 gnd vdd FILL
XFILL_1_OAI21X1_704 gnd vdd FILL
XFILL_1_OAI21X1_726 gnd vdd FILL
XFILL_1_OAI21X1_737 gnd vdd FILL
XFILL_1_OAI21X1_759 gnd vdd FILL
XFILL_0_OAI21X1_566 gnd vdd FILL
XFILL_0_OAI21X1_577 gnd vdd FILL
XFILL_1_OAI21X1_748 gnd vdd FILL
XFILL_0_OAI21X1_599 gnd vdd FILL
XFILL_0_OAI21X1_588 gnd vdd FILL
XFILL_6_DFFPOSX1_980 gnd vdd FILL
XFILL_6_DFFPOSX1_991 gnd vdd FILL
XFILL_0_CLKBUF1_11 gnd vdd FILL
XFILL_0_CLKBUF1_22 gnd vdd FILL
XFILL_13_15_0 gnd vdd FILL
XFILL_0_CLKBUF1_44 gnd vdd FILL
XFILL_0_CLKBUF1_33 gnd vdd FILL
XFILL_0_CLKBUF1_55 gnd vdd FILL
XFILL_0_CLKBUF1_88 gnd vdd FILL
XFILL_0_CLKBUF1_77 gnd vdd FILL
XFILL_0_CLKBUF1_66 gnd vdd FILL
XFILL_1_NAND2X1_710 gnd vdd FILL
XFILL_0_CLKBUF1_99 gnd vdd FILL
XFILL_0_NAND2X1_561 gnd vdd FILL
XFILL_0_DFFPOSX1_900 gnd vdd FILL
XFILL_1_NAND2X1_721 gnd vdd FILL
XFILL_0_NAND2X1_550 gnd vdd FILL
XFILL_0_OAI21X1_1332 gnd vdd FILL
XFILL_0_OAI21X1_1310 gnd vdd FILL
XFILL_0_OAI21X1_1321 gnd vdd FILL
XFILL_1_NAND2X1_743 gnd vdd FILL
XFILL_0_NAND2X1_594 gnd vdd FILL
XFILL_1_NAND2X1_754 gnd vdd FILL
XFILL_24_7_0 gnd vdd FILL
XFILL_0_OAI21X1_1343 gnd vdd FILL
XFILL_0_NAND2X1_583 gnd vdd FILL
XFILL_0_DFFPOSX1_922 gnd vdd FILL
XFILL_0_DFFPOSX1_933 gnd vdd FILL
XFILL_0_OAI21X1_1376 gnd vdd FILL
XFILL_0_OAI21X1_1354 gnd vdd FILL
XFILL_0_OAI21X1_1365 gnd vdd FILL
XFILL_0_NAND2X1_572 gnd vdd FILL
XFILL_0_DFFPOSX1_911 gnd vdd FILL
XFILL_0_OAI21X1_1398 gnd vdd FILL
XFILL_6_DFFPOSX1_70 gnd vdd FILL
XFILL_0_DFFPOSX1_944 gnd vdd FILL
XFILL_0_DFFPOSX1_966 gnd vdd FILL
XFILL_0_OAI21X1_1387 gnd vdd FILL
XFILL_0_DFFPOSX1_955 gnd vdd FILL
XFILL_0_DFFPOSX1_977 gnd vdd FILL
XFILL_6_DFFPOSX1_81 gnd vdd FILL
XFILL_0_DFFPOSX1_999 gnd vdd FILL
XFILL_0_DFFPOSX1_988 gnd vdd FILL
XFILL_0_OR2X2_5 gnd vdd FILL
XFILL_5_DFFPOSX1_570 gnd vdd FILL
XFILL_5_DFFPOSX1_581 gnd vdd FILL
XINVX2_109 INVX2_109/A gnd INVX2_109/Y vdd INVX2
XFILL_5_DFFPOSX1_592 gnd vdd FILL
XFILL_0_BUFX2_309 gnd vdd FILL
XFILL_1_BUFX4_3 gnd vdd FILL
XFILL_18_14_0 gnd vdd FILL
XFILL_7_8_0 gnd vdd FILL
XFILL_31_16_0 gnd vdd FILL
XFILL_2_OAI21X1_1437 gnd vdd FILL
XFILL_4_DFFPOSX1_171 gnd vdd FILL
XCLKBUF1_90 BUFX4_90/Y gnd CLKBUF1_90/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_160 gnd vdd FILL
XFILL_4_DFFPOSX1_182 gnd vdd FILL
XFILL_2_NOR3X1_15 gnd vdd FILL
XFILL_4_DFFPOSX1_193 gnd vdd FILL
XFILL_15_7_0 gnd vdd FILL
XFILL_0_INVX1_7 gnd vdd FILL
XFILL_1_NAND3X1_16 gnd vdd FILL
XFILL_1_NAND3X1_27 gnd vdd FILL
XFILL_1_OAI21X1_1005 gnd vdd FILL
XFILL_1_OAI21X1_1038 gnd vdd FILL
XFILL_0_BUFX2_821 gnd vdd FILL
XFILL_1_NAND3X1_38 gnd vdd FILL
XFILL_1_DFFPOSX1_606 gnd vdd FILL
XFILL_0_BUFX2_810 gnd vdd FILL
XDFFPOSX1_408 BUFX2_441/A CLKBUF1_80/Y OAI21X1_380/Y gnd vdd DFFPOSX1
XFILL_1_NAND3X1_49 gnd vdd FILL
XDFFPOSX1_419 BUFX2_453/A CLKBUF1_44/Y OAI21X1_391/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1016 gnd vdd FILL
XFILL_0_BUFX2_832 gnd vdd FILL
XFILL_0_BUFX2_843 gnd vdd FILL
XFILL_1_OAI21X1_1027 gnd vdd FILL
XINVX1_120 bundle_i[84] gnd INVX1_120/Y vdd INVX1
XINVX1_142 bundle_i[126] gnd INVX1_142/Y vdd INVX1
XFILL_0_BUFX2_865 gnd vdd FILL
XFILL_1_DFFPOSX1_639 gnd vdd FILL
XFILL_1_OAI21X1_1049 gnd vdd FILL
XINVX1_131 bundle_i[73] gnd INVX1_131/Y vdd INVX1
XFILL_1_DFFPOSX1_617 gnd vdd FILL
XFILL_1_DFFPOSX1_628 gnd vdd FILL
XFILL_0_BUFX2_876 gnd vdd FILL
XFILL_0_BUFX2_854 gnd vdd FILL
XFILL_0_BUFX2_887 gnd vdd FILL
XINVX1_186 INVX1_186/A gnd INVX1_186/Y vdd INVX1
XINVX1_164 bundle_i[104] gnd INVX1_164/Y vdd INVX1
XINVX1_175 bundleAddress_i[39] gnd INVX1_175/Y vdd INVX1
XFILL_0_BUFX2_898 gnd vdd FILL
XINVX1_153 bundle_i[115] gnd INVX1_153/Y vdd INVX1
XFILL_6_DFFPOSX1_232 gnd vdd FILL
XFILL_6_DFFPOSX1_243 gnd vdd FILL
XFILL_6_DFFPOSX1_221 gnd vdd FILL
XINVX1_197 INVX1_197/A gnd INVX1_197/Y vdd INVX1
XFILL_36_15_0 gnd vdd FILL
XFILL_6_DFFPOSX1_254 gnd vdd FILL
XFILL_6_DFFPOSX1_276 gnd vdd FILL
XFILL_6_DFFPOSX1_265 gnd vdd FILL
XCLKBUF1_101 BUFX4_85/Y gnd CLKBUF1_101/Y vdd CLKBUF1
XFILL_0_INVX2_30 gnd vdd FILL
XFILL_0_INVX2_63 gnd vdd FILL
XFILL_0_INVX2_41 gnd vdd FILL
XFILL_0_INVX2_52 gnd vdd FILL
XFILL_0_INVX2_96 gnd vdd FILL
XFILL_0_INVX2_74 gnd vdd FILL
XFILL_0_INVX2_85 gnd vdd FILL
XFILL_1_NOR3X1_5 gnd vdd FILL
XFILL_0_DFFPOSX1_218 gnd vdd FILL
XFILL_0_DFFPOSX1_207 gnd vdd FILL
XFILL_0_DFFPOSX1_229 gnd vdd FILL
XOAI21X1_1341 AOI21X1_53/Y OAI21X1_1341/B OAI21X1_1341/C gnd OAI21X1_1341/Y vdd OAI21X1
XOAI21X1_1330 OAI21X1_1330/A AOI21X1_51/Y OAI21X1_1330/C gnd OAI21X1_1330/Y vdd OAI21X1
XFILL_0_BUFX4_191 gnd vdd FILL
XDFFPOSX1_942 BUFX2_249/A CLKBUF1_98/Y OAI21X1_1401/Y gnd vdd DFFPOSX1
XDFFPOSX1_920 BUFX2_172/A CLKBUF1_21/Y OAI21X1_1341/Y gnd vdd DFFPOSX1
XOAI21X1_1374 BUFX4_111/Y BUFX4_348/Y BUFX2_186/A gnd OAI21X1_1375/C vdd OAI21X1
XFILL_0_BUFX4_180 gnd vdd FILL
XDFFPOSX1_931 BUFX2_184/A CLKBUF1_40/Y OAI21X1_1373/Y gnd vdd DFFPOSX1
XOAI21X1_1352 OAI21X1_1352/A AOI21X1_55/Y OAI21X1_1352/C gnd OAI21X1_1352/Y vdd OAI21X1
XFILL_1_OAI21X1_1550 gnd vdd FILL
XOAI21X1_1363 INVX2_104/Y INVX1_215/A OAI21X1_1363/C gnd OAI21X1_1364/A vdd OAI21X1
XFILL_1_OAI21X1_1594 gnd vdd FILL
XFILL_1_BUFX2_91 gnd vdd FILL
XOAI21X1_1385 INVX2_54/Y BUFX4_301/Y OAI21X1_1385/C gnd OAI21X1_1385/Y vdd OAI21X1
XFILL_1_OAI21X1_1583 gnd vdd FILL
XOAI21X1_1396 NOR2X1_215/B INVX2_57/Y INVX2_58/Y gnd OAI21X1_1397/C vdd OAI21X1
XDFFPOSX1_953 BUFX2_202/A CLKBUF1_23/Y OAI21X1_1435/Y gnd vdd DFFPOSX1
XDFFPOSX1_964 BUFX2_214/A CLKBUF1_27/Y OAI21X1_1466/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1572 gnd vdd FILL
XFILL_1_OAI21X1_501 gnd vdd FILL
XFILL_1_OAI21X1_1561 gnd vdd FILL
XFILL_0_OAI21X1_330 gnd vdd FILL
XFILL_1_BUFX2_80 gnd vdd FILL
XDFFPOSX1_975 BUFX2_226/A CLKBUF1_34/Y OAI21X1_1501/Y gnd vdd DFFPOSX1
XFILL_1_NOR2X1_117 gnd vdd FILL
XDFFPOSX1_997 BUFX2_251/A CLKBUF1_36/Y OAI21X1_1569/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_534 gnd vdd FILL
XFILL_0_OAI21X1_341 gnd vdd FILL
XFILL_1_OAI21X1_545 gnd vdd FILL
XDFFPOSX1_986 BUFX2_239/A CLKBUF1_81/Y OAI21X1_1535/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_352 gnd vdd FILL
XFILL_0_OAI21X1_363 gnd vdd FILL
XFILL_1_OAI21X1_523 gnd vdd FILL
XFILL_1_OAI21X1_512 gnd vdd FILL
XFILL_0_OAI21X1_385 gnd vdd FILL
XFILL_2_OAI21X1_738 gnd vdd FILL
XFILL_1_OAI21X1_567 gnd vdd FILL
XFILL_1_OAI21X1_556 gnd vdd FILL
XFILL_1_OAI21X1_578 gnd vdd FILL
XFILL_0_OAI21X1_396 gnd vdd FILL
XFILL_0_OAI21X1_374 gnd vdd FILL
XFILL_1_NOR2X1_139 gnd vdd FILL
XFILL_1_OAI21X1_589 gnd vdd FILL
XFILL_1_OAI21X1_2 gnd vdd FILL
XFILL_1_NAND2X1_551 gnd vdd FILL
XFILL_0_OAI21X1_1151 gnd vdd FILL
XFILL_1_BUFX4_304 gnd vdd FILL
XFILL_1_NAND2X1_540 gnd vdd FILL
XFILL_0_NAND2X1_380 gnd vdd FILL
XFILL_0_OAI21X1_1140 gnd vdd FILL
XFILL_0_DFFPOSX1_741 gnd vdd FILL
XFILL_0_DFFPOSX1_752 gnd vdd FILL
XFILL_0_OAI21X1_1173 gnd vdd FILL
XFILL_1_NAND2X1_584 gnd vdd FILL
XFILL_1_NAND2X1_562 gnd vdd FILL
XFILL_0_OAI21X1_1184 gnd vdd FILL
XFILL_1_NAND2X1_573 gnd vdd FILL
XFILL_0_NAND2X1_391 gnd vdd FILL
XFILL_1_BUFX4_326 gnd vdd FILL
XFILL_1_BUFX4_315 gnd vdd FILL
XFILL_1_BUFX4_337 gnd vdd FILL
XFILL_0_DFFPOSX1_730 gnd vdd FILL
XFILL_0_OAI21X1_1162 gnd vdd FILL
XFILL_0_DFFPOSX1_774 gnd vdd FILL
XFILL_1_BUFX4_359 gnd vdd FILL
XFILL_1_NAND2X1_595 gnd vdd FILL
XFILL_1_BUFX4_348 gnd vdd FILL
XFILL_0_DFFPOSX1_763 gnd vdd FILL
XFILL_0_OAI21X1_1195 gnd vdd FILL
XFILL_0_DFFPOSX1_785 gnd vdd FILL
XFILL_0_DFFPOSX1_796 gnd vdd FILL
XFILL_2_OAI21X1_28 gnd vdd FILL
XFILL_0_BUFX2_106 gnd vdd FILL
XFILL_0_BUFX2_128 gnd vdd FILL
XFILL_0_BUFX2_117 gnd vdd FILL
XFILL_0_BUFX2_139 gnd vdd FILL
XFILL_20_13_1 gnd vdd FILL
XINVX4_50 INVX4_50/A gnd INVX4_50/Y vdd INVX4
XFILL_1_NAND2X1_60 gnd vdd FILL
XFILL_1_NAND2X1_93 gnd vdd FILL
XFILL_1_NAND2X1_82 gnd vdd FILL
XBUFX2_911 BUFX2_911/A gnd tid3_o[49] vdd BUFX2
XBUFX2_922 BUFX2_922/A gnd tid3_o[39] vdd BUFX2
XFILL_2_DFFPOSX1_813 gnd vdd FILL
XFILL_2_DFFPOSX1_824 gnd vdd FILL
XFILL_2_DFFPOSX1_802 gnd vdd FILL
XBUFX2_900 BUFX2_900/A gnd tid2_o[1] vdd BUFX2
XBUFX2_944 BUFX2_944/A gnd tid3_o[19] vdd BUFX2
XBUFX2_933 BUFX2_933/A gnd tid3_o[29] vdd BUFX2
XBUFX2_955 BUFX2_955/A gnd tid3_o[9] vdd BUFX2
XFILL_2_DFFPOSX1_835 gnd vdd FILL
XFILL_2_OAI21X1_1289 gnd vdd FILL
XFILL_2_OAI21X1_1278 gnd vdd FILL
XFILL_2_DFFPOSX1_857 gnd vdd FILL
XFILL_2_DFFPOSX1_846 gnd vdd FILL
XBUFX2_988 BUFX2_988/A gnd tid4_o[37] vdd BUFX2
XFILL_2_DFFPOSX1_879 gnd vdd FILL
XBUFX2_977 BUFX2_977/A gnd tid4_o[47] vdd BUFX2
XBUFX2_966 BUFX2_966/A gnd tid3_o[56] vdd BUFX2
XFILL_2_DFFPOSX1_868 gnd vdd FILL
XBUFX2_999 BUFX2_999/A gnd tid4_o[27] vdd BUFX2
XFILL_30_5_0 gnd vdd FILL
XFILL_25_12_1 gnd vdd FILL
XFILL_1_DFFPOSX1_414 gnd vdd FILL
XFILL_0_BUFX2_651 gnd vdd FILL
XFILL_0_BUFX2_640 gnd vdd FILL
XFILL_1_DFFPOSX1_403 gnd vdd FILL
XFILL_2_AOI21X1_8 gnd vdd FILL
XDFFPOSX1_205 BUFX2_877/A CLKBUF1_38/Y OAI21X1_49/Y gnd vdd DFFPOSX1
XDFFPOSX1_216 BUFX2_889/A CLKBUF1_2/Y OAI21X1_60/Y gnd vdd DFFPOSX1
XDFFPOSX1_227 BUFX2_901/A CLKBUF1_58/Y OAI21X1_71/Y gnd vdd DFFPOSX1
XDFFPOSX1_249 BUFX2_919/A CLKBUF1_98/Y OAI21X1_115/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_662 gnd vdd FILL
XFILL_0_BUFX2_684 gnd vdd FILL
XDFFPOSX1_238 BUFX2_907/A CLKBUF1_35/Y OAI21X1_93/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_673 gnd vdd FILL
XFILL_1_DFFPOSX1_447 gnd vdd FILL
XFILL_1_DFFPOSX1_425 gnd vdd FILL
XFILL_1_DFFPOSX1_436 gnd vdd FILL
XFILL_0_BUFX2_695 gnd vdd FILL
XFILL_1_DFFPOSX1_458 gnd vdd FILL
XFILL_1_DFFPOSX1_469 gnd vdd FILL
XNAND2X1_308 INVX2_52/A NOR2X1_4/Y gnd NOR2X1_105/A vdd NAND2X1
XNAND2X1_319 NOR2X1_16/Y NOR2X1_105/Y gnd NOR2X1_108/B vdd NAND2X1
XFILL_4_DFFPOSX1_918 gnd vdd FILL
XFILL_4_DFFPOSX1_929 gnd vdd FILL
XFILL_4_DFFPOSX1_907 gnd vdd FILL
XFILL_38_6_0 gnd vdd FILL
XNOR3X1_15 INVX2_92/Y INVX4_49/Y NOR3X1_15/C gnd NOR3X1_15/Y vdd NOR3X1
XBUFX4_281 INVX8_7/Y gnd BUFX4_64/A vdd BUFX4
XBUFX4_270 INVX8_7/Y gnd BUFX4_51/A vdd BUFX4
XFILL_0_INVX2_180 gnd vdd FILL
XBUFX4_292 BUFX4_303/A gnd BUFX4_292/Y vdd BUFX4
XFILL_0_13_1 gnd vdd FILL
XFILL_0_INVX2_191 gnd vdd FILL
XFILL_0_XNOR2X1_7 gnd vdd FILL
XFILL_1_BUFX2_808 gnd vdd FILL
XFILL_1_BUFX2_819 gnd vdd FILL
XOAI21X1_803 INVX2_51/Y INVX2_53/Y OAI21X1_803/C gnd OAI21X1_805/A vdd OAI21X1
XFILL_21_5_0 gnd vdd FILL
XOAI21X1_814 BUFX4_142/Y BUFX4_41/Y BUFX2_634/A gnd OAI21X1_815/C vdd OAI21X1
XOAI21X1_858 INVX1_59/Y BUFX4_263/Y OAI21X1_858/C gnd OAI21X1_858/Y vdd OAI21X1
XOAI21X1_836 OAI21X1_839/A INVX4_27/Y BUFX4_288/Y gnd OAI21X1_837/B vdd OAI21X1
XOAI21X1_825 BUFX4_171/Y BUFX4_64/A BUFX2_638/A gnd OAI21X1_826/C vdd OAI21X1
XFILL_3_DFFPOSX1_519 gnd vdd FILL
XOAI21X1_847 INVX1_48/Y INVX8_4/A OAI21X1_847/C gnd OAI21X1_847/Y vdd OAI21X1
XFILL_3_DFFPOSX1_508 gnd vdd FILL
XOAI21X1_869 INVX1_70/Y BUFX4_264/Y OAI21X1_869/C gnd OAI21X1_869/Y vdd OAI21X1
XDFFPOSX1_750 BUFX2_57/A CLKBUF1_31/Y OAI21X1_1042/Y gnd vdd DFFPOSX1
XOAI21X1_1171 INVX1_194/A INVX4_43/Y INVX1_177/Y gnd NAND2X1_554/B vdd OAI21X1
XOAI21X1_1182 NOR3X1_14/C INVX4_44/Y INVX2_84/Y gnd NAND2X1_568/A vdd OAI21X1
XOAI21X1_1160 XNOR2X1_68/Y OAI21X1_9/B NAND2X1_537/Y gnd OAI21X1_1160/Y vdd OAI21X1
XDFFPOSX1_761 BUFX2_10/A CLKBUF1_102/Y OAI21X1_1053/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1391 gnd vdd FILL
XDFFPOSX1_772 BUFX2_22/A CLKBUF1_55/Y OAI21X1_1064/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1380 gnd vdd FILL
XFILL_1_DFFPOSX1_970 gnd vdd FILL
XFILL_1_OAI21X1_320 gnd vdd FILL
XOAI21X1_1193 OAI21X1_1193/A AOI21X1_42/Y NAND2X1_578/Y gnd OAI21X1_1193/Y vdd OAI21X1
XDFFPOSX1_783 BUFX2_34/A CLKBUF1_53/Y OAI21X1_1075/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_160 gnd vdd FILL
XFILL_1_DFFPOSX1_981 gnd vdd FILL
XFILL_1_OAI21X1_353 gnd vdd FILL
XFILL_0_OAI21X1_171 gnd vdd FILL
XFILL_0_OAI21X1_182 gnd vdd FILL
XFILL_1_OAI21X1_331 gnd vdd FILL
XFILL_1_DFFPOSX1_992 gnd vdd FILL
XFILL_1_OAI21X1_342 gnd vdd FILL
XDFFPOSX1_794 BUFX2_47/A CLKBUF1_76/Y OAI21X1_1086/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_386 gnd vdd FILL
XFILL_1_OAI21X1_364 gnd vdd FILL
XFILL_1_OAI21X1_375 gnd vdd FILL
XFILL_2_OAI21X1_546 gnd vdd FILL
XFILL_0_OAI21X1_193 gnd vdd FILL
XFILL_1_CLKBUF1_7 gnd vdd FILL
XFILL_1_OAI21X1_397 gnd vdd FILL
XFILL_5_12_1 gnd vdd FILL
XFILL_29_6_0 gnd vdd FILL
XFILL_0_NAND3X1_13 gnd vdd FILL
XFILL_2_DFFPOSX1_109 gnd vdd FILL
XFILL_0_NAND3X1_35 gnd vdd FILL
XFILL_0_NAND3X1_24 gnd vdd FILL
XBUFX2_207 BUFX2_207/A gnd addr4_o[42] vdd BUFX2
XFILL_4_6_0 gnd vdd FILL
XBUFX2_218 BUFX2_218/A gnd addr4_o[32] vdd BUFX2
XFILL_0_NAND3X1_46 gnd vdd FILL
XFILL_0_NAND3X1_57 gnd vdd FILL
XBUFX2_229 BUFX2_229/A gnd addr4_o[22] vdd BUFX2
XFILL_0_NAND3X1_68 gnd vdd FILL
XFILL_0_BUFX4_70 gnd vdd FILL
XFILL_0_BUFX4_81 gnd vdd FILL
XFILL_1_BUFX4_101 gnd vdd FILL
XFILL_0_BUFX4_92 gnd vdd FILL
XFILL_1_BUFX4_112 gnd vdd FILL
XFILL_1_NAND2X1_392 gnd vdd FILL
XFILL_1_BUFX4_123 gnd vdd FILL
XFILL_1_BUFX4_145 gnd vdd FILL
XFILL_0_DFFPOSX1_560 gnd vdd FILL
XFILL_1_BUFX4_134 gnd vdd FILL
XFILL_1_BUFX4_178 gnd vdd FILL
XFILL_1_BUFX4_156 gnd vdd FILL
XFILL_0_DFFPOSX1_582 gnd vdd FILL
XFILL_0_DFFPOSX1_593 gnd vdd FILL
XFILL_12_5_0 gnd vdd FILL
XFILL_1_BUFX4_167 gnd vdd FILL
XFILL_1_BUFX4_189 gnd vdd FILL
XFILL_0_DFFPOSX1_571 gnd vdd FILL
XFILL_2_CLKBUF1_29 gnd vdd FILL
XFILL_2_CLKBUF1_18 gnd vdd FILL
XBUFX2_730 BUFX2_730/A gnd pid3_o[7] vdd BUFX2
XFILL_2_OAI21X1_1042 gnd vdd FILL
XFILL_2_DFFPOSX1_632 gnd vdd FILL
XFILL_2_DFFPOSX1_621 gnd vdd FILL
XFILL_2_DFFPOSX1_610 gnd vdd FILL
XFILL_11_18_1 gnd vdd FILL
XFILL_2_DFFPOSX1_654 gnd vdd FILL
XBUFX2_752 BUFX2_752/A gnd pid4_o[16] vdd BUFX2
XBUFX2_763 BUFX2_763/A gnd pid4_o[6] vdd BUFX2
XNOR2X1_81 NOR2X1_81/A NOR2X1_89/B gnd NOR2X1_81/Y vdd NOR2X1
XNOR2X1_70 OR2X2_4/A NOR2X1_70/B gnd NOR2X1_71/B vdd NOR2X1
XFILL_2_DFFPOSX1_643 gnd vdd FILL
XFILL_2_DFFPOSX1_665 gnd vdd FILL
XBUFX2_741 BUFX2_741/A gnd pid3_o[25] vdd BUFX2
XBUFX2_796 BUFX2_796/A gnd tid1_o[37] vdd BUFX2
XBUFX2_774 BUFX2_774/A gnd pid4_o[24] vdd BUFX2
XFILL_2_DFFPOSX1_698 gnd vdd FILL
XFILL_3_DFFPOSX1_90 gnd vdd FILL
XBUFX2_785 BUFX2_785/A gnd tid1_o[47] vdd BUFX2
XNOR2X1_92 INVX4_23/Y NOR2X1_97/B gnd NOR2X1_93/B vdd NOR2X1
XFILL_2_DFFPOSX1_687 gnd vdd FILL
XFILL_2_DFFPOSX1_676 gnd vdd FILL
XFILL_0_NOR2X1_103 gnd vdd FILL
XFILL_0_NOR2X1_125 gnd vdd FILL
XFILL_0_NOR2X1_136 gnd vdd FILL
XFILL_0_NOR2X1_114 gnd vdd FILL
XFILL_0_NOR2X1_147 gnd vdd FILL
XFILL_0_NOR2X1_169 gnd vdd FILL
XFILL_0_NOR2X1_158 gnd vdd FILL
XBUFX2_8 BUFX2_8/A gnd addr1_o[48] vdd BUFX2
XFILL_1_DFFPOSX1_211 gnd vdd FILL
XFILL_1_DFFPOSX1_200 gnd vdd FILL
XFILL_1_DFFPOSX1_222 gnd vdd FILL
XFILL_1_DFFPOSX1_255 gnd vdd FILL
XFILL_0_BUFX2_481 gnd vdd FILL
XFILL_1_DFFPOSX1_244 gnd vdd FILL
XFILL_0_BUFX2_470 gnd vdd FILL
XFILL_0_BUFX2_492 gnd vdd FILL
XFILL_1_DFFPOSX1_233 gnd vdd FILL
XFILL_1_DFFPOSX1_266 gnd vdd FILL
XFILL_1_DFFPOSX1_299 gnd vdd FILL
XFILL_1_DFFPOSX1_277 gnd vdd FILL
XNAND2X1_116 BUFX2_432/A BUFX4_372/Y gnd OAI21X1_372/C vdd NAND2X1
XFILL_1_DFFPOSX1_288 gnd vdd FILL
XNAND2X1_105 BUFX2_420/A BUFX4_335/Y gnd OAI21X1_361/C vdd NAND2X1
XFILL_4_DFFPOSX1_704 gnd vdd FILL
XNAND2X1_138 BUFX4_244/Y NOR2X1_2/Y gnd OAI21X1_393/C vdd NAND2X1
XNAND2X1_127 BUFX2_444/A BUFX4_335/Y gnd OAI21X1_383/C vdd NAND2X1
XNAND2X1_149 bundleStartMajId_i[57] bundleStartMajId_i[56] gnd NOR2X1_4/B vdd NAND2X1
XFILL_4_DFFPOSX1_715 gnd vdd FILL
XFILL_1_OAI21X1_25 gnd vdd FILL
XFILL_4_DFFPOSX1_737 gnd vdd FILL
XFILL_1_OAI21X1_14 gnd vdd FILL
XFILL_16_17_1 gnd vdd FILL
XFILL_4_DFFPOSX1_726 gnd vdd FILL
XNAND2X1_3 NAND2X1_3/A OAI21X1_4/A gnd OAI21X1_3/C vdd NAND2X1
XFILL_1_OAI21X1_58 gnd vdd FILL
XFILL_4_DFFPOSX1_759 gnd vdd FILL
XFILL_4_DFFPOSX1_748 gnd vdd FILL
XFILL_1_OAI21X1_47 gnd vdd FILL
XFILL_1_OAI21X1_36 gnd vdd FILL
XFILL_1_OAI21X1_69 gnd vdd FILL
XFILL_10_13_0 gnd vdd FILL
XFILL_0_NAND2X1_90 gnd vdd FILL
XNOR2X1_160 INVX1_224/A NOR2X1_160/B gnd NOR2X1_160/Y vdd NOR2X1
XNOR2X1_182 INVX2_67/Y INVX4_34/Y gnd INVX2_105/A vdd NOR2X1
XNOR2X1_193 OR2X2_19/Y NOR2X1_193/B gnd NOR2X1_193/Y vdd NOR2X1
XNOR2X1_171 INVX4_45/Y INVX2_88/Y gnd INVX2_104/A vdd NOR2X1
XFILL_1_BUFX2_616 gnd vdd FILL
XFILL_1_BUFX2_627 gnd vdd FILL
XOAI21X1_633 AOI21X1_19/Y OAI21X1_633/B OAI21X1_633/C gnd OAI21X1_633/Y vdd OAI21X1
XOAI21X1_611 NOR2X1_85/Y OAI21X1_611/B OAI21X1_611/C gnd OAI21X1_611/Y vdd OAI21X1
XOAI21X1_600 OAI21X1_600/A BUFX4_155/Y OAI21X1_600/C gnd OAI21X1_600/Y vdd OAI21X1
XOAI21X1_622 INVX2_50/Y NOR3X1_3/C NOR2X1_89/B gnd OAI21X1_623/A vdd OAI21X1
XINVX2_8 bundleStartMajId_i[62] gnd INVX2_8/Y vdd INVX2
XFILL_3_DFFPOSX1_316 gnd vdd FILL
XOAI21X1_655 BUFX4_94/A BUFX4_340/Y BUFX2_580/A gnd OAI21X1_657/C vdd OAI21X1
XOAI21X1_644 BUFX4_251/Y BUFX4_328/Y BUFX2_575/A gnd OAI21X1_646/C vdd OAI21X1
XFILL_3_DFFPOSX1_327 gnd vdd FILL
XAOI21X1_8 bundleStartMajId_i[31] OR2X2_7/A BUFX4_175/Y gnd AOI21X1_9/A vdd AOI21X1
XOAI21X1_666 NOR2X1_2/A INVX2_9/Y INVX2_10/Y gnd OAI21X1_667/C vdd OAI21X1
XFILL_3_DFFPOSX1_305 gnd vdd FILL
XFILL_3_DFFPOSX1_349 gnd vdd FILL
XFILL_3_DFFPOSX1_338 gnd vdd FILL
XOAI21X1_699 BUFX4_167/Y BUFX4_69/Y BUFX2_591/A gnd OAI21X1_700/C vdd OAI21X1
XOAI21X1_688 AOI21X1_30/Y OAI21X1_688/B OAI21X1_688/C gnd OAI21X1_688/Y vdd OAI21X1
XOAI21X1_677 BUFX4_163/Y BUFX4_42/Y BUFX2_641/A gnd OAI21X1_678/C vdd OAI21X1
XFILL_6_DFFPOSX1_809 gnd vdd FILL
XDFFPOSX1_591 BUFX2_623/A CLKBUF1_100/Y OAI21X1_782/Y gnd vdd DFFPOSX1
XDFFPOSX1_580 BUFX2_611/A CLKBUF1_9/Y OAI21X1_750/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_161 gnd vdd FILL
XXNOR2X1_38 NOR2X1_94/Y bundleStartMajId_i[12] gnd XNOR2X1_38/Y vdd XNOR2X1
XXNOR2X1_16 NOR2X1_32/Y bundleStartMajId_i[26] gnd XNOR2X1_16/Y vdd XNOR2X1
XFILL_1_OAI21X1_150 gnd vdd FILL
XXNOR2X1_27 XNOR2X1_27/A INVX4_6/Y gnd XNOR2X1_27/Y vdd XNOR2X1
XFILL_1_OAI21X1_172 gnd vdd FILL
XFILL_34_18_1 gnd vdd FILL
XNAND2X1_650 BUFX2_649/A BUFX4_313/Y gnd NAND2X1_650/Y vdd NAND2X1
XNAND2X1_672 BUFX2_664/A OAI21X1_1/A gnd NAND2X1_672/Y vdd NAND2X1
XNAND2X1_661 BUFX2_652/A BUFX4_366/Y gnd NAND2X1_661/Y vdd NAND2X1
XFILL_1_OAI21X1_194 gnd vdd FILL
XXNOR2X1_49 INVX1_41/A OR2X2_8/B gnd XNOR2X1_49/Y vdd XNOR2X1
XFILL_1_OAI21X1_183 gnd vdd FILL
XINVX1_40 NOR3X1_7/C gnd INVX1_40/Y vdd INVX1
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XNAND2X1_683 BUFX2_682/A BUFX4_235/Y gnd NAND2X1_683/Y vdd NAND2X1
XINVX1_84 bundle_i[56] gnd INVX1_84/Y vdd INVX1
XINVX1_62 INVX1_62/A gnd INVX1_62/Y vdd INVX1
XNAND2X1_694 BUFX2_685/A BUFX4_183/Y gnd NAND2X1_694/Y vdd NAND2X1
XFILL_15_12_0 gnd vdd FILL
XFILL_2_OAI21X1_398 gnd vdd FILL
XINVX1_73 INVX1_73/A gnd INVX1_73/Y vdd INVX1
XBUFX2_26 BUFX2_26/A gnd addr1_o[32] vdd BUFX2
XINVX1_95 bundle_i[45] gnd INVX1_95/Y vdd INVX1
XBUFX2_15 BUFX2_15/A gnd addr1_o[42] vdd BUFX2
XBUFX2_59 BUFX2_59/A gnd addr1_o[2] vdd BUFX2
XBUFX2_37 BUFX2_37/A gnd addr1_o[22] vdd BUFX2
XDFFPOSX1_3 BUFX2_674/A CLKBUF1_66/Y DFFPOSX1_3/D gnd vdd DFFPOSX1
XBUFX2_48 BUFX2_48/A gnd addr1_o[12] vdd BUFX2
XFILL_1_BUFX4_26 gnd vdd FILL
XFILL_1_BUFX4_15 gnd vdd FILL
XFILL_0_DFFPOSX1_390 gnd vdd FILL
XFILL_1_BUFX4_48 gnd vdd FILL
XFILL_1_BUFX4_59 gnd vdd FILL
XFILL_1_BUFX4_37 gnd vdd FILL
XFILL_3_DFFPOSX1_850 gnd vdd FILL
XFILL_3_DFFPOSX1_883 gnd vdd FILL
XFILL_3_DFFPOSX1_872 gnd vdd FILL
XFILL_3_DFFPOSX1_861 gnd vdd FILL
XFILL_0_OAI21X1_907 gnd vdd FILL
XFILL_0_OAI21X1_929 gnd vdd FILL
XFILL_3_DFFPOSX1_894 gnd vdd FILL
XNOR2X1_6 OR2X2_1/Y NOR2X1_6/B gnd NOR2X1_6/Y vdd NOR2X1
XFILL_0_OAI21X1_918 gnd vdd FILL
XFILL_33_13_0 gnd vdd FILL
XFILL_36_9_1 gnd vdd FILL
XFILL_35_4_0 gnd vdd FILL
XFILL_1_OR2X2_18 gnd vdd FILL
XFILL_0_OAI21X1_1706 gnd vdd FILL
XFILL_2_DFFPOSX1_440 gnd vdd FILL
XFILL_0_OAI21X1_1739 gnd vdd FILL
XFILL_0_OAI21X1_1728 gnd vdd FILL
XFILL_0_OAI21X1_1717 gnd vdd FILL
XFILL_2_DFFPOSX1_462 gnd vdd FILL
XBUFX2_560 BUFX2_560/A gnd majID3_o[19] vdd BUFX2
XFILL_2_DFFPOSX1_451 gnd vdd FILL
XFILL_2_DFFPOSX1_473 gnd vdd FILL
XBUFX2_571 BUFX2_571/A gnd majID3_o[9] vdd BUFX2
XFILL_4_DFFPOSX1_91 gnd vdd FILL
XFILL_4_DFFPOSX1_80 gnd vdd FILL
XFILL_2_DFFPOSX1_484 gnd vdd FILL
XFILL_2_DFFPOSX1_495 gnd vdd FILL
XBUFX2_582 BUFX2_582/A gnd majID3_o[56] vdd BUFX2
XBUFX2_593 BUFX2_593/A gnd majID4_o[47] vdd BUFX2
XFILL_5_DFFPOSX1_900 gnd vdd FILL
XFILL_5_DFFPOSX1_922 gnd vdd FILL
XFILL_5_DFFPOSX1_911 gnd vdd FILL
XFILL_5_DFFPOSX1_944 gnd vdd FILL
XFILL_5_DFFPOSX1_955 gnd vdd FILL
XFILL_5_DFFPOSX1_933 gnd vdd FILL
XFILL_5_DFFPOSX1_966 gnd vdd FILL
XFILL_5_DFFPOSX1_977 gnd vdd FILL
XAOI21X1_16 INVX1_33/A INVX2_50/A bundleStartMajId_i[16] gnd AOI21X1_16/Y vdd AOI21X1
XFILL_5_DFFPOSX1_988 gnd vdd FILL
XAOI21X1_38 bundleAddress_i[31] NOR2X1_149/B bundleAddress_i[30] gnd AOI21X1_38/Y
+ vdd AOI21X1
XAOI21X1_27 bundleStartMajId_i[0] OR2X2_14/A BUFX4_156/Y gnd AOI21X1_28/A vdd AOI21X1
XAOI21X1_49 bundleAddress_i[32] OR2X2_20/A bundleAddress_i[31] gnd AOI21X1_49/Y vdd
+ AOI21X1
XFILL_5_DFFPOSX1_999 gnd vdd FILL
XFILL_38_12_0 gnd vdd FILL
XFILL_0_AND2X2_2 gnd vdd FILL
XFILL_4_DFFPOSX1_512 gnd vdd FILL
XFILL_4_DFFPOSX1_501 gnd vdd FILL
XFILL_4_DFFPOSX1_545 gnd vdd FILL
XFILL_4_DFFPOSX1_534 gnd vdd FILL
XFILL_4_DFFPOSX1_523 gnd vdd FILL
XFILL_4_DFFPOSX1_578 gnd vdd FILL
XFILL_4_DFFPOSX1_567 gnd vdd FILL
XFILL_4_DFFPOSX1_589 gnd vdd FILL
XFILL_4_DFFPOSX1_556 gnd vdd FILL
XFILL_27_9_1 gnd vdd FILL
XFILL_2_9_1 gnd vdd FILL
XFILL_26_4_0 gnd vdd FILL
XFILL_1_4_0 gnd vdd FILL
XFILL_1_BUFX2_1003 gnd vdd FILL
XFILL_1_BUFX2_1025 gnd vdd FILL
XFILL_1_BUFX2_1014 gnd vdd FILL
XFILL_1_BUFX2_435 gnd vdd FILL
XFILL_1_BUFX2_413 gnd vdd FILL
XFILL_1_BUFX2_424 gnd vdd FILL
XFILL_1_BUFX2_468 gnd vdd FILL
XFILL_10_8_1 gnd vdd FILL
XFILL_1_BUFX2_457 gnd vdd FILL
XFILL_3_DFFPOSX1_102 gnd vdd FILL
XFILL_1_BUFX2_479 gnd vdd FILL
XOAI21X1_430 INVX1_10/A OR2X2_2/Y OAI21X1_430/C gnd OAI21X1_431/A vdd OAI21X1
XOAI21X1_441 OAI21X1_441/A AOI21X1_1/Y OAI21X1_441/C gnd OAI21X1_441/Y vdd OAI21X1
XFILL_3_DFFPOSX1_124 gnd vdd FILL
XFILL_1_CLKBUF1_26 gnd vdd FILL
XOAI21X1_474 NOR3X1_4/C INVX4_22/Y INVX4_23/Y gnd OAI21X1_474/Y vdd OAI21X1
XFILL_3_DFFPOSX1_135 gnd vdd FILL
XOAI21X1_463 OAI21X1_463/A NOR2X1_37/Y OAI21X1_463/C gnd OAI21X1_463/Y vdd OAI21X1
XFILL_3_DFFPOSX1_146 gnd vdd FILL
XFILL_3_DFFPOSX1_113 gnd vdd FILL
XOAI21X1_452 OAI21X1_452/A NOR2X1_24/Y OAI21X1_452/C gnd OAI21X1_452/Y vdd OAI21X1
XFILL_1_CLKBUF1_37 gnd vdd FILL
XFILL_1_CLKBUF1_15 gnd vdd FILL
XFILL_3_DFFPOSX1_157 gnd vdd FILL
XFILL_3_DFFPOSX1_179 gnd vdd FILL
XFILL_3_DFFPOSX1_168 gnd vdd FILL
XFILL_1_CLKBUF1_59 gnd vdd FILL
XOAI21X1_496 OAI21X1_496/A NOR2X1_56/Y OAI21X1_496/C gnd OAI21X1_496/Y vdd OAI21X1
XOAI21X1_485 AOI21X1_3/Y OAI21X1_485/B OAI21X1_485/C gnd OAI21X1_485/Y vdd OAI21X1
XFILL_1_CLKBUF1_48 gnd vdd FILL
XFILL_9_5_0 gnd vdd FILL
XFILL_2_OAI21X1_162 gnd vdd FILL
XNAND2X1_480 bundleAddress_i[56] bundleAddress_i[55] gnd NOR2X1_180/A vdd NAND2X1
XNAND2X1_491 BUFX2_70/A BUFX4_235/Y gnd NAND2X1_491/Y vdd NAND2X1
XFILL_0_INVX1_201 gnd vdd FILL
XFILL_0_INVX1_212 gnd vdd FILL
XFILL_18_9_1 gnd vdd FILL
XFILL_0_NAND2X1_209 gnd vdd FILL
XFILL_17_4_0 gnd vdd FILL
XFILL_0_INVX1_223 gnd vdd FILL
XFILL_5_DFFPOSX1_207 gnd vdd FILL
XFILL_5_DFFPOSX1_218 gnd vdd FILL
XFILL_5_DFFPOSX1_229 gnd vdd FILL
XFILL_0_OAI21X1_22 gnd vdd FILL
XFILL_0_OAI21X1_33 gnd vdd FILL
XFILL_0_OAI21X1_11 gnd vdd FILL
XFILL_0_OAI21X1_55 gnd vdd FILL
XFILL_1_BUFX2_980 gnd vdd FILL
XOAI21X1_1715 INVX2_119/Y BUFX4_293/Y OAI21X1_1715/C gnd DFFPOSX1_70/D vdd OAI21X1
XFILL_0_OAI21X1_44 gnd vdd FILL
XFILL_1_BUFX2_991 gnd vdd FILL
XFILL_22_10_1 gnd vdd FILL
XOAI21X1_1704 BUFX4_12/Y NAND2X1_7/B BUFX2_735/A gnd OAI21X1_1705/C vdd OAI21X1
XFILL_0_OAI21X1_66 gnd vdd FILL
XOAI21X1_1726 BUFX4_123/Y BUFX4_60/Y BUFX2_775/A gnd OAI21X1_1727/C vdd OAI21X1
XOAI21X1_1737 INVX2_130/Y BUFX4_292/Y OAI21X1_1737/C gnd DFFPOSX1_81/D vdd OAI21X1
XOAI21X1_1748 BUFX4_142/Y BUFX4_77/Y BUFX2_756/A gnd OAI21X1_1749/C vdd OAI21X1
XFILL_0_OAI21X1_99 gnd vdd FILL
XFILL_0_OAI21X1_77 gnd vdd FILL
XFILL_0_OAI21X1_88 gnd vdd FILL
XFILL_3_DFFPOSX1_691 gnd vdd FILL
XFILL_3_DFFPOSX1_680 gnd vdd FILL
XOAI21X1_1759 INVX2_141/Y BUFX4_292/Y OAI21X1_1759/C gnd DFFPOSX1_92/D vdd OAI21X1
XFILL_0_OAI21X1_704 gnd vdd FILL
XFILL_1_OAI21X1_908 gnd vdd FILL
XFILL_0_OAI21X1_715 gnd vdd FILL
XFILL_0_OAI21X1_737 gnd vdd FILL
XFILL_0_OAI21X1_748 gnd vdd FILL
XFILL_0_OAI21X1_726 gnd vdd FILL
XFILL_1_OAI21X1_919 gnd vdd FILL
XFILL_0_OAI21X1_759 gnd vdd FILL
XFILL_0_NAND2X1_710 gnd vdd FILL
XFILL_0_NAND2X1_732 gnd vdd FILL
XFILL_0_NAND2X1_754 gnd vdd FILL
XFILL_0_OAI21X1_1525 gnd vdd FILL
XFILL_0_NAND2X1_721 gnd vdd FILL
XFILL_0_OAI21X1_1514 gnd vdd FILL
XFILL_0_NAND2X1_743 gnd vdd FILL
XFILL_0_OAI21X1_1503 gnd vdd FILL
XFILL_0_NAND2X1_765 gnd vdd FILL
XBUFX2_390 BUFX2_390/A gnd is64b2_o vdd BUFX2
XFILL_2_DFFPOSX1_281 gnd vdd FILL
XFILL_2_DFFPOSX1_292 gnd vdd FILL
XFILL_0_OAI21X1_1558 gnd vdd FILL
XFILL_4_NOR3X1_2 gnd vdd FILL
XFILL_0_OAI21X1_1536 gnd vdd FILL
XFILL_0_OAI21X1_1547 gnd vdd FILL
XFILL_2_DFFPOSX1_270 gnd vdd FILL
XFILL_5_DFFPOSX1_70 gnd vdd FILL
XFILL_5_DFFPOSX1_81 gnd vdd FILL
XFILL_0_OAI21X1_1569 gnd vdd FILL
XFILL_5_DFFPOSX1_92 gnd vdd FILL
XFILL_5_DFFPOSX1_730 gnd vdd FILL
XFILL_5_DFFPOSX1_741 gnd vdd FILL
XOAI21X1_90 BUFX4_94/A BUFX4_340/Y BUFX2_968/A gnd OAI21X1_91/C vdd OAI21X1
XFILL_5_DFFPOSX1_752 gnd vdd FILL
XFILL_5_DFFPOSX1_763 gnd vdd FILL
XFILL_5_DFFPOSX1_774 gnd vdd FILL
XFILL_24_18_0 gnd vdd FILL
XFILL_5_DFFPOSX1_785 gnd vdd FILL
XFILL_5_DFFPOSX1_796 gnd vdd FILL
XFILL_4_DFFPOSX1_320 gnd vdd FILL
XFILL_4_DFFPOSX1_342 gnd vdd FILL
XFILL_4_DFFPOSX1_353 gnd vdd FILL
XFILL_4_DFFPOSX1_331 gnd vdd FILL
XFILL_4_DFFPOSX1_364 gnd vdd FILL
XFILL_2_OAI21X1_1619 gnd vdd FILL
XFILL_2_DFFPOSX1_1012 gnd vdd FILL
XFILL_2_DFFPOSX1_1001 gnd vdd FILL
XFILL_4_DFFPOSX1_375 gnd vdd FILL
XFILL_4_DFFPOSX1_397 gnd vdd FILL
XFILL_2_DFFPOSX1_1023 gnd vdd FILL
XFILL_4_DFFPOSX1_386 gnd vdd FILL
XFILL_2_10_1 gnd vdd FILL
XFILL_29_17_0 gnd vdd FILL
XFILL_1_BUFX2_210 gnd vdd FILL
XFILL_1_BUFX2_232 gnd vdd FILL
XFILL_1_BUFX2_221 gnd vdd FILL
XFILL_1_BUFX2_276 gnd vdd FILL
XFILL_1_BUFX2_265 gnd vdd FILL
XOAI21X1_260 BUFX4_164/Y BUFX4_79/Y BUFX2_993/A gnd OAI21X1_261/C vdd OAI21X1
XFILL_1_OAI21X1_1209 gnd vdd FILL
XOAI21X1_282 BUFX4_128/Y BUFX4_38/Y BUFX2_1005/A gnd OAI21X1_283/C vdd OAI21X1
XOAI21X1_271 INVX2_181/Y BUFX4_290/Y OAI21X1_271/C gnd OAI21X1_271/Y vdd OAI21X1
XOAI21X1_293 INVX2_192/Y BUFX4_302/Y OAI21X1_293/C gnd OAI21X1_293/Y vdd OAI21X1
XFILL_6_DFFPOSX1_414 gnd vdd FILL
XFILL_6_DFFPOSX1_403 gnd vdd FILL
XFILL_6_DFFPOSX1_425 gnd vdd FILL
XFILL_6_DFFPOSX1_458 gnd vdd FILL
XFILL_6_DFFPOSX1_447 gnd vdd FILL
XFILL_6_DFFPOSX1_436 gnd vdd FILL
XFILL_4_18_0 gnd vdd FILL
XFILL_36_4 gnd vdd FILL
XFILL_1_NAND3X1_6 gnd vdd FILL
XFILL_0_INVX8_1 gnd vdd FILL
XFILL_33_7_1 gnd vdd FILL
XFILL_32_2_0 gnd vdd FILL
XFILL_29_3 gnd vdd FILL
XFILL_5_DFFPOSX1_1005 gnd vdd FILL
XFILL_5_DFFPOSX1_1016 gnd vdd FILL
XFILL_5_DFFPOSX1_1027 gnd vdd FILL
XDFFPOSX1_27 BUFX2_697/A CLKBUF1_32/Y DFFPOSX1_27/D gnd vdd DFFPOSX1
XFILL_0_BUFX4_340 gnd vdd FILL
XFILL_0_BUFX4_351 gnd vdd FILL
XOAI21X1_1523 BUFX4_128/Y BUFX4_45/Y BUFX2_234/A gnd OAI21X1_1524/C vdd OAI21X1
XDFFPOSX1_16 BUFX2_685/A CLKBUF1_87/Y DFFPOSX1_16/D gnd vdd DFFPOSX1
XOAI21X1_1512 NAND2X1_639/Y BUFX4_297/Y OAI21X1_1512/C gnd OAI21X1_1512/Y vdd OAI21X1
XOAI21X1_1501 XNOR2X1_101/Y INVX8_2/A OAI21X1_1501/C gnd OAI21X1_1501/Y vdd OAI21X1
XFILL_1_OAI21X1_1710 gnd vdd FILL
XDFFPOSX1_38 BUFX2_725/A CLKBUF1_99/Y DFFPOSX1_38/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1743 gnd vdd FILL
XFILL_1_OAI21X1_1732 gnd vdd FILL
XFILL_0_BUFX4_362 gnd vdd FILL
XDFFPOSX1_49 BUFX2_718/A CLKBUF1_77/Y DFFPOSX1_49/D gnd vdd DFFPOSX1
XOAI21X1_1556 INVX1_226/A INVX2_104/Y INVX1_180/Y gnd NAND3X1_68/C vdd OAI21X1
XFILL_0_BUFX4_373 gnd vdd FILL
XFILL_0_BUFX4_384 gnd vdd FILL
XOAI21X1_1534 BUFX4_152/Y BUFX4_28/Y BUFX2_239/A gnd OAI21X1_1535/C vdd OAI21X1
XFILL_1_OAI21X1_1721 gnd vdd FILL
XOAI21X1_1545 BUFX4_152/Y BUFX4_78/Y BUFX2_242/A gnd OAI21X1_1546/C vdd OAI21X1
XFILL_0_BUFX2_1000 gnd vdd FILL
XOAI21X1_1589 BUFX4_349/Y INVX2_125/Y NAND2X1_658/Y gnd OAI21X1_1589/Y vdd OAI21X1
XFILL_1_OAI21X1_1754 gnd vdd FILL
XFILL_1_OAI21X1_1765 gnd vdd FILL
XOAI21X1_1567 OR2X2_21/Y INVX4_49/Y BUFX4_284/Y gnd OAI21X1_1569/B vdd OAI21X1
XOAI21X1_1578 BUFX4_129/Y INVX2_113/Y OAI21X1_1578/C gnd OAI21X1_1578/Y vdd OAI21X1
XFILL_0_OAI21X1_501 gnd vdd FILL
XFILL_1_OAI21X1_1776 gnd vdd FILL
XFILL_0_OAI21X1_512 gnd vdd FILL
XFILL_0_BUFX2_1011 gnd vdd FILL
XFILL_1_OAI21X1_1798 gnd vdd FILL
XFILL_0_BUFX2_1022 gnd vdd FILL
XFILL_0_OAI21X1_556 gnd vdd FILL
XFILL_1_OAI21X1_716 gnd vdd FILL
XFILL_1_OAI21X1_727 gnd vdd FILL
XFILL_0_OAI21X1_534 gnd vdd FILL
XFILL_0_OAI21X1_545 gnd vdd FILL
XFILL_1_OAI21X1_1787 gnd vdd FILL
XFILL_0_OAI21X1_523 gnd vdd FILL
XFILL_1_OAI21X1_705 gnd vdd FILL
XFILL_1_OAI21X1_738 gnd vdd FILL
XFILL_0_OAI21X1_567 gnd vdd FILL
XFILL_1_OAI21X1_749 gnd vdd FILL
XFILL_0_OAI21X1_578 gnd vdd FILL
XFILL_9_17_0 gnd vdd FILL
XFILL_0_OAI21X1_589 gnd vdd FILL
XFILL_0_CLKBUF1_12 gnd vdd FILL
XFILL_0_CLKBUF1_23 gnd vdd FILL
XFILL_0_CLKBUF1_45 gnd vdd FILL
XFILL_13_15_1 gnd vdd FILL
XFILL_0_CLKBUF1_34 gnd vdd FILL
XFILL_0_CLKBUF1_67 gnd vdd FILL
XFILL_0_CLKBUF1_78 gnd vdd FILL
XFILL_0_OAI21X1_1300 gnd vdd FILL
XFILL_0_CLKBUF1_56 gnd vdd FILL
XFILL_0_NAND2X1_551 gnd vdd FILL
XFILL_0_CLKBUF1_89 gnd vdd FILL
XFILL_1_NAND2X1_722 gnd vdd FILL
XFILL_0_OAI21X1_1333 gnd vdd FILL
XFILL_0_DFFPOSX1_901 gnd vdd FILL
XFILL_0_NAND2X1_562 gnd vdd FILL
XFILL_0_OAI21X1_1311 gnd vdd FILL
XFILL_1_NAND2X1_711 gnd vdd FILL
XFILL_0_OAI21X1_1322 gnd vdd FILL
XFILL_0_NAND2X1_540 gnd vdd FILL
XFILL_0_NAND2X1_595 gnd vdd FILL
XFILL_24_7_1 gnd vdd FILL
XFILL_23_2_0 gnd vdd FILL
XFILL_0_DFFPOSX1_934 gnd vdd FILL
XFILL_0_OAI21X1_1344 gnd vdd FILL
XFILL_0_NAND2X1_584 gnd vdd FILL
XFILL_0_OAI21X1_1366 gnd vdd FILL
XFILL_0_DFFPOSX1_923 gnd vdd FILL
XFILL_0_NAND2X1_573 gnd vdd FILL
XFILL_1_NAND2X1_744 gnd vdd FILL
XFILL_1_NAND2X1_755 gnd vdd FILL
XFILL_0_DFFPOSX1_912 gnd vdd FILL
XFILL_0_OAI21X1_1355 gnd vdd FILL
XFILL_0_OAI21X1_1399 gnd vdd FILL
XFILL_0_DFFPOSX1_967 gnd vdd FILL
XFILL_0_OAI21X1_1388 gnd vdd FILL
XFILL_0_DFFPOSX1_945 gnd vdd FILL
XFILL_0_OAI21X1_1377 gnd vdd FILL
XFILL_0_DFFPOSX1_956 gnd vdd FILL
XFILL_0_DFFPOSX1_978 gnd vdd FILL
XFILL_0_DFFPOSX1_989 gnd vdd FILL
XFILL_5_DFFPOSX1_582 gnd vdd FILL
XFILL_5_DFFPOSX1_560 gnd vdd FILL
XFILL_5_DFFPOSX1_571 gnd vdd FILL
XFILL_0_OR2X2_6 gnd vdd FILL
XFILL_5_DFFPOSX1_593 gnd vdd FILL
XFILL_1_BUFX4_4 gnd vdd FILL
XFILL_18_14_1 gnd vdd FILL
XFILL_7_8_1 gnd vdd FILL
XFILL_2_OAI21X1_1405 gnd vdd FILL
XFILL_6_3_0 gnd vdd FILL
XFILL_4_DFFPOSX1_150 gnd vdd FILL
XFILL_31_16_1 gnd vdd FILL
XCLKBUF1_91 BUFX4_83/Y gnd CLKBUF1_91/Y vdd CLKBUF1
XCLKBUF1_80 BUFX4_83/Y gnd CLKBUF1_80/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_161 gnd vdd FILL
XFILL_4_DFFPOSX1_172 gnd vdd FILL
XFILL_4_DFFPOSX1_194 gnd vdd FILL
XFILL_4_DFFPOSX1_183 gnd vdd FILL
XFILL_2_NOR3X1_16 gnd vdd FILL
XFILL_12_10_0 gnd vdd FILL
XFILL_15_7_1 gnd vdd FILL
XFILL_0_INVX1_8 gnd vdd FILL
XFILL_14_2_0 gnd vdd FILL
XFILL_1_NAND3X1_17 gnd vdd FILL
XFILL_1_NAND3X1_28 gnd vdd FILL
XFILL_0_BUFX2_800 gnd vdd FILL
XFILL_0_BUFX2_811 gnd vdd FILL
XFILL_1_OAI21X1_1028 gnd vdd FILL
XINVX1_110 bundle_i[94] gnd INVX1_110/Y vdd INVX1
XFILL_1_NAND3X1_39 gnd vdd FILL
XFILL_1_OAI21X1_1006 gnd vdd FILL
XFILL_0_BUFX2_833 gnd vdd FILL
XDFFPOSX1_409 BUFX2_442/A CLKBUF1_84/Y OAI21X1_381/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1017 gnd vdd FILL
XFILL_0_BUFX2_822 gnd vdd FILL
XFILL_1_INVX4_4 gnd vdd FILL
XFILL_0_BUFX2_844 gnd vdd FILL
XFILL_1_OAI21X1_1039 gnd vdd FILL
XINVX1_121 bundle_i[83] gnd INVX1_121/Y vdd INVX1
XFILL_0_BUFX2_855 gnd vdd FILL
XFILL_0_BUFX2_866 gnd vdd FILL
XFILL_1_DFFPOSX1_607 gnd vdd FILL
XINVX1_143 bundle_i[125] gnd INVX1_143/Y vdd INVX1
XFILL_1_DFFPOSX1_629 gnd vdd FILL
XFILL_1_DFFPOSX1_618 gnd vdd FILL
XINVX1_132 bundle_i[72] gnd INVX1_132/Y vdd INVX1
XINVX1_154 bundle_i[114] gnd INVX1_154/Y vdd INVX1
XFILL_0_BUFX2_877 gnd vdd FILL
XINVX1_165 bundle_i[103] gnd INVX1_165/Y vdd INVX1
XFILL_6_DFFPOSX1_200 gnd vdd FILL
XINVX1_176 bundleAddress_i[35] gnd INVX1_176/Y vdd INVX1
XFILL_0_BUFX2_899 gnd vdd FILL
XFILL_0_BUFX2_888 gnd vdd FILL
XFILL_6_DFFPOSX1_211 gnd vdd FILL
XINVX1_198 OR2X2_21/B gnd INVX1_198/Y vdd INVX1
XINVX1_187 INVX1_187/A gnd INVX1_187/Y vdd INVX1
XFILL_36_15_1 gnd vdd FILL
XCLKBUF1_102 BUFX4_91/Y gnd CLKBUF1_102/Y vdd CLKBUF1
XFILL_6_DFFPOSX1_299 gnd vdd FILL
XFILL_0_INVX2_20 gnd vdd FILL
XFILL_0_INVX2_64 gnd vdd FILL
XFILL_0_INVX2_53 gnd vdd FILL
XFILL_0_INVX2_31 gnd vdd FILL
XFILL_0_INVX2_42 gnd vdd FILL
XFILL_30_11_0 gnd vdd FILL
XFILL_0_INVX2_75 gnd vdd FILL
XFILL_0_INVX2_97 gnd vdd FILL
XFILL_0_INVX2_86 gnd vdd FILL
XFILL_1_NOR3X1_6 gnd vdd FILL
XFILL_0_DFFPOSX1_208 gnd vdd FILL
XFILL_34_1 gnd vdd FILL
XFILL_0_DFFPOSX1_219 gnd vdd FILL
XOAI21X1_1331 BUFX4_109/Y BUFX4_324/Y BUFX2_169/A gnd OAI21X1_1332/C vdd OAI21X1
XOAI21X1_1320 BUFX4_6/A BUFX4_350/Y BUFX2_165/A gnd OAI21X1_1322/C vdd OAI21X1
XFILL_0_BUFX4_170 gnd vdd FILL
XDFFPOSX1_932 BUFX2_186/A CLKBUF1_97/Y OAI21X1_1375/Y gnd vdd DFFPOSX1
XDFFPOSX1_921 BUFX2_173/A CLKBUF1_36/Y OAI21X1_1344/Y gnd vdd DFFPOSX1
XOAI21X1_1342 BUFX4_96/Y BUFX4_342/Y BUFX2_173/A gnd OAI21X1_1344/C vdd OAI21X1
XOAI21X1_1353 BUFX4_1/A BUFX4_342/Y BUFX2_178/A gnd OAI21X1_1354/C vdd OAI21X1
XFILL_1_OAI21X1_1540 gnd vdd FILL
XDFFPOSX1_910 BUFX2_161/A CLKBUF1_28/Y OAI21X1_1313/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1551 gnd vdd FILL
XFILL_0_BUFX4_181 gnd vdd FILL
XFILL_0_BUFX4_192 gnd vdd FILL
XOAI21X1_1364 OAI21X1_1364/A BUFX4_121/Y OAI21X1_1364/C gnd OAI21X1_1364/Y vdd OAI21X1
XFILL_1_BUFX2_70 gnd vdd FILL
XOAI21X1_1397 NOR2X1_215/B INVX1_185/A OAI21X1_1397/C gnd OAI21X1_1399/A vdd OAI21X1
XFILL_1_OAI21X1_1584 gnd vdd FILL
XDFFPOSX1_954 BUFX2_203/A CLKBUF1_16/Y OAI21X1_1438/Y gnd vdd DFFPOSX1
XDFFPOSX1_943 BUFX2_254/A CLKBUF1_72/Y OAI21X1_1405/Y gnd vdd DFFPOSX1
XOAI21X1_1375 AOI21X1_58/Y NAND2X1_623/Y OAI21X1_1375/C gnd OAI21X1_1375/Y vdd OAI21X1
XOAI21X1_1386 BUFX4_125/Y BUFX4_46/Y BUFX2_194/A gnd OAI21X1_1387/C vdd OAI21X1
XFILL_1_OAI21X1_1573 gnd vdd FILL
XDFFPOSX1_965 BUFX2_215/A CLKBUF1_49/Y OAI21X1_1470/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1562 gnd vdd FILL
XFILL_0_OAI21X1_320 gnd vdd FILL
XFILL_0_OAI21X1_331 gnd vdd FILL
XFILL_1_OAI21X1_502 gnd vdd FILL
XFILL_1_BUFX2_81 gnd vdd FILL
XDFFPOSX1_976 BUFX2_228/A CLKBUF1_76/Y OAI21X1_1505/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1595 gnd vdd FILL
XFILL_1_NOR2X1_129 gnd vdd FILL
XDFFPOSX1_998 BUFX2_252/A CLKBUF1_30/Y OAI21X1_1572/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_364 gnd vdd FILL
XFILL_0_OAI21X1_353 gnd vdd FILL
XFILL_1_OAI21X1_535 gnd vdd FILL
XDFFPOSX1_987 BUFX2_240/A CLKBUF1_28/Y OAI21X1_1539/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_513 gnd vdd FILL
XFILL_0_OAI21X1_342 gnd vdd FILL
XFILL_1_OAI21X1_524 gnd vdd FILL
XFILL_0_OAI21X1_386 gnd vdd FILL
XFILL_1_OAI21X1_568 gnd vdd FILL
XFILL_0_OAI21X1_375 gnd vdd FILL
XFILL_0_OAI21X1_397 gnd vdd FILL
XFILL_1_OAI21X1_557 gnd vdd FILL
XFILL_1_OAI21X1_546 gnd vdd FILL
XFILL_35_10_0 gnd vdd FILL
XFILL_1_OAI21X1_579 gnd vdd FILL
XFILL_1_OAI21X1_3 gnd vdd FILL
XFILL_0_OAI21X1_1130 gnd vdd FILL
XFILL_1_NAND2X1_530 gnd vdd FILL
XFILL_0_NAND2X1_370 gnd vdd FILL
XFILL_1_NAND2X1_541 gnd vdd FILL
XFILL_0_OAI21X1_1141 gnd vdd FILL
XFILL_0_NAND2X1_392 gnd vdd FILL
XFILL_0_DFFPOSX1_742 gnd vdd FILL
XFILL_1_BUFX4_316 gnd vdd FILL
XFILL_0_OAI21X1_1152 gnd vdd FILL
XFILL_1_BUFX4_305 gnd vdd FILL
XFILL_0_OAI21X1_1174 gnd vdd FILL
XFILL_1_NAND2X1_563 gnd vdd FILL
XFILL_1_NAND2X1_585 gnd vdd FILL
XFILL_1_BUFX4_327 gnd vdd FILL
XFILL_0_NAND2X1_381 gnd vdd FILL
XFILL_0_DFFPOSX1_720 gnd vdd FILL
XFILL_0_DFFPOSX1_731 gnd vdd FILL
XFILL_1_BUFX4_338 gnd vdd FILL
XFILL_0_OAI21X1_1163 gnd vdd FILL
XFILL_1_NAND2X1_596 gnd vdd FILL
XFILL_1_BUFX4_349 gnd vdd FILL
XFILL_0_DFFPOSX1_753 gnd vdd FILL
XFILL_0_DFFPOSX1_775 gnd vdd FILL
XFILL_0_OAI21X1_1196 gnd vdd FILL
XFILL_0_OAI21X1_1185 gnd vdd FILL
XFILL_0_DFFPOSX1_764 gnd vdd FILL
XFILL_0_DFFPOSX1_786 gnd vdd FILL
XFILL_0_DFFPOSX1_797 gnd vdd FILL
XFILL_5_DFFPOSX1_390 gnd vdd FILL
XFILL_0_BUFX2_129 gnd vdd FILL
XFILL_0_BUFX2_107 gnd vdd FILL
XFILL_0_BUFX2_118 gnd vdd FILL
XFILL_1_NAND2X1_61 gnd vdd FILL
XINVX4_51 INVX4_51/A gnd INVX4_51/Y vdd INVX4
XINVX4_40 bundleAddress_i[29] gnd INVX4_40/Y vdd INVX4
XFILL_1_NAND2X1_94 gnd vdd FILL
XBUFX2_912 BUFX2_912/A gnd tid3_o[48] vdd BUFX2
XFILL_2_DFFPOSX1_814 gnd vdd FILL
XFILL_2_OAI21X1_1224 gnd vdd FILL
XFILL_2_DFFPOSX1_803 gnd vdd FILL
XBUFX2_901 BUFX2_901/A gnd tid2_o[0] vdd BUFX2
XBUFX2_945 BUFX2_945/A gnd tid3_o[18] vdd BUFX2
XBUFX2_923 BUFX2_923/A gnd tid3_o[38] vdd BUFX2
XFILL_2_DFFPOSX1_90 gnd vdd FILL
XFILL_2_DFFPOSX1_825 gnd vdd FILL
XFILL_2_DFFPOSX1_836 gnd vdd FILL
XBUFX2_934 BUFX2_934/A gnd tid3_o[28] vdd BUFX2
XBUFX2_956 BUFX2_956/A gnd tid3_o[8] vdd BUFX2
XFILL_2_DFFPOSX1_847 gnd vdd FILL
XBUFX2_989 BUFX2_989/A gnd tid4_o[36] vdd BUFX2
XBUFX2_978 BUFX2_978/A gnd tid4_o[46] vdd BUFX2
XFILL_2_DFFPOSX1_869 gnd vdd FILL
XFILL_2_DFFPOSX1_858 gnd vdd FILL
XBUFX2_967 BUFX2_967/A gnd tid3_o[55] vdd BUFX2
XFILL_30_5_1 gnd vdd FILL
XFILL_1_INVX2_1 gnd vdd FILL
XDFFPOSX1_217 BUFX2_890/A CLKBUF1_14/Y OAI21X1_61/Y gnd vdd DFFPOSX1
XDFFPOSX1_228 BUFX2_905/A CLKBUF1_102/Y OAI21X1_73/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_404 gnd vdd FILL
XDFFPOSX1_206 BUFX2_878/A CLKBUF1_51/Y OAI21X1_50/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_641 gnd vdd FILL
XFILL_0_BUFX2_630 gnd vdd FILL
XFILL_1_DFFPOSX1_415 gnd vdd FILL
XDFFPOSX1_239 BUFX2_908/A CLKBUF1_14/Y OAI21X1_95/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_663 gnd vdd FILL
XFILL_0_BUFX2_652 gnd vdd FILL
XFILL_0_BUFX2_685 gnd vdd FILL
XFILL_1_DFFPOSX1_426 gnd vdd FILL
XFILL_0_BUFX2_674 gnd vdd FILL
XFILL_1_DFFPOSX1_448 gnd vdd FILL
XFILL_1_DFFPOSX1_437 gnd vdd FILL
XFILL_0_BUFX2_696 gnd vdd FILL
XFILL_1_DFFPOSX1_459 gnd vdd FILL
XNAND2X1_309 NOR2X1_105/A OAI21X1_679/Y gnd OAI21X1_681/A vdd NAND2X1
XFILL_4_DFFPOSX1_919 gnd vdd FILL
XFILL_4_DFFPOSX1_908 gnd vdd FILL
XNOR3X1_16 INVX4_42/Y NOR3X1_16/B NOR3X1_16/C gnd NOR3X1_16/Y vdd NOR3X1
XFILL_38_6_1 gnd vdd FILL
XFILL_37_1_0 gnd vdd FILL
XBUFX4_282 INVX8_7/Y gnd BUFX4_81/A vdd BUFX4
XBUFX4_260 INVX8_5/Y gnd BUFX4_10/A vdd BUFX4
XBUFX4_271 INVX8_7/Y gnd BUFX4_71/A vdd BUFX4
XFILL_0_INVX2_170 gnd vdd FILL
XFILL_2_OAI21X1_1791 gnd vdd FILL
XBUFX4_293 BUFX4_303/A gnd BUFX4_293/Y vdd BUFX4
XFILL_0_INVX2_181 gnd vdd FILL
XFILL_0_INVX2_192 gnd vdd FILL
XFILL_1_BUFX2_809 gnd vdd FILL
XFILL_0_XNOR2X1_8 gnd vdd FILL
XOAI21X1_804 BUFX4_161/Y BUFX4_52/Y BUFX2_631/A gnd OAI21X1_805/C vdd OAI21X1
XFILL_21_5_1 gnd vdd FILL
XFILL_20_0_0 gnd vdd FILL
XOAI21X1_815 XNOR2X1_54/Y BUFX4_300/Y OAI21X1_815/C gnd OAI21X1_815/Y vdd OAI21X1
XOAI21X1_837 NOR2X1_119/Y OAI21X1_837/B OAI21X1_837/C gnd OAI21X1_837/Y vdd OAI21X1
XOAI21X1_826 XNOR2X1_55/Y BUFX4_289/Y OAI21X1_826/C gnd OAI21X1_826/Y vdd OAI21X1
XFILL_3_DFFPOSX1_509 gnd vdd FILL
XOAI21X1_848 INVX1_49/Y BUFX4_262/Y OAI21X1_848/C gnd OAI21X1_848/Y vdd OAI21X1
XOAI21X1_859 INVX1_60/Y BUFX4_262/Y OAI21X1_859/C gnd OAI21X1_859/Y vdd OAI21X1
XFILL_21_16_0 gnd vdd FILL
XDFFPOSX1_740 BUFX2_378/A CLKBUF1_59/Y OAI21X1_1029/Y gnd vdd DFFPOSX1
XOAI21X1_1150 NAND2X1_529/Y NOR2X1_146/Y NAND2X1_530/Y gnd OAI21X1_1150/Y vdd OAI21X1
XOAI21X1_1172 NAND2X1_554/Y NOR2X1_161/Y NAND2X1_552/Y gnd OAI21X1_1172/Y vdd OAI21X1
XOAI21X1_1161 XNOR2X1_69/Y INVX8_1/A NAND2X1_538/Y gnd OAI21X1_1161/Y vdd OAI21X1
XOAI21X1_1183 NAND2X1_568/Y BUFX4_201/Y NAND2X1_569/Y gnd OAI21X1_1183/Y vdd OAI21X1
XDFFPOSX1_751 BUFX2_62/A CLKBUF1_12/Y OAI21X1_1043/Y gnd vdd DFFPOSX1
XDFFPOSX1_773 BUFX2_23/A CLKBUF1_7/Y OAI21X1_1065/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1392 gnd vdd FILL
XDFFPOSX1_762 BUFX2_11/A CLKBUF1_55/Y OAI21X1_1054/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1381 gnd vdd FILL
XFILL_1_DFFPOSX1_960 gnd vdd FILL
XFILL_1_OAI21X1_310 gnd vdd FILL
XOAI21X1_1194 NOR3X1_14/C OR2X2_21/B BUFX4_242/Y gnd OAI21X1_1195/B vdd OAI21X1
XFILL_1_OAI21X1_1370 gnd vdd FILL
XDFFPOSX1_784 BUFX2_36/A CLKBUF1_53/Y OAI21X1_1076/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_172 gnd vdd FILL
XFILL_0_OAI21X1_161 gnd vdd FILL
XFILL_1_DFFPOSX1_982 gnd vdd FILL
XFILL_0_OAI21X1_150 gnd vdd FILL
XFILL_1_OAI21X1_321 gnd vdd FILL
XFILL_1_DFFPOSX1_993 gnd vdd FILL
XFILL_1_OAI21X1_332 gnd vdd FILL
XFILL_1_DFFPOSX1_971 gnd vdd FILL
XFILL_1_OAI21X1_343 gnd vdd FILL
XDFFPOSX1_795 BUFX2_48/A CLKBUF1_76/Y OAI21X1_1087/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_387 gnd vdd FILL
XFILL_0_OAI21X1_194 gnd vdd FILL
XFILL_1_OAI21X1_354 gnd vdd FILL
XFILL_0_OAI21X1_183 gnd vdd FILL
XFILL_2_OAI21X1_558 gnd vdd FILL
XFILL_2_OAI21X1_547 gnd vdd FILL
XFILL_1_OAI21X1_365 gnd vdd FILL
XFILL_1_OAI21X1_376 gnd vdd FILL
XFILL_2_OAI21X1_536 gnd vdd FILL
XFILL_1_CLKBUF1_8 gnd vdd FILL
XFILL_2_OAI21X1_569 gnd vdd FILL
XFILL_1_OAI21X1_398 gnd vdd FILL
XFILL_29_6_1 gnd vdd FILL
XFILL_28_1_0 gnd vdd FILL
XFILL_0_NAND3X1_36 gnd vdd FILL
XFILL_0_NAND3X1_25 gnd vdd FILL
XFILL_4_6_1 gnd vdd FILL
XFILL_0_NAND3X1_14 gnd vdd FILL
XBUFX2_208 BUFX2_208/A gnd addr4_o[41] vdd BUFX2
XBUFX2_219 BUFX2_219/A gnd addr4_o[31] vdd BUFX2
XFILL_0_NAND3X1_69 gnd vdd FILL
XFILL_0_NAND3X1_58 gnd vdd FILL
XFILL_0_NAND3X1_47 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XFILL_0_BUFX4_60 gnd vdd FILL
XFILL_0_BUFX4_71 gnd vdd FILL
XFILL_0_BUFX4_82 gnd vdd FILL
XFILL_0_BUFX4_93 gnd vdd FILL
XFILL_1_BUFX4_102 gnd vdd FILL
XFILL_1_NAND2X1_360 gnd vdd FILL
XFILL_1_BUFX4_146 gnd vdd FILL
XFILL_1_NAND2X1_371 gnd vdd FILL
XFILL_1_BUFX4_113 gnd vdd FILL
XFILL_1_BUFX4_135 gnd vdd FILL
XFILL_0_DFFPOSX1_550 gnd vdd FILL
XFILL_1_NAND2X1_393 gnd vdd FILL
XFILL_1_BUFX4_124 gnd vdd FILL
XFILL_1_BUFX4_168 gnd vdd FILL
XFILL_26_15_0 gnd vdd FILL
XFILL_1_BUFX4_179 gnd vdd FILL
XFILL_0_DFFPOSX1_583 gnd vdd FILL
XFILL_1_BUFX4_157 gnd vdd FILL
XFILL_0_DFFPOSX1_594 gnd vdd FILL
XFILL_0_DFFPOSX1_572 gnd vdd FILL
XFILL_12_5_1 gnd vdd FILL
XFILL_0_DFFPOSX1_561 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XFILL_2_CLKBUF1_19 gnd vdd FILL
XNAND3X1_60 bundleAddress_i[5] INVX2_103/A NOR2X1_172/Y gnd NOR2X1_210/B vdd NAND3X1
XFILL_2_OAI21X1_1032 gnd vdd FILL
XBUFX2_720 BUFX2_720/A gnd pid3_o[16] vdd BUFX2
XFILL_2_DFFPOSX1_600 gnd vdd FILL
XFILL_2_DFFPOSX1_611 gnd vdd FILL
XFILL_19_1_0 gnd vdd FILL
XFILL_2_DFFPOSX1_622 gnd vdd FILL
XFILL_2_DFFPOSX1_655 gnd vdd FILL
XBUFX2_742 BUFX2_742/A gnd pid3_o[24] vdd BUFX2
XBUFX2_753 BUFX2_753/A gnd pid4_o[15] vdd BUFX2
XBUFX2_764 BUFX2_764/A gnd pid4_o[5] vdd BUFX2
XFILL_2_DFFPOSX1_633 gnd vdd FILL
XBUFX2_731 BUFX2_731/A gnd pid3_o[6] vdd BUFX2
XFILL_2_OAI21X1_1098 gnd vdd FILL
XFILL_3_DFFPOSX1_80 gnd vdd FILL
XNOR2X1_82 OR2X2_2/Y NOR2X1_82/B gnd NOR2X1_82/Y vdd NOR2X1
XFILL_1_16_0 gnd vdd FILL
XFILL_2_DFFPOSX1_644 gnd vdd FILL
XFILL_2_DFFPOSX1_666 gnd vdd FILL
XNOR2X1_60 NOR2X1_60/A NOR2X1_60/B gnd NOR2X1_60/Y vdd NOR2X1
XNOR2X1_71 bundleStartMajId_i[36] NOR2X1_71/B gnd NOR2X1_71/Y vdd NOR2X1
XBUFX2_775 BUFX2_775/A gnd pid4_o[23] vdd BUFX2
XBUFX2_797 BUFX2_797/A gnd tid1_o[36] vdd BUFX2
XBUFX2_786 BUFX2_786/A gnd tid1_o[46] vdd BUFX2
XFILL_3_DFFPOSX1_91 gnd vdd FILL
XFILL_2_DFFPOSX1_688 gnd vdd FILL
XNOR2X1_93 bundleStartMajId_i[13] NOR2X1_93/B gnd NOR2X1_93/Y vdd NOR2X1
XFILL_2_DFFPOSX1_677 gnd vdd FILL
XFILL_2_DFFPOSX1_699 gnd vdd FILL
XFILL_0_NOR2X1_104 gnd vdd FILL
XFILL_0_NOR2X1_126 gnd vdd FILL
XFILL_0_NOR2X1_115 gnd vdd FILL
XFILL_0_NOR2X1_137 gnd vdd FILL
XFILL_0_NOR2X1_148 gnd vdd FILL
XFILL_0_NOR2X1_159 gnd vdd FILL
XFILL_1_DFFPOSX1_212 gnd vdd FILL
XBUFX2_9 BUFX2_9/A gnd addr1_o[47] vdd BUFX2
XFILL_1_DFFPOSX1_201 gnd vdd FILL
XFILL_1_DFFPOSX1_223 gnd vdd FILL
XFILL_1_DFFPOSX1_245 gnd vdd FILL
XFILL_1_DFFPOSX1_234 gnd vdd FILL
XFILL_0_BUFX2_493 gnd vdd FILL
XFILL_0_BUFX2_482 gnd vdd FILL
XFILL_0_BUFX2_460 gnd vdd FILL
XFILL_0_BUFX2_471 gnd vdd FILL
XFILL_1_DFFPOSX1_256 gnd vdd FILL
XFILL_1_DFFPOSX1_278 gnd vdd FILL
XFILL_1_DFFPOSX1_289 gnd vdd FILL
XFILL_1_DFFPOSX1_267 gnd vdd FILL
XNAND2X1_117 BUFX2_433/A BUFX4_345/Y gnd OAI21X1_373/C vdd NAND2X1
XNAND2X1_106 BUFX2_421/A BUFX4_335/Y gnd OAI21X1_362/C vdd NAND2X1
XNAND2X1_128 BUFX2_445/A BUFX4_319/Y gnd OAI21X1_384/C vdd NAND2X1
XNAND2X1_139 bundleStartMajId_i[62] bundleStartMajId_i[61] gnd INVX1_24/A vdd NAND2X1
XFILL_4_DFFPOSX1_716 gnd vdd FILL
XFILL_1_OAI21X1_15 gnd vdd FILL
XFILL_4_DFFPOSX1_727 gnd vdd FILL
XNAND2X1_4 NAND2X1_4/A OAI21X1_4/A gnd OAI21X1_4/C vdd NAND2X1
XFILL_4_DFFPOSX1_738 gnd vdd FILL
XFILL_4_DFFPOSX1_705 gnd vdd FILL
XFILL_6_15_0 gnd vdd FILL
XFILL_4_DFFPOSX1_749 gnd vdd FILL
XFILL_1_OAI21X1_26 gnd vdd FILL
XFILL_1_OAI21X1_48 gnd vdd FILL
XFILL_1_OAI21X1_37 gnd vdd FILL
XFILL_1_OAI21X1_59 gnd vdd FILL
XFILL_10_13_1 gnd vdd FILL
XNOR2X1_150 INVX4_39/Y INVX2_74/Y gnd INVX2_99/A vdd NOR2X1
XNOR2X1_161 NOR2X1_204/A INVX1_194/A gnd NOR2X1_161/Y vdd NOR2X1
XFILL_0_NAND2X1_91 gnd vdd FILL
XFILL_0_NAND2X1_80 gnd vdd FILL
XNOR2X1_183 NOR2X1_183/A INVX1_201/A gnd NOR2X1_183/Y vdd NOR2X1
XNOR2X1_194 INVX1_207/A NOR2X1_194/B gnd NOR2X1_195/B vdd NOR2X1
XNOR2X1_172 INVX2_86/Y INVX2_87/Y gnd NOR2X1_172/Y vdd NOR2X1
XFILL_1_BUFX2_606 gnd vdd FILL
XFILL_1_BUFX2_617 gnd vdd FILL
XFILL_1_BUFX2_639 gnd vdd FILL
XOAI21X1_612 BUFX4_2/A BUFX4_362/Y BUFX2_560/A gnd OAI21X1_614/C vdd OAI21X1
XOAI21X1_623 OAI21X1_623/A AOI21X1_16/Y OAI21X1_623/C gnd OAI21X1_623/Y vdd OAI21X1
XINVX2_9 bundleStartMajId_i[61] gnd INVX2_9/Y vdd INVX2
XOAI21X1_601 BUFX4_10/A BUFX4_383/Y BUFX2_553/A gnd OAI21X1_602/C vdd OAI21X1
XFILL_3_DFFPOSX1_306 gnd vdd FILL
XFILL_3_DFFPOSX1_328 gnd vdd FILL
XOAI21X1_656 OAI21X1_656/A INVX4_28/Y BUFX4_305/Y gnd OAI21X1_657/B vdd OAI21X1
XOAI21X1_645 OAI21X1_645/A INVX4_26/Y BUFX4_305/Y gnd OAI21X1_646/A vdd OAI21X1
XOAI21X1_634 BUFX4_8/Y BUFX4_347/Y BUFX2_570/A gnd OAI21X1_635/C vdd OAI21X1
XFILL_3_DFFPOSX1_317 gnd vdd FILL
XFILL_3_DFFPOSX1_339 gnd vdd FILL
XAOI21X1_9 AOI21X1_9/A OR2X2_7/Y NOR2X1_73/Y gnd AOI21X1_9/Y vdd AOI21X1
XOAI21X1_667 NOR2X1_2/A NOR2X1_3/B OAI21X1_667/C gnd OAI21X1_669/A vdd OAI21X1
XOAI21X1_689 INVX1_35/A OR2X2_1/A INVX4_4/Y gnd OAI21X1_690/C vdd OAI21X1
XOAI21X1_678 NOR2X1_103/Y OAI21X1_678/B OAI21X1_678/C gnd OAI21X1_678/Y vdd OAI21X1
XDFFPOSX1_592 BUFX2_624/A CLKBUF1_84/Y OAI21X1_786/Y gnd vdd DFFPOSX1
XDFFPOSX1_570 BUFX2_600/A CLKBUF1_24/Y OAI21X1_724/Y gnd vdd DFFPOSX1
XDFFPOSX1_581 BUFX2_612/A CLKBUF1_24/Y OAI21X1_754/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_162 gnd vdd FILL
XFILL_1_OAI21X1_140 gnd vdd FILL
XFILL_1_DFFPOSX1_790 gnd vdd FILL
XFILL_1_INVX2_102 gnd vdd FILL
XXNOR2X1_17 NOR2X1_33/Y bundleStartMajId_i[25] gnd XNOR2X1_17/Y vdd XNOR2X1
XXNOR2X1_39 NOR2X1_95/Y bundleStartMajId_i[10] gnd XNOR2X1_39/Y vdd XNOR2X1
XFILL_1_OAI21X1_151 gnd vdd FILL
XFILL_2_OAI21X1_311 gnd vdd FILL
XXNOR2X1_28 OR2X2_10/B INVX4_7/Y gnd XNOR2X1_28/Y vdd XNOR2X1
XFILL_2_OAI21X1_333 gnd vdd FILL
XNAND2X1_673 BUFX2_665/A BUFX4_332/Y gnd NAND2X1_673/Y vdd NAND2X1
XNAND2X1_651 BUFX2_650/A BUFX4_316/Y gnd NAND2X1_651/Y vdd NAND2X1
XFILL_1_OAI21X1_173 gnd vdd FILL
XFILL_1_OAI21X1_184 gnd vdd FILL
XFILL_1_OAI21X1_195 gnd vdd FILL
XNAND2X1_640 bundleAddress_i[17] NOR2X1_226/Y gnd INVX1_225/A vdd NAND2X1
XNAND2X1_662 BUFX2_653/A BUFX4_376/Y gnd NAND2X1_662/Y vdd NAND2X1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XINVX1_30 NOR3X1_5/B gnd INVX1_30/Y vdd INVX1
XFILL_2_OAI21X1_344 gnd vdd FILL
XINVX1_85 bundle_i[55] gnd INVX1_85/Y vdd INVX1
XINVX1_74 INVX1_74/A gnd INVX1_74/Y vdd INVX1
XNAND2X1_684 BUFX2_693/A BUFX4_227/Y gnd NAND2X1_684/Y vdd NAND2X1
XINVX1_63 INVX1_63/A gnd INVX1_63/Y vdd INVX1
XFILL_2_OAI21X1_388 gnd vdd FILL
XNAND2X1_695 BUFX2_686/A INVX8_1/A gnd NAND2X1_695/Y vdd NAND2X1
XFILL_15_12_1 gnd vdd FILL
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XBUFX2_27 BUFX2_27/A gnd addr1_o[31] vdd BUFX2
XINVX1_96 bundle_i[44] gnd INVX1_96/Y vdd INVX1
XBUFX2_16 BUFX2_16/A gnd addr1_o[41] vdd BUFX2
XBUFX2_38 BUFX2_38/A gnd addr1_o[21] vdd BUFX2
XBUFX2_49 BUFX2_49/A gnd addr1_o[11] vdd BUFX2
XDFFPOSX1_4 BUFX2_681/A CLKBUF1_86/Y DFFPOSX1_4/D gnd vdd DFFPOSX1
XFILL_1_BUFX4_16 gnd vdd FILL
XFILL_1_BUFX4_27 gnd vdd FILL
XFILL_0_DFFPOSX1_391 gnd vdd FILL
XFILL_0_DFFPOSX1_380 gnd vdd FILL
XFILL_1_BUFX4_38 gnd vdd FILL
XFILL_1_BUFX4_49 gnd vdd FILL
XFILL_3_DFFPOSX1_840 gnd vdd FILL
XFILL_3_DFFPOSX1_884 gnd vdd FILL
XFILL_3_DFFPOSX1_851 gnd vdd FILL
XFILL_3_DFFPOSX1_873 gnd vdd FILL
XFILL_3_DFFPOSX1_862 gnd vdd FILL
XFILL_0_OAI21X1_908 gnd vdd FILL
XFILL_3_DFFPOSX1_895 gnd vdd FILL
XFILL_0_OAI21X1_919 gnd vdd FILL
XNOR2X1_7 OR2X2_1/A NOR2X1_7/B gnd NOR2X1_7/Y vdd NOR2X1
XFILL_33_13_1 gnd vdd FILL
XFILL_1_INVX1_190 gnd vdd FILL
XFILL_1_OR2X2_19 gnd vdd FILL
XFILL_2_DFFPOSX1_430 gnd vdd FILL
XFILL_0_OAI21X1_1707 gnd vdd FILL
XFILL_2_DFFPOSX1_441 gnd vdd FILL
XFILL_35_4_1 gnd vdd FILL
XFILL_0_OAI21X1_1729 gnd vdd FILL
XFILL_2_DFFPOSX1_463 gnd vdd FILL
XBUFX2_572 BUFX2_572/A gnd majID3_o[8] vdd BUFX2
XFILL_0_OAI21X1_1718 gnd vdd FILL
XBUFX2_561 BUFX2_561/A gnd majID3_o[18] vdd BUFX2
XFILL_2_DFFPOSX1_452 gnd vdd FILL
XBUFX2_550 BUFX2_550/A gnd majID3_o[28] vdd BUFX2
XFILL_2_DFFPOSX1_474 gnd vdd FILL
XFILL_4_DFFPOSX1_70 gnd vdd FILL
XFILL_4_DFFPOSX1_92 gnd vdd FILL
XFILL_4_DFFPOSX1_81 gnd vdd FILL
XFILL_2_DFFPOSX1_485 gnd vdd FILL
XBUFX2_594 BUFX2_594/A gnd majID4_o[46] vdd BUFX2
XBUFX2_583 BUFX2_583/A gnd majID3_o[55] vdd BUFX2
XFILL_2_DFFPOSX1_496 gnd vdd FILL
XFILL_5_DFFPOSX1_901 gnd vdd FILL
XFILL_5_DFFPOSX1_912 gnd vdd FILL
XFILL_5_DFFPOSX1_945 gnd vdd FILL
XFILL_5_DFFPOSX1_934 gnd vdd FILL
XFILL_5_DFFPOSX1_956 gnd vdd FILL
XFILL_5_DFFPOSX1_923 gnd vdd FILL
XFILL_5_DFFPOSX1_967 gnd vdd FILL
XFILL_5_DFFPOSX1_978 gnd vdd FILL
XAOI21X1_17 bundleStartMajId_i[15] OR2X2_11/A BUFX4_122/Y gnd AOI21X1_18/A vdd AOI21X1
XFILL_5_DFFPOSX1_989 gnd vdd FILL
XAOI21X1_28 AOI21X1_28/A OR2X2_14/Y NOR2X1_101/Y gnd AOI21X1_28/Y vdd AOI21X1
XAOI21X1_39 INVX2_111/A NOR2X1_160/Y bundleAddress_i[17] gnd AOI21X1_39/Y vdd AOI21X1
XFILL_0_BUFX2_290 gnd vdd FILL
XFILL_0_AND2X2_3 gnd vdd FILL
XFILL_38_12_1 gnd vdd FILL
XFILL_4_DFFPOSX1_513 gnd vdd FILL
XFILL_4_DFFPOSX1_502 gnd vdd FILL
XFILL_4_DFFPOSX1_546 gnd vdd FILL
XFILL_4_DFFPOSX1_535 gnd vdd FILL
XFILL_4_DFFPOSX1_524 gnd vdd FILL
XFILL_4_DFFPOSX1_568 gnd vdd FILL
XFILL_4_DFFPOSX1_579 gnd vdd FILL
XFILL_4_DFFPOSX1_557 gnd vdd FILL
XFILL_26_4_1 gnd vdd FILL
XFILL_1_4_1 gnd vdd FILL
XFILL_1_BUFX2_1004 gnd vdd FILL
XFILL_1_BUFX2_403 gnd vdd FILL
XFILL_1_BUFX2_414 gnd vdd FILL
XFILL_1_BUFX2_447 gnd vdd FILL
XFILL_3_DFFPOSX1_103 gnd vdd FILL
XFILL_1_BUFX2_458 gnd vdd FILL
XOAI21X1_420 XNOR2X1_3/Y BUFX4_225/Y OAI21X1_420/C gnd OAI21X1_420/Y vdd OAI21X1
XOAI21X1_431 OAI21X1_431/A BUFX4_194/Y OAI21X1_431/C gnd OAI21X1_431/Y vdd OAI21X1
XFILL_3_DFFPOSX1_114 gnd vdd FILL
XFILL_3_DFFPOSX1_125 gnd vdd FILL
XFILL_1_CLKBUF1_16 gnd vdd FILL
XFILL_3_DFFPOSX1_136 gnd vdd FILL
XFILL_1_CLKBUF1_27 gnd vdd FILL
XOAI21X1_475 OAI21X1_475/A BUFX4_183/Y OAI21X1_475/C gnd OAI21X1_475/Y vdd OAI21X1
XOAI21X1_464 XNOR2X1_19/Y BUFX4_183/Y OAI21X1_464/C gnd OAI21X1_464/Y vdd OAI21X1
XOAI21X1_453 XNOR2X1_14/Y BUFX4_236/Y OAI21X1_453/C gnd OAI21X1_453/Y vdd OAI21X1
XOAI21X1_442 NAND3X1_2/Y INVX4_12/Y INVX4_13/Y gnd OAI21X1_442/Y vdd OAI21X1
XFILL_3_DFFPOSX1_147 gnd vdd FILL
XFILL_1_CLKBUF1_49 gnd vdd FILL
XOAI21X1_497 OAI21X1_499/A INVX4_28/Y BUFX4_240/Y gnd OAI21X1_498/A vdd OAI21X1
XOAI21X1_486 NOR2X1_52/Y bundleStartMajId_i[7] BUFX4_240/Y gnd OAI21X1_487/B vdd OAI21X1
XFILL_3_DFFPOSX1_158 gnd vdd FILL
XFILL_3_DFFPOSX1_169 gnd vdd FILL
XFILL_1_CLKBUF1_38 gnd vdd FILL
XFILL_6_DFFPOSX1_607 gnd vdd FILL
XFILL_6_DFFPOSX1_618 gnd vdd FILL
XFILL_6_DFFPOSX1_629 gnd vdd FILL
XFILL_9_5_1 gnd vdd FILL
XFILL_8_0_0 gnd vdd FILL
XNAND2X1_481 BUFX4_241/Y NAND2X1_481/B gnd NAND2X1_481/Y vdd NAND2X1
XNAND2X1_470 bundleAddress_i[60] bundleAddress_i[59] gnd INVX1_183/A vdd NAND2X1
XNAND2X1_492 INVX2_66/Y NAND2X1_492/B gnd NAND2X1_492/Y vdd NAND2X1
XFILL_0_INVX1_213 gnd vdd FILL
XFILL_0_INVX1_202 gnd vdd FILL
XFILL_0_INVX1_224 gnd vdd FILL
XFILL_17_4_1 gnd vdd FILL
XFILL_5_DFFPOSX1_208 gnd vdd FILL
XFILL_5_DFFPOSX1_219 gnd vdd FILL
XFILL_0_OAI21X1_23 gnd vdd FILL
XFILL_0_OAI21X1_12 gnd vdd FILL
XFILL_0_OAI21X1_34 gnd vdd FILL
XFILL_0_OAI21X1_56 gnd vdd FILL
XFILL_0_OAI21X1_45 gnd vdd FILL
XOAI21X1_1705 BUFX4_144/Y INVX2_114/Y OAI21X1_1705/C gnd DFFPOSX1_65/D vdd OAI21X1
XFILL_1_BUFX2_970 gnd vdd FILL
XFILL_1_BUFX2_981 gnd vdd FILL
XOAI21X1_1727 INVX2_125/Y BUFX4_293/Y OAI21X1_1727/C gnd DFFPOSX1_76/D vdd OAI21X1
XOAI21X1_1738 BUFX4_128/Y BUFX4_38/Y BUFX2_751/A gnd OAI21X1_1739/C vdd OAI21X1
XOAI21X1_1716 BUFX4_129/Y BUFX4_80/Y BUFX2_768/A gnd OAI21X1_1717/C vdd OAI21X1
XFILL_0_OAI21X1_78 gnd vdd FILL
XFILL_0_OAI21X1_67 gnd vdd FILL
XFILL_0_OAI21X1_89 gnd vdd FILL
XFILL_3_DFFPOSX1_670 gnd vdd FILL
XFILL_3_DFFPOSX1_692 gnd vdd FILL
XFILL_3_DFFPOSX1_681 gnd vdd FILL
XOAI21X1_1749 INVX2_136/Y BUFX4_300/Y OAI21X1_1749/C gnd DFFPOSX1_87/D vdd OAI21X1
XFILL_0_OAI21X1_705 gnd vdd FILL
XFILL_1_OAI21X1_909 gnd vdd FILL
XFILL_0_OAI21X1_738 gnd vdd FILL
XFILL_0_OAI21X1_716 gnd vdd FILL
XFILL_0_OAI21X1_727 gnd vdd FILL
XFILL_0_OAI21X1_749 gnd vdd FILL
XFILL_0_NAND2X1_700 gnd vdd FILL
XFILL_0_NAND2X1_711 gnd vdd FILL
XFILL_0_NAND2X1_733 gnd vdd FILL
XFILL_0_OAI21X1_1515 gnd vdd FILL
XFILL_0_NAND2X1_722 gnd vdd FILL
XFILL_0_NAND2X1_744 gnd vdd FILL
XFILL_0_OAI21X1_1504 gnd vdd FILL
XBUFX2_380 BUFX2_380/A gnd instr4_o[28] vdd BUFX2
XFILL_2_DFFPOSX1_282 gnd vdd FILL
XFILL_2_DFFPOSX1_271 gnd vdd FILL
XFILL_0_OAI21X1_1526 gnd vdd FILL
XFILL_0_NAND2X1_766 gnd vdd FILL
XFILL_4_NOR3X1_3 gnd vdd FILL
XFILL_0_OAI21X1_1537 gnd vdd FILL
XFILL_0_NAND2X1_755 gnd vdd FILL
XFILL_2_DFFPOSX1_260 gnd vdd FILL
XFILL_0_OAI21X1_1548 gnd vdd FILL
XFILL_5_DFFPOSX1_82 gnd vdd FILL
XFILL_5_DFFPOSX1_60 gnd vdd FILL
XFILL_5_DFFPOSX1_71 gnd vdd FILL
XFILL_0_OAI21X1_1559 gnd vdd FILL
XBUFX2_391 BUFX2_391/A gnd is64b3_o vdd BUFX2
XFILL_2_DFFPOSX1_293 gnd vdd FILL
XFILL_5_DFFPOSX1_93 gnd vdd FILL
XFILL_5_DFFPOSX1_720 gnd vdd FILL
XOAI21X1_80 BUFX4_94/Y BUFX4_312/Y BUFX2_939/A gnd OAI21X1_81/C vdd OAI21X1
XFILL_5_DFFPOSX1_742 gnd vdd FILL
XFILL_5_DFFPOSX1_753 gnd vdd FILL
XFILL_5_DFFPOSX1_731 gnd vdd FILL
XFILL_5_DFFPOSX1_764 gnd vdd FILL
XOAI21X1_91 BUFX4_150/Y INVX2_155/Y OAI21X1_91/C gnd OAI21X1_91/Y vdd OAI21X1
XFILL_5_DFFPOSX1_775 gnd vdd FILL
XFILL_24_18_1 gnd vdd FILL
XFILL_5_DFFPOSX1_786 gnd vdd FILL
XFILL_5_DFFPOSX1_797 gnd vdd FILL
XFILL_4_DFFPOSX1_321 gnd vdd FILL
XFILL_4_DFFPOSX1_310 gnd vdd FILL
XFILL_4_DFFPOSX1_343 gnd vdd FILL
XFILL_4_DFFPOSX1_354 gnd vdd FILL
XFILL_4_DFFPOSX1_332 gnd vdd FILL
XFILL_2_DFFPOSX1_1013 gnd vdd FILL
XFILL_2_DFFPOSX1_1002 gnd vdd FILL
XFILL_4_DFFPOSX1_365 gnd vdd FILL
XFILL_4_DFFPOSX1_376 gnd vdd FILL
XFILL_4_DFFPOSX1_387 gnd vdd FILL
XFILL_2_DFFPOSX1_1024 gnd vdd FILL
XFILL_4_DFFPOSX1_398 gnd vdd FILL
XFILL_29_17_1 gnd vdd FILL
XFILL_1_BUFX2_211 gnd vdd FILL
XFILL_1_BUFX2_200 gnd vdd FILL
XFILL_1_BUFX2_244 gnd vdd FILL
XFILL_1_BUFX2_255 gnd vdd FILL
XOAI21X1_250 BUFX4_138/Y BUFX4_40/Y BUFX2_987/A gnd OAI21X1_251/C vdd OAI21X1
XFILL_1_BUFX2_266 gnd vdd FILL
XFILL_23_13_0 gnd vdd FILL
XFILL_1_BUFX2_299 gnd vdd FILL
XOAI21X1_261 INVX2_176/Y BUFX4_291/Y OAI21X1_261/C gnd OAI21X1_261/Y vdd OAI21X1
XOAI21X1_272 BUFX4_148/Y BUFX4_55/Y BUFX2_999/A gnd OAI21X1_273/C vdd OAI21X1
XOAI21X1_283 INVX2_187/Y BUFX4_301/Y OAI21X1_283/C gnd OAI21X1_283/Y vdd OAI21X1
XFILL_1_BUFX2_288 gnd vdd FILL
XOAI21X1_294 BUFX4_159/Y BUFX4_71/Y BUFX2_1011/A gnd OAI21X1_295/C vdd OAI21X1
XFILL_4_18_1 gnd vdd FILL
XFILL_0_INVX8_2 gnd vdd FILL
XFILL_1_NAND3X1_7 gnd vdd FILL
XFILL_29_4 gnd vdd FILL
XFILL_32_2_1 gnd vdd FILL
XFILL_28_12_0 gnd vdd FILL
XFILL_5_DFFPOSX1_1006 gnd vdd FILL
XFILL_5_DFFPOSX1_1017 gnd vdd FILL
XFILL_5_DFFPOSX1_1028 gnd vdd FILL
XFILL_1_OAI21X1_1700 gnd vdd FILL
XFILL_0_BUFX4_352 gnd vdd FILL
XFILL_0_BUFX4_341 gnd vdd FILL
XFILL_0_BUFX4_330 gnd vdd FILL
XDFFPOSX1_17 BUFX2_686/A CLKBUF1_49/Y DFFPOSX1_17/D gnd vdd DFFPOSX1
XOAI21X1_1513 BUFX4_121/Y BUFX4_58/Y BUFX2_231/A gnd OAI21X1_1514/C vdd OAI21X1
XOAI21X1_1502 NAND3X1_65/Y INVX8_3/Y INVX2_79/Y gnd OAI21X1_1503/C vdd OAI21X1
XFILL_1_OAI21X1_1711 gnd vdd FILL
XFILL_0_BUFX4_363 gnd vdd FILL
XFILL_0_BUFX4_385 gnd vdd FILL
XDFFPOSX1_39 BUFX2_736/A CLKBUF1_7/Y DFFPOSX1_39/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1733 gnd vdd FILL
XOAI21X1_1524 NAND2X1_641/Y BUFX4_297/Y OAI21X1_1524/C gnd OAI21X1_1524/Y vdd OAI21X1
XOAI21X1_1557 INVX1_227/Y BUFX4_286/Y NAND3X1_68/Y gnd OAI21X1_1557/Y vdd OAI21X1
XOAI21X1_1546 OAI21X1_1546/A BUFX4_294/Y OAI21X1_1546/C gnd OAI21X1_1546/Y vdd OAI21X1
XOAI21X1_1535 XNOR2X1_103/Y BUFX4_294/Y OAI21X1_1535/C gnd OAI21X1_1535/Y vdd OAI21X1
XDFFPOSX1_28 BUFX2_698/A CLKBUF1_52/Y DFFPOSX1_28/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1722 gnd vdd FILL
XFILL_0_BUFX4_374 gnd vdd FILL
XFILL_0_BUFX2_1001 gnd vdd FILL
XFILL_1_OAI21X1_1755 gnd vdd FILL
XFILL_1_OAI21X1_1744 gnd vdd FILL
XFILL_1_OAI21X1_1766 gnd vdd FILL
XOAI21X1_1568 BUFX4_121/Y BUFX4_47/Y BUFX2_251/A gnd OAI21X1_1569/C vdd OAI21X1
XOAI21X1_1579 BUFX4_129/Y BUFX4_35/Y BUFX2_392/A gnd OAI21X1_1580/C vdd OAI21X1
XFILL_0_OAI21X1_502 gnd vdd FILL
XFILL_0_OAI21X1_513 gnd vdd FILL
XFILL_1_OAI21X1_1788 gnd vdd FILL
XFILL_1_OAI21X1_1799 gnd vdd FILL
XFILL_0_BUFX2_1012 gnd vdd FILL
XFILL_1_OAI21X1_717 gnd vdd FILL
XFILL_0_OAI21X1_535 gnd vdd FILL
XFILL_1_OAI21X1_1777 gnd vdd FILL
XFILL_1_OAI21X1_706 gnd vdd FILL
XFILL_0_OAI21X1_546 gnd vdd FILL
XFILL_0_BUFX2_1023 gnd vdd FILL
XFILL_0_OAI21X1_524 gnd vdd FILL
XFILL_0_OAI21X1_568 gnd vdd FILL
XFILL_0_OAI21X1_579 gnd vdd FILL
XFILL_1_OAI21X1_728 gnd vdd FILL
XFILL_1_OAI21X1_739 gnd vdd FILL
XFILL_0_OAI21X1_557 gnd vdd FILL
XFILL_9_17_1 gnd vdd FILL
XFILL_6_DFFPOSX1_982 gnd vdd FILL
XFILL_6_DFFPOSX1_960 gnd vdd FILL
XFILL_6_DFFPOSX1_971 gnd vdd FILL
XFILL_6_DFFPOSX1_993 gnd vdd FILL
XFILL_0_CLKBUF1_35 gnd vdd FILL
XFILL_0_CLKBUF1_24 gnd vdd FILL
XFILL_0_CLKBUF1_13 gnd vdd FILL
XFILL_0_CLKBUF1_57 gnd vdd FILL
XFILL_0_CLKBUF1_68 gnd vdd FILL
XFILL_0_CLKBUF1_79 gnd vdd FILL
XFILL_3_13_0 gnd vdd FILL
XFILL_0_CLKBUF1_46 gnd vdd FILL
XFILL_1_NAND2X1_734 gnd vdd FILL
XFILL_0_NAND2X1_530 gnd vdd FILL
XFILL_0_NAND2X1_552 gnd vdd FILL
XFILL_0_OAI21X1_1301 gnd vdd FILL
XFILL_0_OAI21X1_1323 gnd vdd FILL
XFILL_0_OAI21X1_1312 gnd vdd FILL
XFILL_0_NAND2X1_541 gnd vdd FILL
XFILL_1_NAND2X1_723 gnd vdd FILL
XFILL_0_NAND2X1_596 gnd vdd FILL
XFILL_0_DFFPOSX1_902 gnd vdd FILL
XFILL_0_OAI21X1_1334 gnd vdd FILL
XFILL_0_NAND2X1_563 gnd vdd FILL
XFILL_0_NAND2X1_585 gnd vdd FILL
XFILL_0_OAI21X1_1345 gnd vdd FILL
XFILL_0_DFFPOSX1_924 gnd vdd FILL
XFILL_0_OAI21X1_1367 gnd vdd FILL
XFILL_0_NAND2X1_574 gnd vdd FILL
XFILL_0_OAI21X1_1356 gnd vdd FILL
XFILL_1_NAND2X1_767 gnd vdd FILL
XFILL_1_NAND2X1_756 gnd vdd FILL
XFILL_0_DFFPOSX1_913 gnd vdd FILL
XFILL_6_DFFPOSX1_50 gnd vdd FILL
XFILL_0_DFFPOSX1_946 gnd vdd FILL
XFILL_0_DFFPOSX1_968 gnd vdd FILL
XFILL_0_OAI21X1_1389 gnd vdd FILL
XFILL_6_DFFPOSX1_61 gnd vdd FILL
XFILL_23_2_1 gnd vdd FILL
XFILL_0_DFFPOSX1_935 gnd vdd FILL
XFILL_0_OAI21X1_1378 gnd vdd FILL
XFILL_0_DFFPOSX1_957 gnd vdd FILL
XFILL_6_DFFPOSX1_94 gnd vdd FILL
XFILL_6_DFFPOSX1_83 gnd vdd FILL
XFILL_6_DFFPOSX1_72 gnd vdd FILL
XFILL_0_DFFPOSX1_979 gnd vdd FILL
XFILL_5_DFFPOSX1_550 gnd vdd FILL
XFILL_5_DFFPOSX1_572 gnd vdd FILL
XFILL_5_DFFPOSX1_561 gnd vdd FILL
XFILL_5_DFFPOSX1_583 gnd vdd FILL
XFILL_0_OR2X2_7 gnd vdd FILL
XFILL_5_DFFPOSX1_594 gnd vdd FILL
XFILL_1_BUFX4_5 gnd vdd FILL
XFILL_1_AOI21X1_1 gnd vdd FILL
XFILL_8_12_0 gnd vdd FILL
XFILL_6_3_1 gnd vdd FILL
XCLKBUF1_70 BUFX4_84/Y gnd CLKBUF1_70/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_151 gnd vdd FILL
XFILL_4_DFFPOSX1_162 gnd vdd FILL
XCLKBUF1_81 BUFX4_89/Y gnd CLKBUF1_81/Y vdd CLKBUF1
XCLKBUF1_92 BUFX4_84/Y gnd CLKBUF1_92/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_140 gnd vdd FILL
XFILL_1_DFFPOSX1_90 gnd vdd FILL
XFILL_4_DFFPOSX1_195 gnd vdd FILL
XFILL_4_DFFPOSX1_173 gnd vdd FILL
XFILL_2_NOR3X1_17 gnd vdd FILL
XFILL_12_10_1 gnd vdd FILL
XFILL_4_DFFPOSX1_184 gnd vdd FILL
XFILL_2_BUFX4_261 gnd vdd FILL
XFILL_0_INVX1_9 gnd vdd FILL
XFILL_14_2_1 gnd vdd FILL
XFILL_1_NAND3X1_18 gnd vdd FILL
XFILL_0_BUFX2_801 gnd vdd FILL
XFILL_1_OAI21X1_1029 gnd vdd FILL
XFILL_0_BUFX2_823 gnd vdd FILL
XFILL_1_OAI21X1_1007 gnd vdd FILL
XFILL_1_OAI21X1_1018 gnd vdd FILL
XFILL_1_NAND3X1_29 gnd vdd FILL
XFILL_0_BUFX2_834 gnd vdd FILL
XINVX1_100 bundle_i[40] gnd INVX1_100/Y vdd INVX1
XFILL_0_BUFX2_812 gnd vdd FILL
XFILL_1_INVX4_5 gnd vdd FILL
XINVX1_133 bundle_i[71] gnd INVX1_133/Y vdd INVX1
XFILL_0_BUFX2_845 gnd vdd FILL
XFILL_0_BUFX2_856 gnd vdd FILL
XFILL_1_DFFPOSX1_608 gnd vdd FILL
XFILL_0_BUFX2_867 gnd vdd FILL
XFILL_1_DFFPOSX1_619 gnd vdd FILL
XINVX1_122 bundle_i[82] gnd INVX1_122/Y vdd INVX1
XINVX1_111 bundle_i[93] gnd INVX1_111/Y vdd INVX1
XINVX1_144 bundle_i[124] gnd INVX1_144/Y vdd INVX1
XINVX1_166 bundle_i[102] gnd INVX1_166/Y vdd INVX1
XINVX1_177 bundleAddress_i[19] gnd INVX1_177/Y vdd INVX1
XINVX1_155 bundle_i[113] gnd INVX1_155/Y vdd INVX1
XFILL_0_BUFX2_889 gnd vdd FILL
XFILL_0_BUFX2_878 gnd vdd FILL
XFILL_6_DFFPOSX1_234 gnd vdd FILL
XINVX1_188 INVX1_188/A gnd INVX1_188/Y vdd INVX1
XINVX1_199 INVX1_199/A gnd INVX1_199/Y vdd INVX1
XFILL_6_DFFPOSX1_245 gnd vdd FILL
XFILL_6_DFFPOSX1_267 gnd vdd FILL
XFILL_6_DFFPOSX1_256 gnd vdd FILL
XFILL_6_DFFPOSX1_278 gnd vdd FILL
XFILL_6_DFFPOSX1_289 gnd vdd FILL
XFILL_0_INVX2_10 gnd vdd FILL
XFILL_0_INVX2_21 gnd vdd FILL
XFILL_0_INVX2_54 gnd vdd FILL
XFILL_0_INVX2_32 gnd vdd FILL
XFILL_14_18_0 gnd vdd FILL
XFILL_0_INVX2_43 gnd vdd FILL
XFILL_30_11_1 gnd vdd FILL
XFILL_0_INVX2_65 gnd vdd FILL
XFILL_0_INVX2_98 gnd vdd FILL
XFILL_0_INVX2_87 gnd vdd FILL
XFILL_0_INVX2_76 gnd vdd FILL
XFILL_1_NOR3X1_7 gnd vdd FILL
XFILL_0_DFFPOSX1_209 gnd vdd FILL
XFILL_34_2 gnd vdd FILL
XFILL_27_1 gnd vdd FILL
XFILL_0_BUFX4_160 gnd vdd FILL
XOAI21X1_1332 XNOR2X1_85/Y BUFX4_157/Y OAI21X1_1332/C gnd OAI21X1_1332/Y vdd OAI21X1
XOAI21X1_1310 BUFX4_6/A BUFX4_370/Y BUFX2_160/A gnd OAI21X1_1311/C vdd OAI21X1
XOAI21X1_1321 NAND2X1_612/Y INVX4_42/Y BUFX4_308/Y gnd OAI21X1_1322/A vdd OAI21X1
XFILL_0_BUFX4_193 gnd vdd FILL
XFILL_0_BUFX4_171 gnd vdd FILL
XDFFPOSX1_900 BUFX2_150/A CLKBUF1_55/Y OAI21X1_1287/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1530 gnd vdd FILL
XOAI21X1_1343 INVX1_213/A INVX2_83/Y BUFX4_310/Y gnd OAI21X1_1344/B vdd OAI21X1
XDFFPOSX1_922 BUFX2_175/A CLKBUF1_85/Y OAI21X1_1347/Y gnd vdd DFFPOSX1
XDFFPOSX1_933 BUFX2_187/A CLKBUF1_69/Y OAI21X1_1378/Y gnd vdd DFFPOSX1
XOAI21X1_1354 XNOR2X1_87/Y BUFX4_121/Y OAI21X1_1354/C gnd OAI21X1_1354/Y vdd OAI21X1
XOAI21X1_1365 BUFX4_1/A BUFX4_357/Y BUFX2_182/A gnd OAI21X1_1367/C vdd OAI21X1
XFILL_1_OAI21X1_1541 gnd vdd FILL
XFILL_0_BUFX4_182 gnd vdd FILL
XDFFPOSX1_911 BUFX2_162/A CLKBUF1_62/Y OAI21X1_1315/Y gnd vdd DFFPOSX1
XFILL_1_BUFX2_71 gnd vdd FILL
XOAI21X1_1398 BUFX4_126/Y BUFX4_29/Y BUFX2_238/A gnd OAI21X1_1399/C vdd OAI21X1
XDFFPOSX1_944 BUFX2_255/A CLKBUF1_31/Y OAI21X1_1408/Y gnd vdd DFFPOSX1
XFILL_1_BUFX2_60 gnd vdd FILL
XDFFPOSX1_966 BUFX2_217/A CLKBUF1_27/Y OAI21X1_1473/Y gnd vdd DFFPOSX1
XOAI21X1_1387 INVX2_55/Y BUFX4_296/Y OAI21X1_1387/C gnd OAI21X1_1387/Y vdd OAI21X1
XFILL_1_OAI21X1_1574 gnd vdd FILL
XDFFPOSX1_955 BUFX2_204/A CLKBUF1_60/Y OAI21X1_1442/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1563 gnd vdd FILL
XFILL_0_OAI21X1_310 gnd vdd FILL
XFILL_1_OAI21X1_1585 gnd vdd FILL
XOAI21X1_1376 BUFX4_105/Y BUFX4_357/Y BUFX2_187/A gnd OAI21X1_1378/C vdd OAI21X1
XFILL_0_OAI21X1_321 gnd vdd FILL
XFILL_1_OAI21X1_1552 gnd vdd FILL
XFILL_1_OAI21X1_1596 gnd vdd FILL
XFILL_1_NOR2X1_119 gnd vdd FILL
XFILL_1_OAI21X1_525 gnd vdd FILL
XDFFPOSX1_999 BUFX2_253/A CLKBUF1_97/Y OAI21X1_1574/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_354 gnd vdd FILL
XDFFPOSX1_977 BUFX2_229/A CLKBUF1_85/Y OAI21X1_1509/Y gnd vdd DFFPOSX1
XDFFPOSX1_988 BUFX2_241/A CLKBUF1_85/Y OAI21X1_1542/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_503 gnd vdd FILL
XFILL_1_BUFX2_93 gnd vdd FILL
XFILL_1_NOR2X1_108 gnd vdd FILL
XFILL_1_OAI21X1_536 gnd vdd FILL
XFILL_1_OAI21X1_514 gnd vdd FILL
XFILL_0_OAI21X1_332 gnd vdd FILL
XFILL_0_OAI21X1_343 gnd vdd FILL
XFILL_0_OAI21X1_387 gnd vdd FILL
XFILL_19_17_0 gnd vdd FILL
XFILL_1_OAI21X1_569 gnd vdd FILL
XFILL_1_OAI21X1_558 gnd vdd FILL
XFILL_0_OAI21X1_398 gnd vdd FILL
XFILL_1_OAI21X1_547 gnd vdd FILL
XFILL_0_OAI21X1_365 gnd vdd FILL
XFILL_0_OAI21X1_376 gnd vdd FILL
XFILL_35_10_1 gnd vdd FILL
XFILL_1_OAI21X1_4 gnd vdd FILL
XFILL_1_NAND2X1_531 gnd vdd FILL
XFILL_0_OAI21X1_1131 gnd vdd FILL
XFILL_0_OAI21X1_1120 gnd vdd FILL
XFILL_0_NAND2X1_371 gnd vdd FILL
XFILL_1_NAND2X1_520 gnd vdd FILL
XFILL_0_NAND2X1_360 gnd vdd FILL
XFILL_0_OAI21X1_1142 gnd vdd FILL
XFILL_1_NAND2X1_542 gnd vdd FILL
XFILL_0_DFFPOSX1_710 gnd vdd FILL
XFILL_0_NAND2X1_382 gnd vdd FILL
XFILL_0_DFFPOSX1_721 gnd vdd FILL
XFILL_0_OAI21X1_1153 gnd vdd FILL
XFILL_1_BUFX4_328 gnd vdd FILL
XFILL_0_OAI21X1_1175 gnd vdd FILL
XFILL_1_BUFX4_317 gnd vdd FILL
XFILL_1_NAND2X1_553 gnd vdd FILL
XFILL_0_DFFPOSX1_743 gnd vdd FILL
XFILL_1_NAND2X1_564 gnd vdd FILL
XFILL_1_BUFX4_306 gnd vdd FILL
XFILL_1_NAND2X1_575 gnd vdd FILL
XFILL_0_NAND2X1_393 gnd vdd FILL
XFILL_0_DFFPOSX1_732 gnd vdd FILL
XFILL_0_OAI21X1_1164 gnd vdd FILL
XFILL_1_NAND2X1_597 gnd vdd FILL
XFILL_0_DFFPOSX1_754 gnd vdd FILL
XFILL_0_DFFPOSX1_776 gnd vdd FILL
XFILL_1_BUFX4_339 gnd vdd FILL
XFILL_0_OAI21X1_1197 gnd vdd FILL
XFILL_1_NAND2X1_586 gnd vdd FILL
XFILL_0_OAI21X1_1186 gnd vdd FILL
XFILL_0_DFFPOSX1_765 gnd vdd FILL
XFILL_0_DFFPOSX1_787 gnd vdd FILL
XFILL_0_DFFPOSX1_798 gnd vdd FILL
XFILL_2_OAI21X1_19 gnd vdd FILL
XFILL_5_DFFPOSX1_380 gnd vdd FILL
XFILL_0_BUFX2_108 gnd vdd FILL
XFILL_0_BUFX2_119 gnd vdd FILL
XFILL_5_DFFPOSX1_391 gnd vdd FILL
XFILL_1_NAND2X1_40 gnd vdd FILL
XFILL_1_NAND2X1_62 gnd vdd FILL
XFILL_1_NAND2X1_51 gnd vdd FILL
XFILL_1_NAND2X1_73 gnd vdd FILL
XFILL_1_NAND2X1_84 gnd vdd FILL
XINVX4_41 bundleAddress_i[26] gnd INVX4_41/Y vdd INVX4
XINVX4_30 INVX4_30/A gnd INVX4_30/Y vdd INVX4
XFILL_1_NAND2X1_95 gnd vdd FILL
XFILL_37_18_0 gnd vdd FILL
XFILL_1_BUFX2_2 gnd vdd FILL
XFILL_2_DFFPOSX1_815 gnd vdd FILL
XBUFX2_913 BUFX2_913/A gnd tid3_o[47] vdd BUFX2
XBUFX2_902 BUFX2_902/A gnd tid2_o[56] vdd BUFX2
XFILL_2_DFFPOSX1_804 gnd vdd FILL
XBUFX2_924 BUFX2_924/A gnd tid3_o[37] vdd BUFX2
XFILL_2_DFFPOSX1_91 gnd vdd FILL
XFILL_2_DFFPOSX1_837 gnd vdd FILL
XBUFX2_935 BUFX2_935/A gnd tid3_o[27] vdd BUFX2
XFILL_2_DFFPOSX1_80 gnd vdd FILL
XBUFX2_946 BUFX2_946/A gnd tid3_o[17] vdd BUFX2
XFILL_2_DFFPOSX1_848 gnd vdd FILL
XFILL_2_DFFPOSX1_826 gnd vdd FILL
XBUFX2_957 BUFX2_957/A gnd tid3_o[7] vdd BUFX2
XBUFX2_968 BUFX2_968/A gnd tid3_o[54] vdd BUFX2
XBUFX2_979 BUFX2_979/A gnd tid4_o[45] vdd BUFX2
XFILL_2_DFFPOSX1_859 gnd vdd FILL
XDFFPOSX1_218 BUFX2_891/A CLKBUF1_98/Y OAI21X1_62/Y gnd vdd DFFPOSX1
XDFFPOSX1_207 BUFX2_879/A CLKBUF1_42/Y OAI21X1_51/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_405 gnd vdd FILL
XFILL_0_BUFX2_631 gnd vdd FILL
XFILL_0_BUFX2_620 gnd vdd FILL
XFILL_0_BUFX2_642 gnd vdd FILL
XFILL_0_BUFX2_664 gnd vdd FILL
XDFFPOSX1_229 BUFX2_906/A CLKBUF1_27/Y OAI21X1_75/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_416 gnd vdd FILL
XFILL_0_BUFX2_653 gnd vdd FILL
XFILL_0_BUFX2_675 gnd vdd FILL
XFILL_1_DFFPOSX1_427 gnd vdd FILL
XFILL_1_DFFPOSX1_438 gnd vdd FILL
XFILL_0_BUFX2_697 gnd vdd FILL
XFILL_0_BUFX2_686 gnd vdd FILL
XFILL_1_DFFPOSX1_449 gnd vdd FILL
XFILL_4_DFFPOSX1_909 gnd vdd FILL
XNOR3X1_17 NOR3X1_18/A NOR3X1_17/B NOR3X1_18/C gnd NOR3X1_17/Y vdd NOR3X1
XFILL_37_1_1 gnd vdd FILL
XBUFX4_250 INVX8_5/Y gnd BUFX4_94/A vdd BUFX4
XBUFX4_272 INVX8_7/Y gnd BUFX4_60/A vdd BUFX4
XBUFX4_261 enable_i gnd BUFX4_261/Y vdd BUFX4
XFILL_0_INVX2_160 gnd vdd FILL
XFILL_0_INVX2_171 gnd vdd FILL
XBUFX4_283 INVX8_7/Y gnd BUFX4_82/A vdd BUFX4
XBUFX4_294 BUFX4_303/A gnd BUFX4_294/Y vdd BUFX4
XFILL_0_INVX2_193 gnd vdd FILL
XFILL_0_INVX2_182 gnd vdd FILL
XFILL_0_XNOR2X1_9 gnd vdd FILL
XOAI21X1_805 OAI21X1_805/A BUFX4_290/Y OAI21X1_805/C gnd OAI21X1_805/Y vdd OAI21X1
XOAI21X1_838 BUFX4_156/Y BUFX4_63/Y BUFX2_644/A gnd OAI21X1_840/C vdd OAI21X1
XOAI21X1_849 INVX1_50/Y BUFX4_265/Y OAI21X1_849/C gnd OAI21X1_849/Y vdd OAI21X1
XOAI21X1_827 XNOR2X1_55/A INVX4_25/Y INVX4_26/Y gnd OAI21X1_828/C vdd OAI21X1
XFILL_20_0_1 gnd vdd FILL
XOAI21X1_816 BUFX4_155/Y BUFX4_37/Y BUFX2_635/A gnd OAI21X1_818/C vdd OAI21X1
XFILL_21_16_1 gnd vdd FILL
XOAI21X1_1140 INVX1_187/A OR2X2_17/Y OAI21X1_1140/C gnd OAI21X1_1141/A vdd OAI21X1
XDFFPOSX1_741 BUFX2_379/A CLKBUF1_17/Y OAI21X1_1031/Y gnd vdd DFFPOSX1
XOAI21X1_1151 NOR2X1_147/Y AOI21X1_37/Y BUFX4_238/Y gnd OAI21X1_1152/C vdd OAI21X1
XOAI21X1_1173 XNOR2X1_73/Y BUFX4_203/Y NAND2X1_555/Y gnd OAI21X1_1173/Y vdd OAI21X1
XFILL_1_OAI21X1_1360 gnd vdd FILL
XDFFPOSX1_730 BUFX2_367/A CLKBUF1_56/Y OAI21X1_1009/Y gnd vdd DFFPOSX1
XOAI21X1_1162 NOR2X1_156/Y bundleAddress_i[25] BUFX4_239/Y gnd OAI21X1_1163/B vdd
+ OAI21X1
XFILL_1_OAI21X1_300 gnd vdd FILL
XDFFPOSX1_752 BUFX2_63/A CLKBUF1_12/Y OAI21X1_1044/Y gnd vdd DFFPOSX1
XDFFPOSX1_774 BUFX2_25/A CLKBUF1_14/Y OAI21X1_1066/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_950 gnd vdd FILL
XFILL_1_OAI21X1_1393 gnd vdd FILL
XFILL_1_DFFPOSX1_961 gnd vdd FILL
XFILL_1_OAI21X1_1382 gnd vdd FILL
XDFFPOSX1_763 BUFX2_12/A CLKBUF1_60/Y OAI21X1_1055/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_311 gnd vdd FILL
XFILL_1_OAI21X1_1371 gnd vdd FILL
XOAI21X1_1184 NOR3X1_14/C NAND2X1_571/Y INVX2_85/Y gnd NAND2X1_572/B vdd OAI21X1
XOAI21X1_1195 AOI21X1_43/Y OAI21X1_1195/B NAND2X1_579/Y gnd OAI21X1_1195/Y vdd OAI21X1
XFILL_0_OAI21X1_162 gnd vdd FILL
XFILL_0_OAI21X1_173 gnd vdd FILL
XFILL_0_OAI21X1_140 gnd vdd FILL
XFILL_1_OAI21X1_322 gnd vdd FILL
XFILL_1_DFFPOSX1_983 gnd vdd FILL
XFILL_1_DFFPOSX1_994 gnd vdd FILL
XFILL_0_OAI21X1_151 gnd vdd FILL
XFILL_1_DFFPOSX1_972 gnd vdd FILL
XDFFPOSX1_785 BUFX2_37/A CLKBUF1_53/Y OAI21X1_1077/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_333 gnd vdd FILL
XFILL_1_OAI21X1_344 gnd vdd FILL
XDFFPOSX1_796 BUFX2_49/A CLKBUF1_76/Y OAI21X1_1088/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_184 gnd vdd FILL
XFILL_0_OAI21X1_195 gnd vdd FILL
XFILL_1_OAI21X1_366 gnd vdd FILL
XFILL_1_OAI21X1_377 gnd vdd FILL
XFILL_1_OAI21X1_355 gnd vdd FILL
XFILL_1_OAI21X1_388 gnd vdd FILL
XFILL_1_CLKBUF1_9 gnd vdd FILL
XFILL_1_OAI21X1_399 gnd vdd FILL
XFILL_0_NAND3X1_26 gnd vdd FILL
XFILL_0_NAND3X1_15 gnd vdd FILL
XFILL_28_1_1 gnd vdd FILL
XFILL_0_NAND3X1_37 gnd vdd FILL
XFILL_0_NAND3X1_59 gnd vdd FILL
XFILL_0_NAND3X1_48 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XBUFX2_209 BUFX2_209/A gnd addr4_o[40] vdd BUFX2
XFILL_0_BUFX4_50 gnd vdd FILL
XFILL_0_BUFX4_72 gnd vdd FILL
XFILL_0_BUFX4_61 gnd vdd FILL
XFILL_0_BUFX4_94 gnd vdd FILL
XFILL_1_BUFX4_103 gnd vdd FILL
XFILL_0_BUFX4_83 gnd vdd FILL
XFILL_1_NAND2X1_361 gnd vdd FILL
XFILL_1_BUFX4_136 gnd vdd FILL
XFILL_1_NAND2X1_372 gnd vdd FILL
XFILL_1_BUFX4_125 gnd vdd FILL
XFILL_0_DFFPOSX1_551 gnd vdd FILL
XFILL_0_DFFPOSX1_540 gnd vdd FILL
XFILL_1_BUFX4_114 gnd vdd FILL
XFILL_0_NAND2X1_190 gnd vdd FILL
XFILL_26_15_1 gnd vdd FILL
XFILL_1_BUFX4_147 gnd vdd FILL
XFILL_0_DFFPOSX1_584 gnd vdd FILL
XFILL_0_DFFPOSX1_573 gnd vdd FILL
XFILL_1_BUFX4_169 gnd vdd FILL
XFILL_1_BUFX4_158 gnd vdd FILL
XFILL_0_DFFPOSX1_562 gnd vdd FILL
XFILL_0_DFFPOSX1_595 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XFILL_20_11_0 gnd vdd FILL
XFILL_0_OR2X2_20 gnd vdd FILL
XNAND3X1_50 AND2X2_24/B INVX1_198/Y AND2X2_24/A gnd NOR3X1_15/C vdd NAND3X1
XNAND3X1_61 INVX1_199/A INVX1_216/A NOR3X1_18/Y gnd INVX1_217/A vdd NAND3X1
XFILL_2_OAI21X1_1011 gnd vdd FILL
XBUFX2_710 BUFX2_710/A gnd pid2_o[24] vdd BUFX2
XBUFX2_721 BUFX2_721/A gnd pid3_o[15] vdd BUFX2
XFILL_19_1_1 gnd vdd FILL
XFILL_2_DFFPOSX1_601 gnd vdd FILL
XFILL_2_DFFPOSX1_612 gnd vdd FILL
XFILL_2_DFFPOSX1_623 gnd vdd FILL
XFILL_2_DFFPOSX1_645 gnd vdd FILL
XFILL_2_DFFPOSX1_634 gnd vdd FILL
XFILL_2_DFFPOSX1_656 gnd vdd FILL
XBUFX2_754 BUFX2_754/A gnd pid4_o[14] vdd BUFX2
XBUFX2_732 BUFX2_732/A gnd pid3_o[5] vdd BUFX2
XFILL_3_DFFPOSX1_70 gnd vdd FILL
XNOR2X1_72 OR2X2_6/B OR2X2_6/A gnd NOR2X1_72/Y vdd NOR2X1
XNOR2X1_50 NOR3X1_8/A INVX4_24/Y gnd NOR2X1_50/Y vdd NOR2X1
XNOR2X1_61 INVX4_5/Y OAI22X1_1/B gnd OAI22X1_1/C vdd NOR2X1
XFILL_2_OAI21X1_1088 gnd vdd FILL
XFILL_1_16_1 gnd vdd FILL
XBUFX2_743 BUFX2_743/A gnd pid3_o[23] vdd BUFX2
XBUFX2_776 BUFX2_776/A gnd pid4_o[22] vdd BUFX2
XBUFX2_787 BUFX2_787/A gnd tid1_o[45] vdd BUFX2
XBUFX2_765 BUFX2_765/A gnd pid4_o[4] vdd BUFX2
XFILL_3_DFFPOSX1_92 gnd vdd FILL
XFILL_3_DFFPOSX1_81 gnd vdd FILL
XNOR2X1_94 INVX2_51/Y NOR2X1_97/B gnd NOR2X1_94/Y vdd NOR2X1
XNOR2X1_83 NOR3X1_5/B NOR2X1_83/B gnd NOR2X1_83/Y vdd NOR2X1
XBUFX2_798 BUFX2_798/A gnd tid1_o[35] vdd BUFX2
XFILL_2_DFFPOSX1_678 gnd vdd FILL
XFILL_2_DFFPOSX1_667 gnd vdd FILL
XFILL_2_DFFPOSX1_689 gnd vdd FILL
XFILL_0_NOR2X1_127 gnd vdd FILL
XFILL_0_NOR2X1_116 gnd vdd FILL
XFILL_0_NOR2X1_105 gnd vdd FILL
XFILL_31_8_0 gnd vdd FILL
XFILL_0_NOR2X1_149 gnd vdd FILL
XFILL_0_NOR2X1_138 gnd vdd FILL
XFILL_25_10_0 gnd vdd FILL
XFILL_1_DFFPOSX1_202 gnd vdd FILL
XFILL_0_BUFX2_450 gnd vdd FILL
XFILL_1_DFFPOSX1_213 gnd vdd FILL
XFILL_1_DFFPOSX1_246 gnd vdd FILL
XFILL_1_DFFPOSX1_235 gnd vdd FILL
XFILL_0_BUFX2_472 gnd vdd FILL
XFILL_0_BUFX2_483 gnd vdd FILL
XFILL_0_BUFX2_461 gnd vdd FILL
XFILL_1_DFFPOSX1_224 gnd vdd FILL
XFILL_0_BUFX2_494 gnd vdd FILL
XFILL_1_DFFPOSX1_279 gnd vdd FILL
XFILL_1_DFFPOSX1_268 gnd vdd FILL
XNAND2X1_107 BUFX2_422/A BUFX4_373/Y gnd OAI21X1_363/C vdd NAND2X1
XFILL_1_DFFPOSX1_257 gnd vdd FILL
XNAND2X1_129 BUFX2_446/A BUFX4_356/Y gnd OAI21X1_385/C vdd NAND2X1
XNAND2X1_118 BUFX2_434/A BUFX4_358/Y gnd OAI21X1_374/C vdd NAND2X1
XNAND2X1_5 NAND2X1_5/A OAI21X1_5/A gnd OAI21X1_5/C vdd NAND2X1
XFILL_4_DFFPOSX1_728 gnd vdd FILL
XFILL_1_OAI21X1_16 gnd vdd FILL
XFILL_4_DFFPOSX1_706 gnd vdd FILL
XFILL_4_DFFPOSX1_717 gnd vdd FILL
XFILL_1_OAI21X1_38 gnd vdd FILL
XFILL_1_OAI21X1_27 gnd vdd FILL
XFILL_1_OAI21X1_49 gnd vdd FILL
XFILL_4_DFFPOSX1_739 gnd vdd FILL
XFILL_6_15_1 gnd vdd FILL
XNOR2X1_151 INVX4_38/Y INVX2_73/Y gnd AND2X2_28/A vdd NOR2X1
XNOR2X1_140 OR2X2_18/A NOR2X1_140/B gnd NOR2X1_140/Y vdd NOR2X1
XFILL_0_NAND2X1_70 gnd vdd FILL
XFILL_0_NAND2X1_81 gnd vdd FILL
XFILL_0_11_0 gnd vdd FILL
XFILL_0_NAND2X1_92 gnd vdd FILL
XNOR2X1_184 INVX2_105/Y NOR2X1_184/B gnd NOR2X1_184/Y vdd NOR2X1
XNOR2X1_162 INVX2_80/Y INVX4_43/Y gnd NOR2X1_162/Y vdd NOR2X1
XNOR2X1_173 INVX2_89/Y NOR3X1_15/C gnd NOR2X1_174/B vdd NOR2X1
XNOR2X1_195 bundleAddress_i[34] NOR2X1_195/B gnd NOR2X1_195/Y vdd NOR2X1
XFILL_22_8_0 gnd vdd FILL
XOAI21X1_613 NOR2X1_87/B INVX2_49/Y NOR2X1_96/B gnd OAI21X1_614/B vdd OAI21X1
XOAI21X1_624 BUFX4_102/Y BUFX4_367/Y BUFX2_565/A gnd OAI21X1_625/C vdd OAI21X1
XFILL_1_BUFX2_629 gnd vdd FILL
XOAI21X1_602 XNOR2X1_35/Y BUFX4_130/Y OAI21X1_602/C gnd OAI21X1_602/Y vdd OAI21X1
XOAI21X1_657 AOI21X1_26/Y OAI21X1_657/B OAI21X1_657/C gnd OAI21X1_657/Y vdd OAI21X1
XFILL_3_DFFPOSX1_318 gnd vdd FILL
XOAI21X1_646 OAI21X1_646/A AOI21X1_24/Y OAI21X1_646/C gnd OAI21X1_646/Y vdd OAI21X1
XFILL_3_DFFPOSX1_307 gnd vdd FILL
XOAI21X1_635 XNOR2X1_39/Y BUFX4_179/Y OAI21X1_635/C gnd OAI21X1_635/Y vdd OAI21X1
XFILL_3_DFFPOSX1_329 gnd vdd FILL
XOAI21X1_668 BUFX4_176/Y BUFX4_52/Y BUFX2_608/A gnd OAI21X1_669/C vdd OAI21X1
XOAI21X1_679 INVX1_34/Y INVX4_2/Y INVX2_13/Y gnd OAI21X1_679/Y vdd OAI21X1
XDFFPOSX1_582 BUFX2_613/A CLKBUF1_9/Y OAI21X1_757/Y gnd vdd DFFPOSX1
XDFFPOSX1_560 BUFX2_589/A CLKBUF1_90/Y OAI21X1_695/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1190 gnd vdd FILL
XDFFPOSX1_571 BUFX2_601/A CLKBUF1_44/Y OAI21X1_726/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_141 gnd vdd FILL
XFILL_1_DFFPOSX1_791 gnd vdd FILL
XXNOR2X1_18 XNOR2X1_18/A INVX4_18/Y gnd XNOR2X1_18/Y vdd XNOR2X1
XNAND2X1_630 NOR2X1_140/Y INVX4_51/A gnd NOR2X1_223/B vdd NAND2X1
XDFFPOSX1_593 BUFX2_625/A CLKBUF1_24/Y OAI21X1_789/Y gnd vdd DFFPOSX1
XFILL_1_INVX2_103 gnd vdd FILL
XFILL_1_OAI21X1_152 gnd vdd FILL
XFILL_1_OAI21X1_130 gnd vdd FILL
XXNOR2X1_29 MUX2X1_1/A INVX2_21/Y gnd XNOR2X1_29/Y vdd XNOR2X1
XFILL_1_DFFPOSX1_780 gnd vdd FILL
XFILL_1_OAI21X1_163 gnd vdd FILL
XNAND2X1_663 BUFX2_654/A BUFX4_363/Y gnd NAND2X1_663/Y vdd NAND2X1
XFILL_1_OAI21X1_185 gnd vdd FILL
XNAND2X1_652 BUFX2_661/A BUFX4_349/Y gnd NAND2X1_652/Y vdd NAND2X1
XNAND2X1_641 NAND2X1_641/A INVX1_225/A gnd NAND2X1_641/Y vdd NAND2X1
XFILL_2_OAI21X1_367 gnd vdd FILL
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XFILL_1_OAI21X1_174 gnd vdd FILL
XFILL_2_OAI21X1_356 gnd vdd FILL
XFILL_1_INVX2_158 gnd vdd FILL
XNAND2X1_696 BUFX2_687/A BUFX4_203/Y gnd NAND2X1_696/Y vdd NAND2X1
XINVX1_53 INVX1_53/A gnd INVX1_53/Y vdd INVX1
XFILL_2_OAI21X1_378 gnd vdd FILL
XFILL_1_OAI21X1_196 gnd vdd FILL
XINVX1_75 INVX1_75/A gnd INVX1_75/Y vdd INVX1
XINVX1_64 INVX1_64/A gnd INVX1_64/Y vdd INVX1
XNAND2X1_674 BUFX2_666/A OAI21X1_4/A gnd NAND2X1_674/Y vdd NAND2X1
XFILL_5_9_0 gnd vdd FILL
XFILL_5_10_0 gnd vdd FILL
XNAND2X1_685 BUFX2_704/A BUFX4_192/Y gnd NAND2X1_685/Y vdd NAND2X1
XINVX1_97 bundle_i[43] gnd INVX1_97/Y vdd INVX1
XINVX1_86 bundle_i[54] gnd INVX1_86/Y vdd INVX1
XBUFX2_17 BUFX2_17/A gnd addr1_o[40] vdd BUFX2
XBUFX2_28 BUFX2_28/A gnd addr1_o[30] vdd BUFX2
XBUFX2_39 BUFX2_39/A gnd addr1_o[20] vdd BUFX2
XDFFPOSX1_5 BUFX2_682/A CLKBUF1_65/Y DFFPOSX1_5/D gnd vdd DFFPOSX1
XFILL_13_8_0 gnd vdd FILL
XFILL_1_NAND2X1_191 gnd vdd FILL
XFILL_1_NAND2X1_180 gnd vdd FILL
XFILL_0_DFFPOSX1_392 gnd vdd FILL
XFILL_0_DFFPOSX1_381 gnd vdd FILL
XFILL_1_BUFX4_17 gnd vdd FILL
XFILL_0_DFFPOSX1_370 gnd vdd FILL
XFILL_1_BUFX4_39 gnd vdd FILL
XFILL_1_BUFX4_28 gnd vdd FILL
XFILL_3_DFFPOSX1_841 gnd vdd FILL
XFILL_3_DFFPOSX1_830 gnd vdd FILL
XFILL_3_DFFPOSX1_874 gnd vdd FILL
XFILL_3_DFFPOSX1_852 gnd vdd FILL
XFILL_3_DFFPOSX1_863 gnd vdd FILL
XFILL_0_OAI21X1_909 gnd vdd FILL
XFILL_3_DFFPOSX1_885 gnd vdd FILL
XFILL_3_DFFPOSX1_896 gnd vdd FILL
XNOR2X1_8 INVX4_5/Y INVX1_1/Y gnd NOR2X1_8/Y vdd NOR2X1
XFILL_11_16_0 gnd vdd FILL
XFILL_2_DFFPOSX1_431 gnd vdd FILL
XFILL_2_DFFPOSX1_420 gnd vdd FILL
XFILL_4_DFFPOSX1_60 gnd vdd FILL
XBUFX2_540 BUFX2_540/A gnd majID3_o[37] vdd BUFX2
XFILL_0_OAI21X1_1719 gnd vdd FILL
XBUFX2_551 BUFX2_551/A gnd majID3_o[27] vdd BUFX2
XBUFX2_562 BUFX2_562/A gnd majID3_o[17] vdd BUFX2
XFILL_2_DFFPOSX1_442 gnd vdd FILL
XFILL_2_DFFPOSX1_453 gnd vdd FILL
XFILL_2_DFFPOSX1_464 gnd vdd FILL
XFILL_0_OAI21X1_1708 gnd vdd FILL
XFILL_4_DFFPOSX1_82 gnd vdd FILL
XBUFX2_584 BUFX2_584/A gnd majID3_o[54] vdd BUFX2
XBUFX2_595 BUFX2_595/A gnd majID4_o[45] vdd BUFX2
XFILL_4_DFFPOSX1_93 gnd vdd FILL
XFILL_4_DFFPOSX1_71 gnd vdd FILL
XFILL_2_DFFPOSX1_486 gnd vdd FILL
XFILL_2_DFFPOSX1_497 gnd vdd FILL
XBUFX2_573 NOR2X1_96/A gnd majID3_o[7] vdd BUFX2
XFILL_2_DFFPOSX1_475 gnd vdd FILL
XFILL_5_DFFPOSX1_902 gnd vdd FILL
XFILL_5_DFFPOSX1_913 gnd vdd FILL
XFILL_5_DFFPOSX1_946 gnd vdd FILL
XFILL_5_DFFPOSX1_935 gnd vdd FILL
XFILL_5_DFFPOSX1_924 gnd vdd FILL
XFILL_5_DFFPOSX1_968 gnd vdd FILL
XFILL_5_DFFPOSX1_979 gnd vdd FILL
XFILL_5_DFFPOSX1_957 gnd vdd FILL
XAOI21X1_18 AOI21X1_18/A OR2X2_11/Y NOR2X1_89/Y gnd AOI21X1_18/Y vdd AOI21X1
XAOI21X1_29 INVX4_1/Y INVX2_8/Y NOR2X1_3/B gnd INVX2_52/A vdd AOI21X1
XFILL_0_BUFX2_291 gnd vdd FILL
XFILL_0_BUFX2_280 gnd vdd FILL
XFILL_0_AND2X2_4 gnd vdd FILL
XFILL_4_DFFPOSX1_503 gnd vdd FILL
XFILL_4_DFFPOSX1_525 gnd vdd FILL
XFILL_4_DFFPOSX1_536 gnd vdd FILL
XFILL_4_DFFPOSX1_514 gnd vdd FILL
XFILL_16_15_0 gnd vdd FILL
XFILL_4_DFFPOSX1_547 gnd vdd FILL
XFILL_4_DFFPOSX1_569 gnd vdd FILL
XFILL_4_DFFPOSX1_558 gnd vdd FILL
XFILL_1_BUFX2_1016 gnd vdd FILL
XFILL_1_BUFX2_1027 gnd vdd FILL
XFILL_1_BUFX2_426 gnd vdd FILL
XFILL_1_BUFX2_448 gnd vdd FILL
XFILL_1_BUFX2_437 gnd vdd FILL
XOAI21X1_421 XNOR2X1_4/Y BUFX4_215/Y OAI21X1_421/C gnd OAI21X1_421/Y vdd OAI21X1
XOAI21X1_432 XNOR2X1_7/Y BUFX4_236/Y OAI21X1_432/C gnd OAI21X1_432/Y vdd OAI21X1
XOAI21X1_410 AND2X2_1/Y bundleStartMajId_i[55] BUFX4_244/Y gnd OAI21X1_411/A vdd OAI21X1
XFILL_3_DFFPOSX1_104 gnd vdd FILL
XFILL_3_DFFPOSX1_126 gnd vdd FILL
XFILL_3_DFFPOSX1_115 gnd vdd FILL
XFILL_3_DFFPOSX1_137 gnd vdd FILL
XFILL_1_CLKBUF1_17 gnd vdd FILL
XOAI21X1_454 XNOR2X1_15/Y BUFX4_224/Y OAI21X1_454/C gnd OAI21X1_454/Y vdd OAI21X1
XOAI21X1_465 NOR3X1_2/C NOR3X1_2/B NOR3X1_2/A gnd OAI21X1_465/Y vdd OAI21X1
XOAI21X1_443 OAI21X1_443/A BUFX4_214/Y OAI21X1_443/C gnd OAI21X1_443/Y vdd OAI21X1
XFILL_1_CLKBUF1_28 gnd vdd FILL
XFILL_1_CLKBUF1_39 gnd vdd FILL
XFILL_3_DFFPOSX1_148 gnd vdd FILL
XOAI21X1_498 OAI21X1_498/A AOI21X1_6/Y OAI21X1_498/C gnd OAI21X1_498/Y vdd OAI21X1
XOAI21X1_476 OAI21X1_476/A INVX2_33/Y BUFX4_241/Y gnd OAI21X1_477/A vdd OAI21X1
XOAI21X1_487 INVX1_22/Y OAI21X1_487/B OAI21X1_487/C gnd OAI21X1_487/Y vdd OAI21X1
XFILL_3_DFFPOSX1_159 gnd vdd FILL
XDFFPOSX1_390 BUFX2_421/A CLKBUF1_44/Y OAI21X1_362/Y gnd vdd DFFPOSX1
XFILL_2_OAI21X1_142 gnd vdd FILL
XFILL_8_0_1 gnd vdd FILL
XNAND2X1_471 BUFX2_99/A BUFX4_216/Y gnd NAND2X1_471/Y vdd NAND2X1
XFILL_34_16_0 gnd vdd FILL
XNAND2X1_460 BUFX2_55/A BUFX4_330/Y gnd NAND2X1_460/Y vdd NAND2X1
XFILL_2_OAI21X1_175 gnd vdd FILL
XNAND2X1_493 BUFX2_71/A BUFX4_235/Y gnd NAND2X1_493/Y vdd NAND2X1
XNAND2X1_482 bundleAddress_i[55] bundleAddress_i[54] gnd NOR2X1_127/B vdd NAND2X1
XFILL_0_INVX1_203 gnd vdd FILL
XFILL_0_INVX1_225 gnd vdd FILL
XFILL_0_INVX1_214 gnd vdd FILL
XFILL_5_DFFPOSX1_209 gnd vdd FILL
XFILL_0_OAI21X1_24 gnd vdd FILL
XFILL_0_OAI21X1_13 gnd vdd FILL
XFILL_0_OAI21X1_35 gnd vdd FILL
XFILL_0_OAI21X1_46 gnd vdd FILL
XFILL_0_OAI21X1_57 gnd vdd FILL
XOAI21X1_1706 BUFX4_7/Y BUFX4_388/Y BUFX2_737/A gnd OAI21X1_1707/C vdd OAI21X1
XFILL_1_BUFX2_960 gnd vdd FILL
XFILL_1_BUFX2_993 gnd vdd FILL
XOAI21X1_1739 INVX2_131/Y BUFX4_301/Y OAI21X1_1739/C gnd DFFPOSX1_82/D vdd OAI21X1
XOAI21X1_1728 BUFX4_178/Y BUFX4_55/Y BUFX2_776/A gnd OAI21X1_1729/C vdd OAI21X1
XOAI21X1_1717 INVX2_120/Y INVX8_2/A OAI21X1_1717/C gnd DFFPOSX1_71/D vdd OAI21X1
XFILL_0_OAI21X1_79 gnd vdd FILL
XFILL_0_OAI21X1_68 gnd vdd FILL
XFILL_3_DFFPOSX1_660 gnd vdd FILL
XFILL_3_DFFPOSX1_671 gnd vdd FILL
XFILL_3_DFFPOSX1_682 gnd vdd FILL
XFILL_0_OAI21X1_717 gnd vdd FILL
XFILL_0_OAI21X1_728 gnd vdd FILL
XFILL_0_OAI21X1_739 gnd vdd FILL
XFILL_0_OAI21X1_706 gnd vdd FILL
XFILL_3_DFFPOSX1_693 gnd vdd FILL
XFILL_0_NAND2X1_701 gnd vdd FILL
XFILL_0_NAND2X1_734 gnd vdd FILL
XFILL_36_7_0 gnd vdd FILL
XFILL_0_NAND2X1_745 gnd vdd FILL
XFILL_0_OAI21X1_1516 gnd vdd FILL
XFILL_0_NAND2X1_712 gnd vdd FILL
XFILL_0_NAND2X1_723 gnd vdd FILL
XFILL_0_OAI21X1_1505 gnd vdd FILL
XFILL_2_DFFPOSX1_261 gnd vdd FILL
XBUFX2_381 BUFX2_381/A gnd instr4_o[1] vdd BUFX2
XFILL_2_DFFPOSX1_272 gnd vdd FILL
XFILL_0_OAI21X1_1527 gnd vdd FILL
XFILL_2_DFFPOSX1_250 gnd vdd FILL
XFILL_2_DFFPOSX1_283 gnd vdd FILL
XFILL_0_OAI21X1_1538 gnd vdd FILL
XBUFX2_370 BUFX2_370/A gnd instr4_o[11] vdd BUFX2
XFILL_0_NAND2X1_767 gnd vdd FILL
XFILL_0_NAND2X1_756 gnd vdd FILL
XFILL_0_OAI21X1_1549 gnd vdd FILL
XFILL_5_DFFPOSX1_50 gnd vdd FILL
XFILL_5_DFFPOSX1_61 gnd vdd FILL
XFILL_5_DFFPOSX1_72 gnd vdd FILL
XFILL_2_DFFPOSX1_294 gnd vdd FILL
XBUFX2_392 BUFX2_392/A gnd is64b4_o vdd BUFX2
XFILL_5_DFFPOSX1_710 gnd vdd FILL
XFILL_5_DFFPOSX1_94 gnd vdd FILL
XFILL_5_DFFPOSX1_83 gnd vdd FILL
XFILL_5_DFFPOSX1_721 gnd vdd FILL
XOAI21X1_81 BUFX4_132/Y INVX2_150/Y OAI21X1_81/C gnd OAI21X1_81/Y vdd OAI21X1
XFILL_5_DFFPOSX1_754 gnd vdd FILL
XFILL_5_DFFPOSX1_743 gnd vdd FILL
XOAI21X1_70 INVX2_6/Y BUFX4_217/Y OAI21X1_70/C gnd OAI21X1_70/Y vdd OAI21X1
XFILL_5_DFFPOSX1_732 gnd vdd FILL
XFILL_5_DFFPOSX1_776 gnd vdd FILL
XFILL_5_DFFPOSX1_787 gnd vdd FILL
XOAI21X1_92 BUFX4_6/A BUFX4_324/Y BUFX2_907/A gnd OAI21X1_93/C vdd OAI21X1
XFILL_5_DFFPOSX1_798 gnd vdd FILL
XFILL_5_DFFPOSX1_765 gnd vdd FILL
XFILL_4_DFFPOSX1_311 gnd vdd FILL
XFILL_4_DFFPOSX1_300 gnd vdd FILL
XFILL_4_DFFPOSX1_322 gnd vdd FILL
XFILL_4_DFFPOSX1_333 gnd vdd FILL
XFILL_4_DFFPOSX1_344 gnd vdd FILL
XFILL_2_DFFPOSX1_1014 gnd vdd FILL
XFILL_0_DFFPOSX1_90 gnd vdd FILL
XFILL_2_DFFPOSX1_1003 gnd vdd FILL
XFILL_4_DFFPOSX1_388 gnd vdd FILL
XFILL_4_DFFPOSX1_377 gnd vdd FILL
XFILL_4_DFFPOSX1_366 gnd vdd FILL
XFILL_4_DFFPOSX1_355 gnd vdd FILL
XFILL_2_DFFPOSX1_1025 gnd vdd FILL
XFILL_27_7_0 gnd vdd FILL
XFILL_4_DFFPOSX1_399 gnd vdd FILL
XFILL_2_7_0 gnd vdd FILL
XFILL_1_BUFX2_201 gnd vdd FILL
XFILL_1_BUFX2_234 gnd vdd FILL
XFILL_1_BUFX2_245 gnd vdd FILL
XFILL_1_BUFX2_223 gnd vdd FILL
XFILL_1_BUFX2_278 gnd vdd FILL
XOAI21X1_240 BUFX4_156/Y BUFX4_62/Y BUFX2_982/A gnd OAI21X1_241/C vdd OAI21X1
XFILL_10_6_0 gnd vdd FILL
XOAI21X1_273 INVX2_182/Y BUFX4_292/Y OAI21X1_273/C gnd OAI21X1_273/Y vdd OAI21X1
XOAI21X1_262 BUFX4_151/Y BUFX4_75/Y BUFX2_994/A gnd OAI21X1_263/C vdd OAI21X1
XOAI21X1_251 INVX2_171/Y BUFX4_292/Y OAI21X1_251/C gnd OAI21X1_251/Y vdd OAI21X1
XFILL_23_13_1 gnd vdd FILL
XFILL_1_BUFX2_289 gnd vdd FILL
XOAI21X1_295 INVX2_193/Y BUFX4_292/Y OAI21X1_295/C gnd OAI21X1_295/Y vdd OAI21X1
XOAI21X1_284 BUFX4_133/Y BUFX4_31/Y BUFX2_1006/A gnd OAI21X1_285/C vdd OAI21X1
XFILL_6_DFFPOSX1_416 gnd vdd FILL
XFILL_6_DFFPOSX1_427 gnd vdd FILL
XFILL_6_DFFPOSX1_449 gnd vdd FILL
XFILL_6_DFFPOSX1_438 gnd vdd FILL
XNAND2X1_290 bundleStartMajId_i[28] bundleStartMajId_i[27] gnd NOR2X1_77/B vdd NAND2X1
XFILL_18_7_0 gnd vdd FILL
XFILL_1_NAND3X1_8 gnd vdd FILL
XFILL_0_INVX8_3 gnd vdd FILL
XFILL_28_12_1 gnd vdd FILL
XFILL_5_DFFPOSX1_1007 gnd vdd FILL
XFILL_5_DFFPOSX1_1018 gnd vdd FILL
XFILL_5_DFFPOSX1_1029 gnd vdd FILL
XDFFPOSX1_18 BUFX2_687/A CLKBUF1_86/Y DFFPOSX1_18/D gnd vdd DFFPOSX1
XFILL_0_BUFX4_342 gnd vdd FILL
XOAI21X1_1514 XNOR2X1_102/Y BUFX4_297/Y OAI21X1_1514/C gnd OAI21X1_1514/Y vdd OAI21X1
XFILL_0_BUFX4_331 gnd vdd FILL
XFILL_1_BUFX2_790 gnd vdd FILL
XFILL_0_BUFX4_320 gnd vdd FILL
XOAI21X1_1503 NOR3X1_16/B NAND3X1_65/Y OAI21X1_1503/C gnd OAI21X1_1505/A vdd OAI21X1
XFILL_1_OAI21X1_1712 gnd vdd FILL
XFILL_0_BUFX4_353 gnd vdd FILL
XFILL_1_OAI21X1_1701 gnd vdd FILL
XFILL_0_BUFX4_375 gnd vdd FILL
XOAI21X1_1525 BUFX4_128/Y BUFX4_39/Y BUFX2_235/A gnd OAI21X1_1527/C vdd OAI21X1
XDFFPOSX1_29 BUFX2_699/A CLKBUF1_47/Y DFFPOSX1_29/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1734 gnd vdd FILL
XOAI21X1_1536 OR2X2_21/A INVX4_44/Y INVX2_84/Y gnd OAI21X1_1537/C vdd OAI21X1
XOAI21X1_1547 OR2X2_21/A INVX4_48/Y INVX2_87/Y gnd NAND2X1_644/A vdd OAI21X1
XFILL_0_BUFX4_364 gnd vdd FILL
XFILL_1_OAI21X1_1723 gnd vdd FILL
XFILL_1_OAI21X1_1756 gnd vdd FILL
XFILL_0_BUFX4_386 gnd vdd FILL
XFILL_1_OAI21X1_1745 gnd vdd FILL
XFILL_1_OAI21X1_1767 gnd vdd FILL
XOAI21X1_1569 AOI21X1_66/Y OAI21X1_1569/B OAI21X1_1569/C gnd OAI21X1_1569/Y vdd OAI21X1
XOAI21X1_1558 OR2X2_21/A OR2X2_21/B INVX2_89/Y gnd NAND2X1_646/A vdd OAI21X1
XFILL_0_OAI21X1_503 gnd vdd FILL
XFILL_3_DFFPOSX1_490 gnd vdd FILL
XFILL_1_OAI21X1_1778 gnd vdd FILL
XFILL_1_OAI21X1_1789 gnd vdd FILL
XFILL_0_BUFX2_1013 gnd vdd FILL
XFILL_0_BUFX2_1002 gnd vdd FILL
XFILL_0_OAI21X1_525 gnd vdd FILL
XFILL_1_OAI21X1_718 gnd vdd FILL
XFILL_1_OAI21X1_707 gnd vdd FILL
XFILL_0_OAI21X1_547 gnd vdd FILL
XFILL_0_OAI21X1_536 gnd vdd FILL
XFILL_0_OAI21X1_514 gnd vdd FILL
XFILL_0_BUFX2_1024 gnd vdd FILL
XFILL_0_OAI21X1_569 gnd vdd FILL
XFILL_0_OAI21X1_558 gnd vdd FILL
XFILL_1_OAI21X1_729 gnd vdd FILL
XFILL_0_CLKBUF1_25 gnd vdd FILL
XFILL_0_CLKBUF1_14 gnd vdd FILL
XFILL_0_CLKBUF1_36 gnd vdd FILL
XFILL_0_CLKBUF1_47 gnd vdd FILL
XFILL_0_NAND2X1_520 gnd vdd FILL
XFILL_0_CLKBUF1_69 gnd vdd FILL
XFILL_3_13_1 gnd vdd FILL
XFILL_0_CLKBUF1_58 gnd vdd FILL
XFILL_0_NAND2X1_531 gnd vdd FILL
XFILL_0_OAI21X1_1302 gnd vdd FILL
XFILL_1_NAND2X1_702 gnd vdd FILL
XFILL_1_NAND2X1_724 gnd vdd FILL
XFILL_0_NAND2X1_553 gnd vdd FILL
XFILL_0_OAI21X1_1324 gnd vdd FILL
XFILL_0_OAI21X1_1313 gnd vdd FILL
XFILL_0_NAND2X1_542 gnd vdd FILL
XFILL_0_DFFPOSX1_903 gnd vdd FILL
XFILL_0_OAI21X1_1335 gnd vdd FILL
XFILL_0_NAND2X1_564 gnd vdd FILL
XFILL_0_NAND2X1_586 gnd vdd FILL
XFILL_0_DFFPOSX1_914 gnd vdd FILL
XFILL_0_OAI21X1_1346 gnd vdd FILL
XFILL_0_DFFPOSX1_925 gnd vdd FILL
XFILL_0_OAI21X1_1357 gnd vdd FILL
XFILL_0_NAND2X1_575 gnd vdd FILL
XFILL_1_NAND2X1_735 gnd vdd FILL
XFILL_1_NAND2X1_757 gnd vdd FILL
XFILL_1_NAND2X1_768 gnd vdd FILL
XFILL_0_DFFPOSX1_936 gnd vdd FILL
XFILL_0_NAND2X1_597 gnd vdd FILL
XFILL_0_DFFPOSX1_947 gnd vdd FILL
XFILL_0_OAI21X1_1379 gnd vdd FILL
XFILL_0_OAI21X1_1368 gnd vdd FILL
XFILL_0_DFFPOSX1_958 gnd vdd FILL
XFILL_0_DFFPOSX1_969 gnd vdd FILL
XFILL_5_DFFPOSX1_551 gnd vdd FILL
XFILL_5_DFFPOSX1_540 gnd vdd FILL
XFILL_5_DFFPOSX1_562 gnd vdd FILL
XFILL_5_DFFPOSX1_595 gnd vdd FILL
XFILL_5_DFFPOSX1_584 gnd vdd FILL
XFILL_5_DFFPOSX1_573 gnd vdd FILL
XFILL_0_OR2X2_8 gnd vdd FILL
XFILL_1_BUFX4_6 gnd vdd FILL
XFILL_1_AOI21X1_2 gnd vdd FILL
XFILL_8_12_1 gnd vdd FILL
XCLKBUF1_60 BUFX4_86/Y gnd CLKBUF1_60/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_130 gnd vdd FILL
XCLKBUF1_93 BUFX4_86/Y gnd CLKBUF1_93/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_163 gnd vdd FILL
XFILL_4_DFFPOSX1_152 gnd vdd FILL
XCLKBUF1_82 BUFX4_89/Y gnd CLKBUF1_82/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_141 gnd vdd FILL
XCLKBUF1_71 BUFX4_89/Y gnd CLKBUF1_71/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_91 gnd vdd FILL
XFILL_4_DFFPOSX1_185 gnd vdd FILL
XFILL_1_DFFPOSX1_80 gnd vdd FILL
XFILL_2_NOR3X1_18 gnd vdd FILL
XFILL_4_DFFPOSX1_196 gnd vdd FILL
XFILL_4_DFFPOSX1_174 gnd vdd FILL
XFILL_1_NAND3X1_19 gnd vdd FILL
XINVX1_101 bundle_i[39] gnd INVX1_101/Y vdd INVX1
XFILL_0_BUFX2_802 gnd vdd FILL
XFILL_0_BUFX2_824 gnd vdd FILL
XFILL_1_OAI21X1_1019 gnd vdd FILL
XFILL_0_BUFX2_813 gnd vdd FILL
XFILL_1_INVX4_6 gnd vdd FILL
XFILL_1_OAI21X1_1008 gnd vdd FILL
XINVX1_112 bundle_i[92] gnd INVX1_112/Y vdd INVX1
XINVX1_123 bundle_i[81] gnd INVX1_123/Y vdd INVX1
XFILL_0_BUFX2_857 gnd vdd FILL
XFILL_1_DFFPOSX1_609 gnd vdd FILL
XFILL_0_BUFX2_846 gnd vdd FILL
XINVX1_134 bundle_i[70] gnd INVX1_134/Y vdd INVX1
XFILL_0_BUFX2_835 gnd vdd FILL
XFILL_0_BUFX2_868 gnd vdd FILL
XFILL_0_BUFX2_879 gnd vdd FILL
XINVX1_145 bundle_i[123] gnd INVX1_145/Y vdd INVX1
XINVX1_156 bundle_i[112] gnd INVX1_156/Y vdd INVX1
XINVX1_167 bundle_i[101] gnd INVX1_167/Y vdd INVX1
XFILL_6_DFFPOSX1_202 gnd vdd FILL
XFILL_6_DFFPOSX1_213 gnd vdd FILL
XINVX1_189 INVX1_189/A gnd INVX1_189/Y vdd INVX1
XINVX1_178 bundleAddress_i[17] gnd INVX1_178/Y vdd INVX1
XFILL_6_DFFPOSX1_224 gnd vdd FILL
XFILL_0_INVX2_11 gnd vdd FILL
XFILL_0_INVX2_33 gnd vdd FILL
XFILL_0_INVX2_55 gnd vdd FILL
XFILL_0_INVX2_44 gnd vdd FILL
XFILL_14_18_1 gnd vdd FILL
XFILL_0_INVX2_22 gnd vdd FILL
XFILL_0_INVX2_66 gnd vdd FILL
XFILL_0_INVX2_88 gnd vdd FILL
XFILL_0_INVX2_77 gnd vdd FILL
XFILL_0_INVX2_99 gnd vdd FILL
XFILL_0_CLKBUF1_1 gnd vdd FILL
XFILL_1_NOR3X1_8 gnd vdd FILL
XFILL_34_3 gnd vdd FILL
XFILL_33_5_0 gnd vdd FILL
XFILL_27_2 gnd vdd FILL
XFILL_0_BUFX4_150 gnd vdd FILL
XOAI21X1_1300 AND2X2_30/A INVX2_75/Y INVX4_40/Y gnd OAI21X1_1301/C vdd OAI21X1
XOAI21X1_1311 XNOR2X1_83/Y BUFX4_157/Y OAI21X1_1311/C gnd OAI21X1_1311/Y vdd OAI21X1
XOAI21X1_1322 OAI21X1_1322/A AOI21X1_50/Y OAI21X1_1322/C gnd OAI21X1_1322/Y vdd OAI21X1
XFILL_0_BUFX4_172 gnd vdd FILL
XFILL_0_BUFX4_161 gnd vdd FILL
XFILL_1_OAI21X1_1520 gnd vdd FILL
XOAI21X1_1333 BUFX4_105/Y BUFX4_360/Y BUFX2_170/A gnd OAI21X1_1335/C vdd OAI21X1
XFILL_0_BUFX4_183 gnd vdd FILL
XFILL_1_OAI21X1_1531 gnd vdd FILL
XDFFPOSX1_901 BUFX2_151/A CLKBUF1_35/Y OAI21X1_1290/Y gnd vdd DFFPOSX1
XOAI21X1_1344 NOR2X1_206/Y OAI21X1_1344/B OAI21X1_1344/C gnd OAI21X1_1344/Y vdd OAI21X1
XFILL_1_OAI21X1_1542 gnd vdd FILL
XDFFPOSX1_923 BUFX2_176/A CLKBUF1_38/Y OAI21X1_1349/Y gnd vdd DFFPOSX1
XFILL_0_BUFX4_194 gnd vdd FILL
XDFFPOSX1_912 BUFX2_164/A CLKBUF1_53/Y OAI21X1_1319/Y gnd vdd DFFPOSX1
XOAI21X1_1355 BUFX4_1/A BUFX4_364/Y BUFX2_179/A gnd OAI21X1_1357/C vdd OAI21X1
XFILL_0_OAI21X1_300 gnd vdd FILL
XOAI21X1_1399 OAI21X1_1399/A BUFX4_290/Y OAI21X1_1399/C gnd OAI21X1_1399/Y vdd OAI21X1
XFILL_1_OAI21X1_1575 gnd vdd FILL
XOAI21X1_1388 BUFX4_179/Y BUFX4_42/Y BUFX2_205/A gnd OAI21X1_1389/C vdd OAI21X1
XFILL_0_OAI21X1_322 gnd vdd FILL
XDFFPOSX1_945 BUFX2_256/A CLKBUF1_91/Y OAI21X1_1412/Y gnd vdd DFFPOSX1
XDFFPOSX1_934 BUFX2_188/A CLKBUF1_30/Y OAI21X1_1381/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1564 gnd vdd FILL
XFILL_0_OAI21X1_311 gnd vdd FILL
XOAI21X1_1377 INVX1_217/A INVX2_91/Y BUFX4_308/Y gnd OAI21X1_1378/B vdd OAI21X1
XOAI21X1_1366 INVX1_215/A INVX1_197/A BUFX4_308/Y gnd OAI21X1_1367/B vdd OAI21X1
XDFFPOSX1_956 BUFX2_206/A CLKBUF1_83/Y OAI21X1_1445/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1553 gnd vdd FILL
XFILL_1_BUFX2_50 gnd vdd FILL
XFILL_1_OAI21X1_1597 gnd vdd FILL
XFILL_1_BUFX2_83 gnd vdd FILL
XDFFPOSX1_967 BUFX2_218/A CLKBUF1_21/Y OAI21X1_1475/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_526 gnd vdd FILL
XDFFPOSX1_978 BUFX2_230/A CLKBUF1_85/Y OAI21X1_1512/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_504 gnd vdd FILL
XFILL_1_OAI21X1_515 gnd vdd FILL
XDFFPOSX1_989 BUFX2_242/A CLKBUF1_28/Y OAI21X1_1546/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_355 gnd vdd FILL
XFILL_1_BUFX2_94 gnd vdd FILL
XFILL_1_OAI21X1_1586 gnd vdd FILL
XFILL_0_OAI21X1_333 gnd vdd FILL
XFILL_0_OAI21X1_344 gnd vdd FILL
XFILL_0_OAI21X1_366 gnd vdd FILL
XFILL_0_OAI21X1_388 gnd vdd FILL
XFILL_0_OAI21X1_377 gnd vdd FILL
XFILL_19_17_1 gnd vdd FILL
XFILL_1_OAI21X1_559 gnd vdd FILL
XFILL_1_OAI21X1_548 gnd vdd FILL
XFILL_1_OAI21X1_537 gnd vdd FILL
XFILL_0_OAI21X1_399 gnd vdd FILL
XFILL_6_DFFPOSX1_780 gnd vdd FILL
XFILL_6_DFFPOSX1_791 gnd vdd FILL
XFILL_1_OAI21X1_5 gnd vdd FILL
XFILL_13_13_0 gnd vdd FILL
XFILL_0_DFFPOSX1_700 gnd vdd FILL
XFILL_0_NAND2X1_361 gnd vdd FILL
XFILL_0_OAI21X1_1110 gnd vdd FILL
XFILL_1_NAND2X1_532 gnd vdd FILL
XFILL_0_OAI21X1_1121 gnd vdd FILL
XFILL_0_OAI21X1_1132 gnd vdd FILL
XFILL_0_NAND2X1_350 gnd vdd FILL
XFILL_0_NAND2X1_394 gnd vdd FILL
XFILL_0_NAND2X1_383 gnd vdd FILL
XFILL_0_DFFPOSX1_711 gnd vdd FILL
XFILL_0_OAI21X1_1143 gnd vdd FILL
XFILL_0_DFFPOSX1_722 gnd vdd FILL
XFILL_0_OAI21X1_1154 gnd vdd FILL
XFILL_0_NAND2X1_372 gnd vdd FILL
XFILL_1_BUFX4_318 gnd vdd FILL
XFILL_24_5_0 gnd vdd FILL
XFILL_1_BUFX4_307 gnd vdd FILL
XFILL_1_NAND2X1_565 gnd vdd FILL
XFILL_0_DFFPOSX1_733 gnd vdd FILL
XFILL_0_OAI21X1_1165 gnd vdd FILL
XFILL_0_DFFPOSX1_755 gnd vdd FILL
XFILL_0_DFFPOSX1_744 gnd vdd FILL
XFILL_1_BUFX4_329 gnd vdd FILL
XFILL_0_OAI21X1_1176 gnd vdd FILL
XFILL_1_NAND2X1_598 gnd vdd FILL
XFILL_1_NAND2X1_587 gnd vdd FILL
XFILL_0_OAI21X1_1198 gnd vdd FILL
XFILL_0_OAI21X1_1187 gnd vdd FILL
XFILL_0_DFFPOSX1_766 gnd vdd FILL
XFILL_0_DFFPOSX1_788 gnd vdd FILL
XFILL_0_DFFPOSX1_777 gnd vdd FILL
XFILL_0_DFFPOSX1_799 gnd vdd FILL
XFILL_5_DFFPOSX1_381 gnd vdd FILL
XFILL_5_DFFPOSX1_370 gnd vdd FILL
XFILL_5_DFFPOSX1_392 gnd vdd FILL
XFILL_0_BUFX2_109 gnd vdd FILL
XFILL_1_NAND2X1_30 gnd vdd FILL
XINVX4_20 bundleStartMajId_i[22] gnd INVX4_20/Y vdd INVX4
XFILL_1_NAND2X1_52 gnd vdd FILL
XINVX4_31 INVX4_31/A gnd INVX4_31/Y vdd INVX4
XFILL_1_NAND2X1_74 gnd vdd FILL
XINVX4_42 bundleAddress_i[22] gnd INVX4_42/Y vdd INVX4
XFILL_37_18_1 gnd vdd FILL
XFILL_1_BUFX2_3 gnd vdd FILL
XFILL_18_12_0 gnd vdd FILL
XFILL_7_6_0 gnd vdd FILL
XFILL_31_14_0 gnd vdd FILL
XFILL_2_DFFPOSX1_805 gnd vdd FILL
XBUFX2_903 BUFX2_903/A gnd tid2_o[55] vdd BUFX2
XBUFX2_914 BUFX2_914/A gnd tid3_o[46] vdd BUFX2
XBUFX2_947 BUFX2_947/A gnd tid3_o[16] vdd BUFX2
XBUFX2_925 BUFX2_925/A gnd tid3_o[36] vdd BUFX2
XBUFX2_936 BUFX2_936/A gnd tid3_o[26] vdd BUFX2
XFILL_2_DFFPOSX1_816 gnd vdd FILL
XFILL_2_DFFPOSX1_70 gnd vdd FILL
XFILL_2_DFFPOSX1_838 gnd vdd FILL
XFILL_2_DFFPOSX1_81 gnd vdd FILL
XFILL_2_DFFPOSX1_827 gnd vdd FILL
XBUFX2_958 BUFX2_958/A gnd tid3_o[6] vdd BUFX2
XBUFX2_969 BUFX2_969/A gnd tid4_o[63] vdd BUFX2
XFILL_2_DFFPOSX1_92 gnd vdd FILL
XFILL_2_DFFPOSX1_849 gnd vdd FILL
XFILL_15_5_0 gnd vdd FILL
XDFFPOSX1_208 BUFX2_880/A CLKBUF1_3/Y OAI21X1_52/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_632 gnd vdd FILL
XDFFPOSX1_219 BUFX2_892/A CLKBUF1_87/Y OAI21X1_63/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_621 gnd vdd FILL
XFILL_0_BUFX2_610 gnd vdd FILL
XFILL_0_BUFX2_665 gnd vdd FILL
XFILL_0_BUFX2_654 gnd vdd FILL
XFILL_0_BUFX2_643 gnd vdd FILL
XFILL_1_DFFPOSX1_406 gnd vdd FILL
XFILL_1_DFFPOSX1_439 gnd vdd FILL
XFILL_1_DFFPOSX1_428 gnd vdd FILL
XFILL_0_BUFX2_676 gnd vdd FILL
XFILL_1_DFFPOSX1_417 gnd vdd FILL
XFILL_0_BUFX2_687 gnd vdd FILL
XFILL_0_BUFX2_698 gnd vdd FILL
XFILL_36_13_0 gnd vdd FILL
XNOR3X1_18 NOR3X1_18/A NOR3X1_18/B NOR3X1_18/C gnd NOR3X1_18/Y vdd NOR3X1
XBUFX4_240 INVX8_1/Y gnd BUFX4_240/Y vdd BUFX4
XBUFX4_251 INVX8_5/Y gnd BUFX4_251/Y vdd BUFX4
XBUFX4_273 INVX8_7/Y gnd BUFX4_55/A vdd BUFX4
XBUFX4_262 enable_i gnd BUFX4_262/Y vdd BUFX4
XFILL_0_INVX2_150 gnd vdd FILL
XFILL_0_INVX2_161 gnd vdd FILL
XBUFX4_295 BUFX4_303/A gnd BUFX4_295/Y vdd BUFX4
XBUFX4_284 INVX8_2/Y gnd BUFX4_284/Y vdd BUFX4
XFILL_0_INVX2_172 gnd vdd FILL
XFILL_0_INVX2_194 gnd vdd FILL
XFILL_0_INVX2_183 gnd vdd FILL
XOAI21X1_806 NOR3X1_8/C INVX2_45/A INVX2_34/Y gnd OAI21X1_807/C vdd OAI21X1
XOAI21X1_839 OAI21X1_839/A INVX4_28/Y BUFX4_288/Y gnd OAI21X1_840/B vdd OAI21X1
XOAI21X1_828 INVX1_43/Y XNOR2X1_55/A OAI21X1_828/C gnd OAI21X1_830/A vdd OAI21X1
XOAI21X1_817 NAND3X1_33/Y INVX2_46/Y BUFX4_285/Y gnd OAI21X1_818/A vdd OAI21X1
XOAI21X1_1130 XNOR2X1_58/Y OAI21X1_8/B NAND2X1_498/Y gnd OAI21X1_1130/Y vdd OAI21X1
XOAI21X1_1152 INVX1_191/Y BUFX4_238/Y OAI21X1_1152/C gnd OAI21X1_1152/Y vdd OAI21X1
XOAI21X1_1174 NAND2X1_557/Y AOI21X1_39/Y NAND2X1_558/Y gnd OAI21X1_1174/Y vdd OAI21X1
XFILL_1_OAI21X1_1350 gnd vdd FILL
XDFFPOSX1_720 BUFX2_387/A CLKBUF1_15/Y OAI21X1_989/Y gnd vdd DFFPOSX1
XDFFPOSX1_731 BUFX2_368/A CLKBUF1_81/Y OAI21X1_1011/Y gnd vdd DFFPOSX1
XOAI21X1_1141 OAI21X1_1141/A BUFX4_186/Y NAND2X1_510/Y gnd OAI21X1_1141/Y vdd OAI21X1
XOAI21X1_1163 INVX1_193/Y OAI21X1_1163/B NAND2X1_543/Y gnd OAI21X1_1163/Y vdd OAI21X1
XFILL_1_OAI21X1_301 gnd vdd FILL
XDFFPOSX1_742 BUFX2_381/A CLKBUF1_57/Y OAI21X1_1033/Y gnd vdd DFFPOSX1
XDFFPOSX1_753 BUFX2_64/A CLKBUF1_12/Y OAI21X1_1045/Y gnd vdd DFFPOSX1
XDFFPOSX1_775 BUFX2_26/A CLKBUF1_89/Y OAI21X1_1067/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_951 gnd vdd FILL
XFILL_1_DFFPOSX1_940 gnd vdd FILL
XFILL_1_OAI21X1_1383 gnd vdd FILL
XFILL_1_OAI21X1_1372 gnd vdd FILL
XOAI21X1_1196 NOR3X1_14/C OR2X2_21/B INVX2_89/Y gnd NAND2X1_581/B vdd OAI21X1
XOAI21X1_1185 NAND2X1_572/Y NOR3X1_12/Y NAND2X1_570/Y gnd OAI21X1_1185/Y vdd OAI21X1
XFILL_0_OAI21X1_130 gnd vdd FILL
XFILL_1_OAI21X1_1361 gnd vdd FILL
XDFFPOSX1_764 BUFX2_14/A CLKBUF1_83/Y OAI21X1_1056/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_163 gnd vdd FILL
XFILL_1_OAI21X1_312 gnd vdd FILL
XFILL_0_OAI21X1_141 gnd vdd FILL
XFILL_1_DFFPOSX1_962 gnd vdd FILL
XFILL_1_OAI21X1_323 gnd vdd FILL
XFILL_1_DFFPOSX1_984 gnd vdd FILL
XFILL_1_OAI21X1_1394 gnd vdd FILL
XDFFPOSX1_786 BUFX2_38/A CLKBUF1_36/Y OAI21X1_1078/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_973 gnd vdd FILL
XDFFPOSX1_797 BUFX2_50/A CLKBUF1_38/Y OAI21X1_1089/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_152 gnd vdd FILL
XFILL_1_OAI21X1_334 gnd vdd FILL
XFILL_2_OAI21X1_516 gnd vdd FILL
XFILL_0_OAI21X1_185 gnd vdd FILL
XFILL_1_OAI21X1_378 gnd vdd FILL
XFILL_1_OAI21X1_367 gnd vdd FILL
XFILL_1_DFFPOSX1_995 gnd vdd FILL
XFILL_0_OAI21X1_196 gnd vdd FILL
XFILL_0_OAI21X1_174 gnd vdd FILL
XFILL_2_OAI21X1_527 gnd vdd FILL
XFILL_1_OAI21X1_345 gnd vdd FILL
XFILL_1_OAI21X1_356 gnd vdd FILL
XFILL_1_OAI21X1_389 gnd vdd FILL
XFILL_0_NAND3X1_16 gnd vdd FILL
XFILL_0_NAND3X1_27 gnd vdd FILL
XFILL_0_NAND3X1_38 gnd vdd FILL
XFILL_0_NAND3X1_49 gnd vdd FILL
XFILL_0_BUFX4_40 gnd vdd FILL
XFILL_0_BUFX4_62 gnd vdd FILL
XFILL_0_BUFX4_51 gnd vdd FILL
XFILL_0_BUFX4_95 gnd vdd FILL
XFILL_0_BUFX4_84 gnd vdd FILL
XFILL_1_NAND2X1_340 gnd vdd FILL
XFILL_0_BUFX4_73 gnd vdd FILL
XFILL_1_NAND2X1_351 gnd vdd FILL
XFILL_1_NAND2X1_384 gnd vdd FILL
XFILL_1_NAND2X1_373 gnd vdd FILL
XFILL_1_BUFX4_137 gnd vdd FILL
XFILL_1_BUFX4_126 gnd vdd FILL
XFILL_0_DFFPOSX1_541 gnd vdd FILL
XFILL_1_BUFX4_115 gnd vdd FILL
XFILL_1_BUFX4_104 gnd vdd FILL
XFILL_0_DFFPOSX1_530 gnd vdd FILL
XFILL_0_NAND2X1_191 gnd vdd FILL
XFILL_0_NAND2X1_180 gnd vdd FILL
XFILL_1_BUFX4_148 gnd vdd FILL
XFILL_1_BUFX4_159 gnd vdd FILL
XFILL_0_DFFPOSX1_585 gnd vdd FILL
XFILL_0_DFFPOSX1_563 gnd vdd FILL
XFILL_0_DFFPOSX1_574 gnd vdd FILL
XFILL_0_DFFPOSX1_552 gnd vdd FILL
XFILL_0_DFFPOSX1_596 gnd vdd FILL
XFILL_20_11_1 gnd vdd FILL
XFILL_0_OR2X2_21 gnd vdd FILL
XFILL_0_OR2X2_10 gnd vdd FILL
XFILL_1_OAI21X1_890 gnd vdd FILL
XNAND3X1_40 bundleAddress_i[37] bundleAddress_i[36] bundleAddress_i[35] gnd INVX2_98/A
+ vdd NAND3X1
XNAND3X1_62 INVX1_216/A NOR2X1_214/Y NOR3X1_18/Y gnd XNOR2X1_89/A vdd NAND3X1
XNAND3X1_51 bundleAddress_i[5] INVX1_198/Y AND2X2_24/Y gnd NAND3X1_51/Y vdd NAND3X1
XFILL_2_OAI21X1_1001 gnd vdd FILL
XBUFX2_700 BUFX2_700/A gnd pid2_o[5] vdd BUFX2
XFILL_2_DFFPOSX1_613 gnd vdd FILL
XBUFX2_711 BUFX2_711/A gnd pid2_o[23] vdd BUFX2
XFILL_2_DFFPOSX1_602 gnd vdd FILL
XBUFX2_722 BUFX2_722/A gnd pid3_o[14] vdd BUFX2
XBUFX2_733 BUFX2_733/A gnd pid3_o[4] vdd BUFX2
XFILL_2_DFFPOSX1_624 gnd vdd FILL
XFILL_2_OAI21X1_1067 gnd vdd FILL
XFILL_3_DFFPOSX1_60 gnd vdd FILL
XBUFX2_744 BUFX2_744/A gnd pid3_o[22] vdd BUFX2
XNOR2X1_51 INVX2_34/Y NOR3X1_8/A gnd NOR2X1_51/Y vdd NOR2X1
XBUFX2_755 BUFX2_755/A gnd pid4_o[13] vdd BUFX2
XFILL_3_DFFPOSX1_71 gnd vdd FILL
XNOR2X1_73 NOR2X1_73/A INVX8_6/A gnd NOR2X1_73/Y vdd NOR2X1
XFILL_2_DFFPOSX1_635 gnd vdd FILL
XFILL_2_DFFPOSX1_657 gnd vdd FILL
XFILL_2_DFFPOSX1_646 gnd vdd FILL
XNOR2X1_40 bundleStartMajId_i[16] AND2X2_8/Y gnd NOR2X1_40/Y vdd NOR2X1
XNOR2X1_62 OR2X2_1/Y NOR2X1_62/B gnd NOR2X1_62/Y vdd NOR2X1
XFILL_2_DFFPOSX1_679 gnd vdd FILL
XBUFX2_788 BUFX2_788/A gnd tid1_o[44] vdd BUFX2
XFILL_2_DFFPOSX1_668 gnd vdd FILL
XFILL_3_DFFPOSX1_82 gnd vdd FILL
XBUFX2_777 BUFX2_777/A gnd tid1_o[63] vdd BUFX2
XBUFX2_766 BUFX2_766/A gnd pid4_o[3] vdd BUFX2
XFILL_3_DFFPOSX1_93 gnd vdd FILL
XNOR2X1_95 OR2X2_13/B NOR2X1_97/B gnd NOR2X1_95/Y vdd NOR2X1
XNOR2X1_84 INVX1_31/A OR2X2_9/A gnd NOR2X1_84/Y vdd NOR2X1
XFILL_0_NOR2X1_128 gnd vdd FILL
XFILL_0_NOR2X1_117 gnd vdd FILL
XFILL_0_NOR2X1_106 gnd vdd FILL
XBUFX2_799 BUFX2_799/A gnd tid1_o[34] vdd BUFX2
XFILL_31_8_1 gnd vdd FILL
XFILL_0_NOR2X1_139 gnd vdd FILL
XFILL_30_3_0 gnd vdd FILL
XFILL_25_10_1 gnd vdd FILL
XFILL_1_DFFPOSX1_214 gnd vdd FILL
XFILL_0_BUFX2_440 gnd vdd FILL
XFILL_1_DFFPOSX1_203 gnd vdd FILL
XFILL_1_DFFPOSX1_247 gnd vdd FILL
XFILL_1_DFFPOSX1_225 gnd vdd FILL
XFILL_0_BUFX2_473 gnd vdd FILL
XFILL_0_BUFX2_484 gnd vdd FILL
XFILL_0_BUFX2_451 gnd vdd FILL
XFILL_0_BUFX2_462 gnd vdd FILL
XFILL_1_DFFPOSX1_236 gnd vdd FILL
XFILL_1_DFFPOSX1_258 gnd vdd FILL
XNAND2X1_108 BUFX2_423/A BUFX4_351/Y gnd OAI21X1_364/C vdd NAND2X1
XFILL_0_BUFX2_495 gnd vdd FILL
XFILL_1_DFFPOSX1_269 gnd vdd FILL
XNAND2X1_119 BUFX2_435/A BUFX4_362/Y gnd OAI21X1_375/C vdd NAND2X1
XFILL_4_DFFPOSX1_718 gnd vdd FILL
XFILL_4_DFFPOSX1_729 gnd vdd FILL
XNAND2X1_6 NAND2X1_6/A OAI21X1_6/A gnd OAI21X1_6/C vdd NAND2X1
XFILL_4_DFFPOSX1_707 gnd vdd FILL
XFILL_1_OAI21X1_39 gnd vdd FILL
XFILL_1_OAI21X1_17 gnd vdd FILL
XFILL_1_OAI21X1_28 gnd vdd FILL
XFILL_38_4_0 gnd vdd FILL
XNOR2X1_130 INVX2_96/A NOR2X1_130/B gnd NOR2X1_130/Y vdd NOR2X1
XNOR2X1_152 INVX1_189/A NOR2X1_152/B gnd AND2X2_23/B vdd NOR2X1
XNOR2X1_141 INVX1_202/A NOR2X1_141/B gnd XNOR2X1_62/A vdd NOR2X1
XFILL_0_11_1 gnd vdd FILL
XFILL_0_NAND2X1_60 gnd vdd FILL
XFILL_0_NAND2X1_71 gnd vdd FILL
XFILL_0_NAND2X1_82 gnd vdd FILL
XNOR2X1_185 NOR2X1_185/A NOR2X1_185/B gnd AND2X2_26/A vdd NOR2X1
XNOR2X1_163 NOR2X1_204/A NOR2X1_163/B gnd INVX2_111/A vdd NOR2X1
XNOR2X1_174 bundleAddress_i[4] NOR2X1_174/B gnd NOR2X1_174/Y vdd NOR2X1
XFILL_0_NAND2X1_93 gnd vdd FILL
XFILL_27_18_0 gnd vdd FILL
XNOR2X1_196 INVX4_40/Y INVX1_192/A gnd NOR2X1_196/Y vdd NOR2X1
XFILL_22_8_1 gnd vdd FILL
XFILL_1_BUFX2_608 gnd vdd FILL
XFILL_1_BUFX2_619 gnd vdd FILL
XFILL_21_3_0 gnd vdd FILL
XOAI21X1_614 AOI21X1_14/Y OAI21X1_614/B OAI21X1_614/C gnd OAI21X1_614/Y vdd OAI21X1
XOAI21X1_603 AOI21X1_10/Y NOR3X1_5/Y NOR2X1_89/B gnd OAI21X1_604/C vdd OAI21X1
XFILL_3_DFFPOSX1_319 gnd vdd FILL
XOAI21X1_647 BUFX4_3/A BUFX4_386/Y BUFX2_576/A gnd OAI21X1_649/C vdd OAI21X1
XFILL_3_DFFPOSX1_308 gnd vdd FILL
XOAI21X1_636 BUFX4_3/Y BUFX4_346/Y BUFX2_571/A gnd OAI21X1_637/C vdd OAI21X1
XOAI21X1_625 XNOR2X1_37/Y BUFX4_134/Y OAI21X1_625/C gnd OAI21X1_625/Y vdd OAI21X1
XOAI21X1_658 BUFX4_145/Y BUFX4_63/Y BUFX2_585/A gnd OAI21X1_659/C vdd OAI21X1
XOAI21X1_669 OAI21X1_669/A BUFX4_296/Y OAI21X1_669/C gnd OAI21X1_669/Y vdd OAI21X1
XDFFPOSX1_550 BUFX2_597/A CLKBUF1_80/Y OAI21X1_665/Y gnd vdd DFFPOSX1
XDFFPOSX1_583 BUFX2_614/A CLKBUF1_19/Y OAI21X1_759/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1180 gnd vdd FILL
XDFFPOSX1_572 BUFX2_602/A CLKBUF1_63/Y OAI21X1_729/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1191 gnd vdd FILL
XDFFPOSX1_561 BUFX2_590/A CLKBUF1_46/Y OAI21X1_697/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_120 gnd vdd FILL
XFILL_1_DFFPOSX1_792 gnd vdd FILL
XFILL_1_OAI21X1_142 gnd vdd FILL
XFILL_1_DFFPOSX1_770 gnd vdd FILL
XXNOR2X1_19 XNOR2X1_19/A INVX4_21/Y gnd XNOR2X1_19/Y vdd XNOR2X1
XNAND2X1_620 AND2X2_33/B INVX2_107/Y gnd NOR3X1_18/B vdd NAND2X1
XDFFPOSX1_594 BUFX2_626/A CLKBUF1_90/Y OAI21X1_792/Y gnd vdd DFFPOSX1
XFILL_2_OAI21X1_324 gnd vdd FILL
XFILL_1_OAI21X1_153 gnd vdd FILL
XFILL_1_OAI21X1_131 gnd vdd FILL
XFILL_1_DFFPOSX1_781 gnd vdd FILL
XFILL_1_OAI21X1_186 gnd vdd FILL
XNAND2X1_664 BUFX2_655/A BUFX4_313/Y gnd NAND2X1_664/Y vdd NAND2X1
XNAND2X1_653 BUFX2_672/A BUFX4_311/Y gnd NAND2X1_653/Y vdd NAND2X1
XNAND2X1_642 OR2X2_21/A NAND2X1_642/B gnd NAND2X1_642/Y vdd NAND2X1
XNAND2X1_631 bundleAddress_i[39] XNOR2X1_96/A gnd XNOR2X1_97/A vdd NAND2X1
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XFILL_1_OAI21X1_164 gnd vdd FILL
XFILL_1_OAI21X1_175 gnd vdd FILL
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XNAND2X1_697 BUFX2_688/A BUFX4_218/Y gnd NAND2X1_697/Y vdd NAND2X1
XINVX1_65 INVX1_65/A gnd INVX1_65/Y vdd INVX1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XNAND2X1_686 BUFX2_707/A BUFX4_180/Y gnd NAND2X1_686/Y vdd NAND2X1
XFILL_1_OAI21X1_197 gnd vdd FILL
XINVX1_76 INVX1_76/A gnd INVX1_76/Y vdd INVX1
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XFILL_5_9_1 gnd vdd FILL
XNAND2X1_675 BUFX2_667/A BUFX4_326/Y gnd NAND2X1_675/Y vdd NAND2X1
XFILL_29_4_0 gnd vdd FILL
XINVX1_98 bundle_i[42] gnd INVX1_98/Y vdd INVX1
XINVX1_87 bundle_i[53] gnd INVX1_87/Y vdd INVX1
XBUFX2_18 BUFX2_18/A gnd addr1_o[39] vdd BUFX2
XFILL_4_4_0 gnd vdd FILL
XFILL_5_10_1 gnd vdd FILL
XBUFX2_29 BUFX2_29/A gnd addr1_o[29] vdd BUFX2
XDFFPOSX1_6 BUFX2_693/A CLKBUF1_99/Y DFFPOSX1_6/D gnd vdd DFFPOSX1
XFILL_13_8_1 gnd vdd FILL
XFILL_1_NAND2X1_192 gnd vdd FILL
XFILL_0_DFFPOSX1_360 gnd vdd FILL
XFILL_1_NAND2X1_181 gnd vdd FILL
XFILL_1_BUFX4_18 gnd vdd FILL
XFILL_0_DFFPOSX1_382 gnd vdd FILL
XFILL_12_3_0 gnd vdd FILL
XFILL_0_DFFPOSX1_393 gnd vdd FILL
XFILL_0_DFFPOSX1_371 gnd vdd FILL
XFILL_1_BUFX4_29 gnd vdd FILL
XFILL_3_DFFPOSX1_820 gnd vdd FILL
XFILL_3_DFFPOSX1_831 gnd vdd FILL
XFILL_3_DFFPOSX1_875 gnd vdd FILL
XFILL_3_DFFPOSX1_853 gnd vdd FILL
XFILL_3_DFFPOSX1_842 gnd vdd FILL
XFILL_3_DFFPOSX1_864 gnd vdd FILL
XFILL_3_DFFPOSX1_886 gnd vdd FILL
XFILL_3_DFFPOSX1_897 gnd vdd FILL
XNOR2X1_9 NOR2X1_9/A NOR2X1_9/B gnd NOR2X1_9/Y vdd NOR2X1
XFILL_7_18_0 gnd vdd FILL
XFILL_2_DFFPOSX1_421 gnd vdd FILL
XFILL_11_16_1 gnd vdd FILL
XFILL_2_DFFPOSX1_410 gnd vdd FILL
XFILL_2_DFFPOSX1_432 gnd vdd FILL
XBUFX2_530 BUFX2_530/A gnd majID3_o[46] vdd BUFX2
XFILL_4_DFFPOSX1_50 gnd vdd FILL
XBUFX2_563 BUFX2_563/A gnd majID3_o[16] vdd BUFX2
XFILL_2_DFFPOSX1_443 gnd vdd FILL
XFILL_2_DFFPOSX1_465 gnd vdd FILL
XBUFX2_552 BUFX2_552/A gnd majID3_o[26] vdd BUFX2
XBUFX2_541 BUFX2_541/A gnd majID3_o[36] vdd BUFX2
XFILL_2_DFFPOSX1_454 gnd vdd FILL
XFILL_0_OAI21X1_1709 gnd vdd FILL
XBUFX2_574 BUFX2_574/A gnd majID3_o[6] vdd BUFX2
XFILL_4_DFFPOSX1_83 gnd vdd FILL
XBUFX2_596 BUFX2_596/A gnd majID4_o[44] vdd BUFX2
XFILL_4_DFFPOSX1_61 gnd vdd FILL
XBUFX2_585 BUFX2_585/A gnd majID4_o[63] vdd BUFX2
XFILL_2_DFFPOSX1_476 gnd vdd FILL
XFILL_4_DFFPOSX1_72 gnd vdd FILL
XFILL_2_DFFPOSX1_498 gnd vdd FILL
XFILL_2_DFFPOSX1_487 gnd vdd FILL
XFILL_4_DFFPOSX1_94 gnd vdd FILL
XFILL_5_DFFPOSX1_903 gnd vdd FILL
XFILL_5_DFFPOSX1_936 gnd vdd FILL
XFILL_5_DFFPOSX1_947 gnd vdd FILL
XFILL_5_DFFPOSX1_914 gnd vdd FILL
XFILL_5_DFFPOSX1_925 gnd vdd FILL
XFILL_5_DFFPOSX1_969 gnd vdd FILL
XFILL_5_DFFPOSX1_958 gnd vdd FILL
XAOI21X1_19 bundleStartMajId_i[12] NOR2X1_94/Y bundleStartMajId_i[11] gnd AOI21X1_19/Y
+ vdd AOI21X1
XFILL_0_BUFX2_270 gnd vdd FILL
XFILL_0_AND2X2_5 gnd vdd FILL
XFILL_0_BUFX2_281 gnd vdd FILL
XFILL_0_BUFX2_292 gnd vdd FILL
XFILL_4_DFFPOSX1_515 gnd vdd FILL
XFILL_4_DFFPOSX1_537 gnd vdd FILL
XFILL_4_DFFPOSX1_526 gnd vdd FILL
XFILL_16_15_1 gnd vdd FILL
XFILL_4_DFFPOSX1_504 gnd vdd FILL
XFILL_4_DFFPOSX1_548 gnd vdd FILL
XFILL_4_DFFPOSX1_559 gnd vdd FILL
XFILL_10_11_0 gnd vdd FILL
XFILL_1_BUFX2_1017 gnd vdd FILL
XFILL_1_BUFX2_1006 gnd vdd FILL
XFILL_1_BUFX2_416 gnd vdd FILL
XFILL_1_BUFX2_405 gnd vdd FILL
XFILL_1_BUFX2_427 gnd vdd FILL
XOAI21X1_411 OAI21X1_411/A NOR2X1_5/Y OAI21X1_411/C gnd OAI21X1_411/Y vdd OAI21X1
XOAI21X1_422 XNOR2X1_5/Y BUFX4_215/Y OAI21X1_422/C gnd OAI21X1_422/Y vdd OAI21X1
XOAI21X1_400 NOR2X1_3/Y bundleStartMajId_i[59] BUFX4_244/Y gnd OAI21X1_401/B vdd OAI21X1
XFILL_3_DFFPOSX1_127 gnd vdd FILL
XFILL_3_DFFPOSX1_116 gnd vdd FILL
XOAI21X1_455 XNOR2X1_16/Y BUFX4_221/Y OAI21X1_455/C gnd OAI21X1_455/Y vdd OAI21X1
XFILL_1_CLKBUF1_18 gnd vdd FILL
XFILL_3_DFFPOSX1_105 gnd vdd FILL
XOAI21X1_444 XNOR2X1_11/Y BUFX4_214/Y OAI21X1_444/C gnd OAI21X1_444/Y vdd OAI21X1
XOAI21X1_433 XNOR2X1_8/Y BUFX4_194/Y OAI21X1_433/C gnd OAI21X1_433/Y vdd OAI21X1
XOAI21X1_466 OAI21X1_466/A NOR3X1_2/Y OAI21X1_466/C gnd OAI21X1_466/Y vdd OAI21X1
XFILL_3_DFFPOSX1_138 gnd vdd FILL
XFILL_3_DFFPOSX1_149 gnd vdd FILL
XFILL_1_CLKBUF1_29 gnd vdd FILL
XOAI21X1_477 OAI21X1_477/A NOR2X1_45/Y OAI21X1_477/C gnd OAI21X1_477/Y vdd OAI21X1
XOAI21X1_499 OAI21X1_499/A INVX4_28/Y INVX2_39/Y gnd NAND3X1_13/C vdd OAI21X1
XOAI21X1_488 OAI21X1_493/A INVX2_37/Y INVX4_25/Y gnd OAI21X1_488/Y vdd OAI21X1
XFILL_3_XNOR2X1_90 gnd vdd FILL
XFILL_6_DFFPOSX1_609 gnd vdd FILL
XDFFPOSX1_391 BUFX2_422/A CLKBUF1_92/Y OAI21X1_363/Y gnd vdd DFFPOSX1
XDFFPOSX1_380 BUFX2_410/A CLKBUF1_15/Y OAI21X1_352/Y gnd vdd DFFPOSX1
XFILL_2_OAI21X1_110 gnd vdd FILL
XFILL_34_16_1 gnd vdd FILL
XNAND2X1_472 bundleAddress_i[59] bundleAddress_i[58] gnd INVX1_185/A vdd NAND2X1
XNAND2X1_450 BUFX2_44/A BUFX4_348/Y gnd NAND2X1_450/Y vdd NAND2X1
XNAND2X1_461 BUFX2_56/A BUFX4_348/Y gnd NAND2X1_461/Y vdd NAND2X1
XNAND2X1_494 bundleAddress_i[53] bundleAddress_i[50] gnd NOR2X1_130/B vdd NAND2X1
XNAND2X1_483 BUFX2_128/A BUFX4_204/Y gnd NAND2X1_483/Y vdd NAND2X1
XFILL_15_10_0 gnd vdd FILL
XFILL_0_INVX1_204 gnd vdd FILL
XFILL_0_INVX1_215 gnd vdd FILL
XFILL_0_INVX1_226 gnd vdd FILL
XFILL_0_DFFPOSX1_190 gnd vdd FILL
XFILL_0_OAI21X1_14 gnd vdd FILL
XFILL_0_OAI21X1_25 gnd vdd FILL
XFILL_1_BUFX2_972 gnd vdd FILL
XFILL_1_BUFX2_983 gnd vdd FILL
XFILL_0_OAI21X1_47 gnd vdd FILL
XFILL_0_OAI21X1_36 gnd vdd FILL
XFILL_0_OAI21X1_58 gnd vdd FILL
XOAI21X1_1729 INVX2_126/Y BUFX4_301/Y OAI21X1_1729/C gnd DFFPOSX1_77/D vdd OAI21X1
XFILL_1_BUFX2_994 gnd vdd FILL
XFILL_3_DFFPOSX1_650 gnd vdd FILL
XFILL_0_OAI21X1_69 gnd vdd FILL
XOAI21X1_1718 BUFX4_134/Y BUFX4_76/Y BUFX2_771/A gnd OAI21X1_1719/C vdd OAI21X1
XOAI21X1_1707 BUFX4_163/Y INVX2_115/Y OAI21X1_1707/C gnd DFFPOSX1_66/D vdd OAI21X1
XFILL_3_DFFPOSX1_672 gnd vdd FILL
XFILL_3_DFFPOSX1_683 gnd vdd FILL
XFILL_3_DFFPOSX1_661 gnd vdd FILL
XFILL_3_DFFPOSX1_694 gnd vdd FILL
XFILL_0_OAI21X1_718 gnd vdd FILL
XFILL_0_OAI21X1_707 gnd vdd FILL
XFILL_0_OAI21X1_729 gnd vdd FILL
XFILL_8_1 gnd vdd FILL
XFILL_33_11_0 gnd vdd FILL
XFILL_0_NAND2X1_702 gnd vdd FILL
XFILL_36_7_1 gnd vdd FILL
XFILL_2_DFFPOSX1_240 gnd vdd FILL
XFILL_0_NAND2X1_724 gnd vdd FILL
XFILL_0_OAI21X1_1506 gnd vdd FILL
XFILL_0_NAND2X1_735 gnd vdd FILL
XFILL_0_NAND2X1_713 gnd vdd FILL
XFILL_2_DFFPOSX1_273 gnd vdd FILL
XFILL_0_NAND2X1_768 gnd vdd FILL
XFILL_2_DFFPOSX1_262 gnd vdd FILL
XFILL_35_2_0 gnd vdd FILL
XFILL_2_DFFPOSX1_251 gnd vdd FILL
XFILL_0_NAND2X1_746 gnd vdd FILL
XFILL_0_OAI21X1_1528 gnd vdd FILL
XFILL_0_OAI21X1_1517 gnd vdd FILL
XFILL_0_OAI21X1_1539 gnd vdd FILL
XBUFX2_360 BUFX2_360/A gnd instr4_o[20] vdd BUFX2
XBUFX2_371 BUFX2_371/A gnd instr4_o[10] vdd BUFX2
XFILL_0_NAND2X1_757 gnd vdd FILL
XFILL_2_DFFPOSX1_284 gnd vdd FILL
XFILL_5_DFFPOSX1_51 gnd vdd FILL
XFILL_5_DFFPOSX1_62 gnd vdd FILL
XFILL_1_NOR3X1_10 gnd vdd FILL
XBUFX2_382 BUFX2_382/A gnd instr4_o[0] vdd BUFX2
XFILL_5_DFFPOSX1_40 gnd vdd FILL
XBUFX2_393 BUFX2_393/A gnd majID1_o[63] vdd BUFX2
XFILL_2_DFFPOSX1_295 gnd vdd FILL
XFILL_5_DFFPOSX1_73 gnd vdd FILL
XFILL_5_DFFPOSX1_700 gnd vdd FILL
XFILL_5_DFFPOSX1_84 gnd vdd FILL
XFILL_5_DFFPOSX1_711 gnd vdd FILL
XFILL_5_DFFPOSX1_95 gnd vdd FILL
XFILL_5_DFFPOSX1_755 gnd vdd FILL
XFILL_5_DFFPOSX1_744 gnd vdd FILL
XFILL_5_DFFPOSX1_722 gnd vdd FILL
XFILL_5_DFFPOSX1_733 gnd vdd FILL
XOAI21X1_60 INVX2_198/Y BUFX4_190/Y OAI21X1_60/C gnd OAI21X1_60/Y vdd OAI21X1
XOAI21X1_71 INVX2_7/Y BUFX4_196/Y OAI21X1_71/C gnd OAI21X1_71/Y vdd OAI21X1
XFILL_5_DFFPOSX1_788 gnd vdd FILL
XFILL_5_DFFPOSX1_777 gnd vdd FILL
XOAI21X1_93 BUFX4_129/Y INVX2_156/Y OAI21X1_93/C gnd OAI21X1_93/Y vdd OAI21X1
XFILL_5_DFFPOSX1_766 gnd vdd FILL
XOAI21X1_82 BUFX4_12/Y BUFX4_374/Y BUFX2_950/A gnd OAI21X1_83/C vdd OAI21X1
XFILL_5_DFFPOSX1_799 gnd vdd FILL
XFILL_38_10_0 gnd vdd FILL
XFILL_4_DFFPOSX1_301 gnd vdd FILL
XFILL_4_DFFPOSX1_312 gnd vdd FILL
XFILL_4_DFFPOSX1_345 gnd vdd FILL
XFILL_4_DFFPOSX1_323 gnd vdd FILL
XFILL_0_DFFPOSX1_80 gnd vdd FILL
XFILL_4_DFFPOSX1_334 gnd vdd FILL
XFILL_0_DFFPOSX1_91 gnd vdd FILL
XFILL_2_DFFPOSX1_1004 gnd vdd FILL
XFILL_4_DFFPOSX1_356 gnd vdd FILL
XFILL_4_DFFPOSX1_378 gnd vdd FILL
XFILL_4_DFFPOSX1_367 gnd vdd FILL
XFILL_2_DFFPOSX1_1026 gnd vdd FILL
XFILL_27_7_1 gnd vdd FILL
XFILL_2_DFFPOSX1_1015 gnd vdd FILL
XFILL_2_7_1 gnd vdd FILL
XFILL_4_DFFPOSX1_389 gnd vdd FILL
XFILL_26_2_0 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XFILL_1_BUFX2_213 gnd vdd FILL
XFILL_1_BUFX2_224 gnd vdd FILL
XOAI21X1_230 BUFX4_132/Y BUFX4_82/Y BUFX2_976/A gnd OAI21X1_231/C vdd OAI21X1
XOAI21X1_241 INVX2_166/Y BUFX4_289/Y OAI21X1_241/C gnd OAI21X1_241/Y vdd OAI21X1
XFILL_10_6_1 gnd vdd FILL
XFILL_1_BUFX2_268 gnd vdd FILL
XFILL_1_BUFX2_257 gnd vdd FILL
XOAI21X1_252 BUFX4_148/Y BUFX4_36/Y BUFX2_988/A gnd OAI21X1_253/C vdd OAI21X1
XOAI21X1_274 BUFX4_150/Y BUFX4_52/Y BUFX2_1000/A gnd OAI21X1_275/C vdd OAI21X1
XOAI21X1_263 INVX2_177/Y BUFX4_296/Y OAI21X1_263/C gnd OAI21X1_263/Y vdd OAI21X1
XFILL_1_BUFX2_279 gnd vdd FILL
XOAI21X1_296 BUFX4_138/Y BUFX4_67/Y BUFX2_1012/A gnd OAI21X1_297/C vdd OAI21X1
XOAI21X1_285 INVX2_188/Y INVX8_2/A OAI21X1_285/C gnd OAI21X1_285/Y vdd OAI21X1
XAND2X2_30 AND2X2_30/A INVX2_75/Y gnd AND2X2_30/Y vdd AND2X2
XFILL_6_DFFPOSX1_406 gnd vdd FILL
XFILL_9_3_0 gnd vdd FILL
XNAND2X1_280 bundleStartMajId_i[40] NOR2X1_68/Y gnd XNOR2X1_31/A vdd NAND2X1
XNAND2X1_291 INVX2_48/A NOR2X1_75/Y gnd NOR3X1_5/C vdd NAND2X1
XFILL_4_DFFPOSX1_890 gnd vdd FILL
XFILL_18_7_1 gnd vdd FILL
XFILL_17_2_0 gnd vdd FILL
XFILL_1_NAND3X1_9 gnd vdd FILL
XFILL_0_INVX8_4 gnd vdd FILL
XFILL_5_DFFPOSX1_1019 gnd vdd FILL
XFILL_5_DFFPOSX1_1008 gnd vdd FILL
XFILL_1_BUFX2_780 gnd vdd FILL
XFILL_1_BUFX2_791 gnd vdd FILL
XFILL_0_BUFX4_332 gnd vdd FILL
XFILL_0_BUFX4_310 gnd vdd FILL
XFILL_0_BUFX4_321 gnd vdd FILL
XOAI21X1_1504 BUFX4_158/Y BUFX4_68/Y BUFX2_228/A gnd OAI21X1_1505/C vdd OAI21X1
XFILL_0_BUFX4_343 gnd vdd FILL
XDFFPOSX1_19 BUFX2_688/A CLKBUF1_57/Y DFFPOSX1_19/D gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1713 gnd vdd FILL
XFILL_1_OAI21X1_1724 gnd vdd FILL
XOAI21X1_1526 INVX1_225/A INVX2_82/Y BUFX4_284/Y gnd OAI21X1_1527/B vdd OAI21X1
XOAI21X1_1515 BUFX4_170/Y BUFX4_53/Y BUFX2_232/A gnd OAI21X1_1517/C vdd OAI21X1
XFILL_1_OAI21X1_1702 gnd vdd FILL
XFILL_0_BUFX4_376 gnd vdd FILL
XFILL_0_BUFX4_365 gnd vdd FILL
XOAI21X1_1537 NAND2X1_571/Y OR2X2_21/A OAI21X1_1537/C gnd OAI21X1_1539/A vdd OAI21X1
XOAI21X1_1548 BUFX4_139/Y BUFX4_73/Y BUFX2_243/A gnd OAI21X1_1549/C vdd OAI21X1
XFILL_0_BUFX4_354 gnd vdd FILL
XFILL_1_OAI21X1_1757 gnd vdd FILL
XFILL_1_OAI21X1_1746 gnd vdd FILL
XFILL_3_DFFPOSX1_480 gnd vdd FILL
XFILL_1_OAI21X1_1735 gnd vdd FILL
XOAI21X1_1559 BUFX4_121/Y BUFX4_59/Y BUFX2_247/A gnd OAI21X1_1560/C vdd OAI21X1
XFILL_0_OAI21X1_504 gnd vdd FILL
XFILL_3_DFFPOSX1_491 gnd vdd FILL
XFILL_0_BUFX4_387 gnd vdd FILL
XFILL_0_BUFX2_1003 gnd vdd FILL
XFILL_0_OAI21X1_526 gnd vdd FILL
XFILL_1_OAI21X1_1768 gnd vdd FILL
XFILL_1_OAI21X1_708 gnd vdd FILL
XFILL_0_BUFX2_1025 gnd vdd FILL
XFILL_0_OAI21X1_537 gnd vdd FILL
XFILL_0_OAI21X1_515 gnd vdd FILL
XFILL_0_BUFX2_1014 gnd vdd FILL
XFILL_1_OAI21X1_1779 gnd vdd FILL
XFILL_0_OAI21X1_559 gnd vdd FILL
XFILL_1_OAI21X1_719 gnd vdd FILL
XFILL_0_OAI21X1_548 gnd vdd FILL
XFILL_6_DFFPOSX1_962 gnd vdd FILL
XFILL_6_DFFPOSX1_973 gnd vdd FILL
XFILL_6_DFFPOSX1_984 gnd vdd FILL
XFILL_6_DFFPOSX1_995 gnd vdd FILL
XFILL_0_CLKBUF1_26 gnd vdd FILL
XFILL_0_CLKBUF1_15 gnd vdd FILL
XFILL_0_CLKBUF1_59 gnd vdd FILL
XFILL_0_CLKBUF1_48 gnd vdd FILL
XFILL_0_NAND2X1_510 gnd vdd FILL
XFILL_0_CLKBUF1_37 gnd vdd FILL
XFILL_0_NAND2X1_532 gnd vdd FILL
XFILL_1_NAND2X1_703 gnd vdd FILL
XFILL_0_NAND2X1_521 gnd vdd FILL
XFILL_1_NAND2X1_714 gnd vdd FILL
XFILL_0_OAI21X1_1303 gnd vdd FILL
XFILL_0_OAI21X1_1314 gnd vdd FILL
XFILL_0_NAND2X1_543 gnd vdd FILL
XFILL_1_NAND2X1_736 gnd vdd FILL
XFILL_0_OAI21X1_1336 gnd vdd FILL
XFILL_0_DFFPOSX1_904 gnd vdd FILL
XFILL_0_NAND2X1_554 gnd vdd FILL
XFILL_0_DFFPOSX1_915 gnd vdd FILL
XFILL_0_NAND2X1_587 gnd vdd FILL
XFILL_0_NAND2X1_565 gnd vdd FILL
XFILL_0_OAI21X1_1325 gnd vdd FILL
XFILL_0_OAI21X1_1347 gnd vdd FILL
XFILL_0_OAI21X1_1358 gnd vdd FILL
XFILL_1_NAND2X1_747 gnd vdd FILL
XFILL_0_NAND2X1_576 gnd vdd FILL
XBUFX2_190 BUFX2_190/A gnd addr3_o[56] vdd BUFX2
XFILL_1_NAND2X1_769 gnd vdd FILL
XFILL_6_DFFPOSX1_52 gnd vdd FILL
XFILL_0_DFFPOSX1_948 gnd vdd FILL
XFILL_0_NAND2X1_598 gnd vdd FILL
XFILL_0_DFFPOSX1_937 gnd vdd FILL
XFILL_0_OAI21X1_1369 gnd vdd FILL
XFILL_0_DFFPOSX1_959 gnd vdd FILL
XFILL_0_DFFPOSX1_926 gnd vdd FILL
XFILL_6_DFFPOSX1_85 gnd vdd FILL
XFILL_6_DFFPOSX1_63 gnd vdd FILL
XFILL_6_DFFPOSX1_96 gnd vdd FILL
XFILL_5_DFFPOSX1_530 gnd vdd FILL
XFILL_6_DFFPOSX1_74 gnd vdd FILL
XFILL_5_DFFPOSX1_541 gnd vdd FILL
XFILL_5_DFFPOSX1_563 gnd vdd FILL
XFILL_5_DFFPOSX1_552 gnd vdd FILL
XFILL_5_DFFPOSX1_585 gnd vdd FILL
XFILL_5_DFFPOSX1_596 gnd vdd FILL
XFILL_24_16_0 gnd vdd FILL
XFILL_5_DFFPOSX1_574 gnd vdd FILL
XFILL_0_OR2X2_9 gnd vdd FILL
XFILL_1_BUFX4_7 gnd vdd FILL
XFILL_1_AOI21X1_3 gnd vdd FILL
XCLKBUF1_50 BUFX4_91/Y gnd CLKBUF1_50/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_120 gnd vdd FILL
XFILL_4_DFFPOSX1_153 gnd vdd FILL
XFILL_4_DFFPOSX1_131 gnd vdd FILL
XCLKBUF1_61 BUFX4_83/Y gnd CLKBUF1_61/Y vdd CLKBUF1
XCLKBUF1_72 BUFX4_85/Y gnd CLKBUF1_72/Y vdd CLKBUF1
XCLKBUF1_83 BUFX4_86/Y gnd CLKBUF1_83/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_142 gnd vdd FILL
XFILL_4_DFFPOSX1_175 gnd vdd FILL
XFILL_4_DFFPOSX1_164 gnd vdd FILL
XFILL_1_DFFPOSX1_70 gnd vdd FILL
XFILL_4_DFFPOSX1_186 gnd vdd FILL
XFILL_1_DFFPOSX1_92 gnd vdd FILL
XFILL_1_DFFPOSX1_81 gnd vdd FILL
XCLKBUF1_94 BUFX4_90/Y gnd CLKBUF1_94/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_197 gnd vdd FILL
XFILL_2_BUFX4_241 gnd vdd FILL
XFILL_2_BUFX4_274 gnd vdd FILL
XFILL_2_BUFX4_285 gnd vdd FILL
XFILL_29_15_0 gnd vdd FILL
XFILL_0_BUFX2_814 gnd vdd FILL
XFILL_0_BUFX2_825 gnd vdd FILL
XFILL_0_BUFX2_803 gnd vdd FILL
XFILL_1_OAI21X1_1009 gnd vdd FILL
XFILL_0_BUFX2_847 gnd vdd FILL
XFILL_0_BUFX2_858 gnd vdd FILL
XINVX1_124 bundle_i[80] gnd INVX1_124/Y vdd INVX1
XFILL_0_BUFX2_836 gnd vdd FILL
XINVX1_102 bundle_i[38] gnd INVX1_102/Y vdd INVX1
XINVX1_113 bundle_i[91] gnd INVX1_113/Y vdd INVX1
XFILL_0_BUFX2_869 gnd vdd FILL
XINVX1_157 bundle_i[111] gnd INVX1_157/Y vdd INVX1
XFILL_3_XNOR2X1_1 gnd vdd FILL
XINVX1_146 bundle_i[122] gnd INVX1_146/Y vdd INVX1
XINVX1_168 bundle_i[100] gnd INVX1_168/Y vdd INVX1
XINVX1_135 bundle_i[69] gnd INVX1_135/Y vdd INVX1
XINVX1_179 bundleAddress_i[15] gnd INVX1_179/Y vdd INVX1
XFILL_6_DFFPOSX1_258 gnd vdd FILL
XFILL_6_DFFPOSX1_247 gnd vdd FILL
XFILL_6_DFFPOSX1_269 gnd vdd FILL
XFILL_0_INVX2_12 gnd vdd FILL
XFILL_0_INVX2_34 gnd vdd FILL
XFILL_0_INVX2_45 gnd vdd FILL
XFILL_0_INVX2_23 gnd vdd FILL
XFILL_0_INVX2_67 gnd vdd FILL
XFILL_0_INVX2_56 gnd vdd FILL
XFILL_0_INVX2_89 gnd vdd FILL
XFILL_0_INVX2_78 gnd vdd FILL
XFILL_4_16_0 gnd vdd FILL
XFILL_1_NOR3X1_9 gnd vdd FILL
XFILL_34_4 gnd vdd FILL
XFILL_0_CLKBUF1_2 gnd vdd FILL
XFILL_33_5_1 gnd vdd FILL
XFILL_32_0_0 gnd vdd FILL
XFILL_4_CLKBUF1_1 gnd vdd FILL
XFILL_0_BUFX4_140 gnd vdd FILL
XFILL_0_BUFX4_151 gnd vdd FILL
XOAI21X1_1301 NOR3X1_18/C NOR3X1_18/A OAI21X1_1301/C gnd OAI21X1_1303/A vdd OAI21X1
XOAI21X1_1323 NOR3X1_16/Y bundleAddress_i[21] NOR2X1_202/Y gnd OAI21X1_1324/C vdd
+ OAI21X1
XOAI21X1_1312 BUFX4_6/A BUFX4_370/Y BUFX2_161/A gnd OAI21X1_1313/C vdd OAI21X1
XFILL_0_BUFX4_184 gnd vdd FILL
XFILL_1_OAI21X1_1532 gnd vdd FILL
XDFFPOSX1_902 BUFX2_153/A CLKBUF1_27/Y OAI21X1_1292/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1521 gnd vdd FILL
XFILL_0_BUFX4_162 gnd vdd FILL
XOAI21X1_1334 NOR2X1_203/B INVX1_211/Y BUFX4_310/Y gnd OAI21X1_1335/B vdd OAI21X1
XFILL_1_OAI21X1_1510 gnd vdd FILL
XOAI21X1_1345 BUFX4_12/Y BUFX4_342/Y BUFX2_175/A gnd OAI21X1_1347/C vdd OAI21X1
XDFFPOSX1_924 BUFX2_177/A CLKBUF1_69/Y OAI21X1_1352/Y gnd vdd DFFPOSX1
XOAI21X1_1356 NOR2X1_211/B INVX1_214/A BUFX4_308/Y gnd OAI21X1_1357/B vdd OAI21X1
XFILL_0_BUFX4_173 gnd vdd FILL
XDFFPOSX1_913 BUFX2_165/A CLKBUF1_28/Y OAI21X1_1322/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_301 gnd vdd FILL
XFILL_1_BUFX2_62 gnd vdd FILL
XFILL_0_OAI21X1_312 gnd vdd FILL
XFILL_1_BUFX2_73 gnd vdd FILL
XDFFPOSX1_946 BUFX2_195/A CLKBUF1_72/Y OAI21X1_1415/Y gnd vdd DFFPOSX1
XOAI21X1_1389 bundleAddress_i[61] BUFX4_290/Y OAI21X1_1389/C gnd OAI21X1_1389/Y vdd
+ OAI21X1
XFILL_0_BUFX4_195 gnd vdd FILL
XFILL_1_OAI21X1_1576 gnd vdd FILL
XDFFPOSX1_935 BUFX2_189/A CLKBUF1_97/Y OAI21X1_1383/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1565 gnd vdd FILL
XOAI21X1_1378 NOR2X1_212/Y OAI21X1_1378/B OAI21X1_1378/C gnd OAI21X1_1378/Y vdd OAI21X1
XOAI21X1_1367 AOI21X1_57/Y OAI21X1_1367/B OAI21X1_1367/C gnd OAI21X1_1367/Y vdd OAI21X1
XFILL_1_OAI21X1_1543 gnd vdd FILL
XDFFPOSX1_957 BUFX2_207/A CLKBUF1_34/Y OAI21X1_1447/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1554 gnd vdd FILL
XFILL_1_OAI21X1_1598 gnd vdd FILL
XFILL_1_BUFX2_84 gnd vdd FILL
XDFFPOSX1_968 BUFX2_219/A CLKBUF1_89/Y OAI21X1_1479/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_323 gnd vdd FILL
XDFFPOSX1_979 BUFX2_231/A CLKBUF1_36/Y OAI21X1_1514/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_505 gnd vdd FILL
XFILL_1_OAI21X1_527 gnd vdd FILL
XFILL_0_OAI21X1_345 gnd vdd FILL
XFILL_0_OAI21X1_334 gnd vdd FILL
XFILL_1_OAI21X1_516 gnd vdd FILL
XFILL_1_OAI21X1_1587 gnd vdd FILL
XFILL_0_OAI21X1_378 gnd vdd FILL
XFILL_0_OAI21X1_367 gnd vdd FILL
XFILL_1_OAI21X1_549 gnd vdd FILL
XFILL_1_OAI21X1_538 gnd vdd FILL
XFILL_0_OAI21X1_356 gnd vdd FILL
XFILL_0_OAI21X1_389 gnd vdd FILL
XFILL_9_15_0 gnd vdd FILL
XFILL_6_DFFPOSX1_770 gnd vdd FILL
XFILL_1_OAI21X1_6 gnd vdd FILL
XFILL_13_13_1 gnd vdd FILL
XFILL_0_OAI21X1_1111 gnd vdd FILL
XFILL_0_OAI21X1_1100 gnd vdd FILL
XFILL_0_NAND2X1_362 gnd vdd FILL
XFILL_1_NAND2X1_522 gnd vdd FILL
XFILL_0_OAI21X1_1122 gnd vdd FILL
XFILL_1_NAND2X1_500 gnd vdd FILL
XFILL_0_NAND2X1_340 gnd vdd FILL
XFILL_0_OAI21X1_1133 gnd vdd FILL
XFILL_0_NAND2X1_351 gnd vdd FILL
XFILL_0_NAND2X1_384 gnd vdd FILL
XFILL_0_NAND2X1_373 gnd vdd FILL
XFILL_0_DFFPOSX1_701 gnd vdd FILL
XFILL_0_OAI21X1_1155 gnd vdd FILL
XFILL_0_OAI21X1_1144 gnd vdd FILL
XFILL_24_5_1 gnd vdd FILL
XFILL_1_BUFX4_319 gnd vdd FILL
XFILL_1_BUFX4_308 gnd vdd FILL
XFILL_1_NAND2X1_566 gnd vdd FILL
XFILL_0_DFFPOSX1_734 gnd vdd FILL
XFILL_0_NAND2X1_395 gnd vdd FILL
XFILL_0_DFFPOSX1_712 gnd vdd FILL
XFILL_1_NAND2X1_544 gnd vdd FILL
XFILL_0_DFFPOSX1_723 gnd vdd FILL
XFILL_0_OAI21X1_1166 gnd vdd FILL
XFILL_0_DFFPOSX1_756 gnd vdd FILL
XFILL_0_OAI21X1_1177 gnd vdd FILL
XFILL_23_0_0 gnd vdd FILL
XFILL_0_DFFPOSX1_745 gnd vdd FILL
XFILL_1_NAND2X1_588 gnd vdd FILL
XFILL_0_OAI21X1_1199 gnd vdd FILL
XFILL_1_NAND2X1_599 gnd vdd FILL
XFILL_0_OAI21X1_1188 gnd vdd FILL
XFILL_0_DFFPOSX1_767 gnd vdd FILL
XFILL_1_NAND2X1_577 gnd vdd FILL
XFILL_0_DFFPOSX1_789 gnd vdd FILL
XFILL_0_DFFPOSX1_778 gnd vdd FILL
XFILL_5_DFFPOSX1_360 gnd vdd FILL
XFILL_5_DFFPOSX1_371 gnd vdd FILL
XFILL_5_DFFPOSX1_382 gnd vdd FILL
XFILL_5_DFFPOSX1_393 gnd vdd FILL
XFILL_1_NAND2X1_31 gnd vdd FILL
XINVX4_10 bundleStartMajId_i[39] gnd INVX4_10/Y vdd INVX4
XFILL_1_NAND2X1_64 gnd vdd FILL
XFILL_1_NAND2X1_53 gnd vdd FILL
XINVX4_32 bundleAddress_i[61] gnd INVX4_32/Y vdd INVX4
XINVX4_43 bundleAddress_i[20] gnd INVX4_43/Y vdd INVX4
XINVX4_21 bundleStartMajId_i[20] gnd INVX4_21/Y vdd INVX4
XFILL_1_NAND2X1_75 gnd vdd FILL
XFILL_1_NAND2X1_97 gnd vdd FILL
XFILL_0_OAI21X1_890 gnd vdd FILL
XFILL_18_12_1 gnd vdd FILL
XFILL_7_6_1 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XFILL_2_OAI21X1_1227 gnd vdd FILL
XBUFX2_904 BUFX2_904/A gnd tid2_o[54] vdd BUFX2
XFILL_31_14_1 gnd vdd FILL
XFILL_2_DFFPOSX1_806 gnd vdd FILL
XBUFX2_915 BUFX2_915/A gnd tid3_o[45] vdd BUFX2
XBUFX2_937 BUFX2_937/A gnd tid3_o[25] vdd BUFX2
XFILL_2_DFFPOSX1_82 gnd vdd FILL
XFILL_2_DFFPOSX1_60 gnd vdd FILL
XFILL_2_DFFPOSX1_839 gnd vdd FILL
XFILL_2_DFFPOSX1_817 gnd vdd FILL
XFILL_2_DFFPOSX1_71 gnd vdd FILL
XBUFX2_926 BUFX2_926/A gnd tid3_o[35] vdd BUFX2
XFILL_2_DFFPOSX1_828 gnd vdd FILL
XBUFX2_948 BUFX2_948/A gnd tid3_o[15] vdd BUFX2
XFILL_2_DFFPOSX1_93 gnd vdd FILL
XBUFX2_959 BUFX2_959/A gnd tid3_o[5] vdd BUFX2
XFILL_15_5_1 gnd vdd FILL
XFILL_14_0_0 gnd vdd FILL
XDFFPOSX1_209 BUFX2_881/A CLKBUF1_74/Y OAI21X1_53/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_633 gnd vdd FILL
XFILL_0_BUFX2_611 gnd vdd FILL
XFILL_0_BUFX2_622 gnd vdd FILL
XFILL_0_BUFX2_600 gnd vdd FILL
XFILL_0_BUFX2_644 gnd vdd FILL
XFILL_0_BUFX2_655 gnd vdd FILL
XFILL_1_DFFPOSX1_418 gnd vdd FILL
XFILL_1_DFFPOSX1_407 gnd vdd FILL
XFILL_0_BUFX2_666 gnd vdd FILL
XFILL_1_DFFPOSX1_429 gnd vdd FILL
XFILL_0_BUFX2_688 gnd vdd FILL
XFILL_0_BUFX2_699 gnd vdd FILL
XFILL_0_BUFX2_677 gnd vdd FILL
XFILL_36_13_1 gnd vdd FILL
XBUFX4_230 BUFX4_24/Y gnd BUFX4_230/Y vdd BUFX4
XBUFX4_263 enable_i gnd BUFX4_263/Y vdd BUFX4
XBUFX4_252 INVX8_5/Y gnd BUFX4_9/A vdd BUFX4
XBUFX4_241 INVX8_1/Y gnd BUFX4_241/Y vdd BUFX4
XFILL_0_INVX2_140 gnd vdd FILL
XFILL_0_INVX2_162 gnd vdd FILL
XBUFX4_296 BUFX4_303/A gnd BUFX4_296/Y vdd BUFX4
XBUFX4_274 INVX8_7/Y gnd BUFX4_72/A vdd BUFX4
XBUFX4_285 INVX8_2/Y gnd BUFX4_285/Y vdd BUFX4
XFILL_0_INVX2_151 gnd vdd FILL
XFILL_0_INVX2_173 gnd vdd FILL
XFILL_32_1 gnd vdd FILL
XFILL_0_INVX2_184 gnd vdd FILL
XFILL_0_INVX2_195 gnd vdd FILL
XOAI21X1_829 BUFX4_156/Y BUFX4_82/Y BUFX2_639/A gnd OAI21X1_830/C vdd OAI21X1
XOAI21X1_807 NOR3X1_8/B NOR3X1_8/C OAI21X1_807/C gnd OAI21X1_809/A vdd OAI21X1
XOAI21X1_818 OAI21X1_818/A AOI21X1_34/Y OAI21X1_818/C gnd OAI21X1_818/Y vdd OAI21X1
XOAI21X1_1131 XNOR2X1_59/Y OAI21X1_8/B NAND2X1_499/Y gnd OAI21X1_1131/Y vdd OAI21X1
XOAI21X1_1120 INVX1_186/Y bundleAddress_i[53] BUFX4_241/Y gnd OAI21X1_1121/A vdd OAI21X1
XDFFPOSX1_710 BUFX2_349/A CLKBUF1_99/Y OAI21X1_969/Y gnd vdd DFFPOSX1
XDFFPOSX1_721 BUFX2_388/A CLKBUF1_98/Y OAI21X1_991/Y gnd vdd DFFPOSX1
XOAI21X1_1153 NOR2X1_148/B INVX2_99/Y BUFX4_238/Y gnd OAI21X1_1154/B vdd OAI21X1
XFILL_1_OAI21X1_1340 gnd vdd FILL
XFILL_1_OAI21X1_1351 gnd vdd FILL
XDFFPOSX1_732 BUFX2_370/A CLKBUF1_71/Y OAI21X1_1013/Y gnd vdd DFFPOSX1
XOAI21X1_1164 XNOR2X1_70/Y BUFX4_226/Y NAND2X1_544/Y gnd OAI21X1_1164/Y vdd OAI21X1
XOAI21X1_1142 XNOR2X1_61/Y BUFX4_192/Y NAND2X1_511/Y gnd OAI21X1_1142/Y vdd OAI21X1
XFILL_0_OAI21X1_120 gnd vdd FILL
XFILL_1_OAI21X1_1384 gnd vdd FILL
XFILL_1_DFFPOSX1_952 gnd vdd FILL
XDFFPOSX1_754 BUFX2_3/A CLKBUF1_5/Y OAI21X1_1046/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_941 gnd vdd FILL
XOAI21X1_1175 INVX2_102/A INVX2_82/Y BUFX4_243/Y gnd OAI21X1_1176/B vdd OAI21X1
XDFFPOSX1_743 BUFX2_382/A CLKBUF1_38/Y OAI21X1_1035/Y gnd vdd DFFPOSX1
XOAI21X1_1197 NAND2X1_581/Y NOR2X1_174/B NAND2X1_582/Y gnd OAI21X1_1197/Y vdd OAI21X1
XFILL_1_OAI21X1_1373 gnd vdd FILL
XFILL_1_OAI21X1_302 gnd vdd FILL
XFILL_1_DFFPOSX1_930 gnd vdd FILL
XOAI21X1_1186 NOR3X1_12/Y bundleAddress_i[10] BUFX4_242/Y gnd OAI21X1_1187/B vdd OAI21X1
XFILL_1_OAI21X1_1362 gnd vdd FILL
XDFFPOSX1_765 BUFX2_15/A CLKBUF1_83/Y OAI21X1_1057/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_313 gnd vdd FILL
XFILL_1_DFFPOSX1_985 gnd vdd FILL
XDFFPOSX1_776 BUFX2_27/A CLKBUF1_89/Y OAI21X1_1068/Y gnd vdd DFFPOSX1
XDFFPOSX1_787 BUFX2_39/A CLKBUF1_49/Y OAI21X1_1079/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_963 gnd vdd FILL
XFILL_0_OAI21X1_142 gnd vdd FILL
XFILL_1_OAI21X1_1395 gnd vdd FILL
XFILL_0_OAI21X1_164 gnd vdd FILL
XFILL_1_OAI21X1_324 gnd vdd FILL
XFILL_0_OAI21X1_153 gnd vdd FILL
XFILL_1_OAI21X1_335 gnd vdd FILL
XFILL_0_OAI21X1_131 gnd vdd FILL
XDFFPOSX1_798 BUFX2_51/A CLKBUF1_37/Y OAI21X1_1090/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_974 gnd vdd FILL
XFILL_0_OAI21X1_186 gnd vdd FILL
XFILL_1_OAI21X1_346 gnd vdd FILL
XFILL_1_DFFPOSX1_996 gnd vdd FILL
XFILL_1_OAI21X1_368 gnd vdd FILL
XFILL_0_OAI21X1_197 gnd vdd FILL
XFILL_0_OAI21X1_175 gnd vdd FILL
XFILL_1_OAI21X1_357 gnd vdd FILL
XFILL_1_OAI21X1_379 gnd vdd FILL
XFILL_0_NAND3X1_17 gnd vdd FILL
XFILL_0_NAND3X1_39 gnd vdd FILL
XFILL_0_NAND3X1_28 gnd vdd FILL
XFILL_0_BUFX4_63 gnd vdd FILL
XFILL_0_BUFX4_52 gnd vdd FILL
XFILL_0_BUFX4_41 gnd vdd FILL
XFILL_0_BUFX4_30 gnd vdd FILL
XFILL_0_BUFX4_85 gnd vdd FILL
XFILL_0_BUFX4_96 gnd vdd FILL
XFILL_0_BUFX4_74 gnd vdd FILL
XFILL_1_NAND2X1_341 gnd vdd FILL
XFILL_0_NAND2X1_170 gnd vdd FILL
XFILL_1_NAND2X1_352 gnd vdd FILL
XFILL_0_DFFPOSX1_542 gnd vdd FILL
XFILL_1_BUFX4_127 gnd vdd FILL
XFILL_1_BUFX4_116 gnd vdd FILL
XFILL_1_BUFX4_105 gnd vdd FILL
XFILL_0_DFFPOSX1_520 gnd vdd FILL
XFILL_0_DFFPOSX1_531 gnd vdd FILL
XFILL_0_NAND2X1_192 gnd vdd FILL
XFILL_1_NAND2X1_374 gnd vdd FILL
XFILL_0_NAND2X1_181 gnd vdd FILL
XFILL_1_BUFX4_149 gnd vdd FILL
XFILL_1_BUFX4_138 gnd vdd FILL
XFILL_0_DFFPOSX1_575 gnd vdd FILL
XFILL_0_DFFPOSX1_564 gnd vdd FILL
XFILL_1_NAND2X1_385 gnd vdd FILL
XFILL_0_DFFPOSX1_553 gnd vdd FILL
XFILL_0_DFFPOSX1_586 gnd vdd FILL
XFILL_0_DFFPOSX1_597 gnd vdd FILL
XFILL_5_DFFPOSX1_190 gnd vdd FILL
XFILL_0_OR2X2_11 gnd vdd FILL
XNAND3X1_41 bundleAddress_i[32] bundleAddress_i[31] bundleAddress_i[30] gnd INVX1_192/A
+ vdd NAND3X1
XNAND3X1_30 AND2X2_7/Y NOR2X1_105/Y NOR2X1_30/Y gnd NOR2X1_114/B vdd NAND3X1
XFILL_1_OAI21X1_880 gnd vdd FILL
XFILL_1_OAI21X1_891 gnd vdd FILL
XNAND3X1_63 bundleAddress_i[50] INVX2_96/Y INVX2_108/A gnd INVX1_220/A vdd NAND3X1
XNAND3X1_52 bundleAddress_i[46] bundleAddress_i[45] INVX2_105/A gnd NOR2X1_185/B vdd
+ NAND3X1
XBUFX2_712 BUFX2_712/A gnd pid2_o[22] vdd BUFX2
XFILL_2_DFFPOSX1_603 gnd vdd FILL
XNOR2X1_30 NOR2X1_30/A NOR2X1_30/B gnd NOR2X1_30/Y vdd NOR2X1
XBUFX2_701 BUFX2_701/A gnd pid2_o[4] vdd BUFX2
XFILL_2_DFFPOSX1_614 gnd vdd FILL
XBUFX2_745 BUFX2_745/A gnd pid4_o[31] vdd BUFX2
XFILL_3_DFFPOSX1_50 gnd vdd FILL
XFILL_2_DFFPOSX1_636 gnd vdd FILL
XBUFX2_734 BUFX2_734/A gnd pid3_o[3] vdd BUFX2
XFILL_3_DFFPOSX1_61 gnd vdd FILL
XBUFX2_723 BUFX2_723/A gnd pid3_o[13] vdd BUFX2
XNOR2X1_52 NOR3X1_4/A NOR3X1_4/C gnd NOR2X1_52/Y vdd NOR2X1
XNOR2X1_63 OR2X2_5/Y OR2X2_10/B gnd NOR2X1_64/B vdd NOR2X1
XNOR2X1_41 NOR3X1_3/B NOR3X1_3/A gnd NOR2X1_41/Y vdd NOR2X1
XFILL_2_DFFPOSX1_647 gnd vdd FILL
XFILL_2_DFFPOSX1_625 gnd vdd FILL
XFILL_3_DFFPOSX1_94 gnd vdd FILL
XFILL_3_DFFPOSX1_83 gnd vdd FILL
XBUFX2_756 BUFX2_756/A gnd pid4_o[12] vdd BUFX2
XBUFX2_767 BUFX2_767/A gnd pid4_o[2] vdd BUFX2
XNOR2X1_96 NOR2X1_96/A NOR2X1_96/B gnd NOR2X1_96/Y vdd NOR2X1
XNOR2X1_85 bundleStartMajId_i[20] NOR2X1_85/B gnd NOR2X1_85/Y vdd NOR2X1
XFILL_3_DFFPOSX1_72 gnd vdd FILL
XNOR2X1_74 NOR2X1_74/A NOR2X1_74/B gnd NOR2X1_74/Y vdd NOR2X1
XBUFX2_778 BUFX2_778/A gnd tid1_o[62] vdd BUFX2
XBUFX2_789 BUFX2_789/A gnd tid1_o[61] vdd BUFX2
XFILL_2_DFFPOSX1_658 gnd vdd FILL
XFILL_2_DFFPOSX1_669 gnd vdd FILL
XFILL_0_NOR2X1_118 gnd vdd FILL
XFILL_0_NOR2X1_107 gnd vdd FILL
XFILL_0_NOR2X1_129 gnd vdd FILL
XFILL_30_3_1 gnd vdd FILL
XFILL_0_BUFX2_430 gnd vdd FILL
XFILL_0_BUFX2_441 gnd vdd FILL
XFILL_1_DFFPOSX1_204 gnd vdd FILL
XFILL_1_DFFPOSX1_237 gnd vdd FILL
XFILL_0_BUFX2_452 gnd vdd FILL
XFILL_1_DFFPOSX1_215 gnd vdd FILL
XFILL_1_DFFPOSX1_226 gnd vdd FILL
XFILL_0_BUFX2_463 gnd vdd FILL
XFILL_0_BUFX2_474 gnd vdd FILL
XFILL_1_DFFPOSX1_248 gnd vdd FILL
XFILL_1_DFFPOSX1_259 gnd vdd FILL
XFILL_0_BUFX2_485 gnd vdd FILL
XFILL_0_BUFX2_496 gnd vdd FILL
XNAND2X1_109 BUFX2_424/A BUFX4_319/Y gnd OAI21X1_365/C vdd NAND2X1
XNAND2X1_7 NAND2X1_7/A NAND2X1_7/B gnd OAI21X1_7/C vdd NAND2X1
XFILL_4_DFFPOSX1_719 gnd vdd FILL
XFILL_4_DFFPOSX1_708 gnd vdd FILL
XFILL_1_OAI21X1_29 gnd vdd FILL
XFILL_1_OAI21X1_18 gnd vdd FILL
XFILL_38_4_1 gnd vdd FILL
XFILL_0_NAND2X1_61 gnd vdd FILL
XNOR2X1_131 INVX2_66/Y OR2X2_16/A gnd XNOR2X1_57/A vdd NOR2X1
XNOR2X1_120 INVX2_39/Y NOR2X1_120/B gnd NOR2X1_120/Y vdd NOR2X1
XNOR2X1_142 INVX1_202/A NOR2X1_142/B gnd NOR2X1_142/Y vdd NOR2X1
XFILL_0_NAND2X1_72 gnd vdd FILL
XFILL_0_NAND2X1_83 gnd vdd FILL
XFILL_0_NAND2X1_50 gnd vdd FILL
XNOR2X1_164 bundleAddress_i[16] INVX2_102/Y gnd NOR2X1_164/Y vdd NOR2X1
XNOR2X1_175 INVX2_90/Y INVX1_181/Y gnd INVX1_199/A vdd NOR2X1
XNOR2X1_153 INVX4_40/Y NOR2X1_160/B gnd XNOR2X1_67/A vdd NOR2X1
XFILL_0_NAND2X1_94 gnd vdd FILL
XFILL_1_BUFX2_609 gnd vdd FILL
XNOR2X1_197 NOR3X1_18/A NOR3X1_18/C gnd INVX2_106/A vdd NOR2X1
XNOR2X1_186 OR2X2_18/Y NOR3X1_18/C gnd NOR2X1_187/B vdd NOR2X1
XFILL_27_18_1 gnd vdd FILL
XFILL_21_3_1 gnd vdd FILL
XOAI21X1_615 BUFX4_10/A BUFX4_345/Y BUFX2_561/A gnd OAI21X1_617/C vdd OAI21X1
XOAI21X1_604 INVX1_29/Y NOR2X1_89/B OAI21X1_604/C gnd OAI21X1_604/Y vdd OAI21X1
XFILL_3_DFFPOSX1_309 gnd vdd FILL
XOAI21X1_648 OAI21X1_648/A INVX1_4/Y BUFX4_305/Y gnd OAI21X1_649/B vdd OAI21X1
XOAI21X1_626 BUFX4_100/Y BUFX4_347/Y BUFX2_567/A gnd OAI21X1_628/C vdd OAI21X1
XOAI21X1_637 OAI21X1_637/A AOI21X1_20/Y OAI21X1_637/C gnd OAI21X1_637/Y vdd OAI21X1
XOAI21X1_659 bundleStartMajId_i[63] BUFX4_290/Y OAI21X1_659/C gnd OAI21X1_659/Y vdd
+ OAI21X1
XFILL_21_14_0 gnd vdd FILL
XDFFPOSX1_540 NOR2X1_96/A CLKBUF1_9/Y AOI21X1_23/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1170 gnd vdd FILL
XFILL_1_OAI21X1_110 gnd vdd FILL
XFILL_1_DFFPOSX1_760 gnd vdd FILL
XDFFPOSX1_551 BUFX2_608/A CLKBUF1_22/Y OAI21X1_669/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1181 gnd vdd FILL
XDFFPOSX1_573 BUFX2_603/A CLKBUF1_60/Y OAI21X1_733/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1192 gnd vdd FILL
XDFFPOSX1_562 BUFX2_591/A CLKBUF1_46/Y OAI21X1_700/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_121 gnd vdd FILL
XFILL_1_OAI21X1_132 gnd vdd FILL
XFILL_1_DFFPOSX1_771 gnd vdd FILL
XDFFPOSX1_595 BUFX2_627/A CLKBUF1_72/Y OAI21X1_796/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_143 gnd vdd FILL
XFILL_1_DFFPOSX1_793 gnd vdd FILL
XDFFPOSX1_584 BUFX2_615/A CLKBUF1_9/Y OAI21X1_763/Y gnd vdd DFFPOSX1
XNAND2X1_610 AND2X2_31/B INVX2_106/A gnd NOR3X1_16/C vdd NAND2X1
XNAND2X1_621 INVX2_103/A NOR2X1_172/Y gnd INVX1_214/A vdd NAND2X1
XFILL_1_DFFPOSX1_782 gnd vdd FILL
XNAND2X1_632 bundleAddress_i[37] INVX2_109/A gnd XNOR2X1_98/A vdd NAND2X1
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XNAND2X1_654 BUFX2_675/A BUFX4_367/Y gnd NAND2X1_654/Y vdd NAND2X1
XFILL_1_OAI21X1_165 gnd vdd FILL
XINVX1_11 NOR3X1_1/C gnd INVX1_11/Y vdd INVX1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XNAND2X1_643 bundleAddress_i[9] NOR2X1_229/Y gnd INVX1_226/A vdd NAND2X1
XFILL_1_INVX2_116 gnd vdd FILL
XFILL_1_OAI21X1_154 gnd vdd FILL
XFILL_1_OAI21X1_176 gnd vdd FILL
XNAND2X1_665 BUFX2_656/A BUFX4_380/Y gnd NAND2X1_665/Y vdd NAND2X1
XFILL_1_OAI21X1_187 gnd vdd FILL
XNAND2X1_676 BUFX2_668/A BUFX4_349/Y gnd NAND2X1_676/Y vdd NAND2X1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XFILL_1_OAI21X1_198 gnd vdd FILL
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XINVX1_66 INVX1_66/A gnd INVX1_66/Y vdd INVX1
XNAND2X1_687 BUFX2_708/A BUFX4_206/Y gnd NAND2X1_687/Y vdd NAND2X1
XINVX1_99 bundle_i[41] gnd INVX1_99/Y vdd INVX1
XNAND2X1_698 BUFX2_689/A BUFX4_231/Y gnd NAND2X1_698/Y vdd NAND2X1
XFILL_29_4_1 gnd vdd FILL
XINVX1_77 bundle_i[63] gnd INVX1_77/Y vdd INVX1
XINVX1_88 bundle_i[52] gnd INVX1_88/Y vdd INVX1
XFILL_4_4_1 gnd vdd FILL
XBUFX2_19 BUFX2_19/A gnd addr1_o[38] vdd BUFX2
XDFFPOSX1_7 BUFX2_704/A CLKBUF1_51/Y DFFPOSX1_7/D gnd vdd DFFPOSX1
XFILL_0_DFFPOSX1_350 gnd vdd FILL
XFILL_1_NAND2X1_193 gnd vdd FILL
XFILL_26_13_0 gnd vdd FILL
XFILL_12_3_1 gnd vdd FILL
XFILL_0_DFFPOSX1_361 gnd vdd FILL
XFILL_0_DFFPOSX1_372 gnd vdd FILL
XFILL_0_DFFPOSX1_383 gnd vdd FILL
XFILL_0_DFFPOSX1_394 gnd vdd FILL
XFILL_1_BUFX4_19 gnd vdd FILL
XFILL_3_DFFPOSX1_821 gnd vdd FILL
XFILL_3_DFFPOSX1_810 gnd vdd FILL
XFILL_3_DFFPOSX1_832 gnd vdd FILL
XFILL_3_DFFPOSX1_854 gnd vdd FILL
XFILL_3_DFFPOSX1_843 gnd vdd FILL
XFILL_3_DFFPOSX1_865 gnd vdd FILL
XFILL_3_DFFPOSX1_887 gnd vdd FILL
XFILL_3_DFFPOSX1_876 gnd vdd FILL
XFILL_3_DFFPOSX1_898 gnd vdd FILL
XFILL_7_18_1 gnd vdd FILL
XFILL_2_OAI21X1_881 gnd vdd FILL
XFILL_2_DFFPOSX1_422 gnd vdd FILL
XFILL_2_DFFPOSX1_400 gnd vdd FILL
XBUFX2_520 BUFX2_520/A gnd majID2_o[54] vdd BUFX2
XFILL_2_DFFPOSX1_411 gnd vdd FILL
XFILL_4_DFFPOSX1_51 gnd vdd FILL
XBUFX2_542 INVX1_28/A gnd majID3_o[35] vdd BUFX2
XFILL_4_DFFPOSX1_40 gnd vdd FILL
XFILL_1_14_0 gnd vdd FILL
XFILL_2_DFFPOSX1_433 gnd vdd FILL
XBUFX2_531 BUFX2_531/A gnd majID3_o[45] vdd BUFX2
XBUFX2_553 BUFX2_553/A gnd majID3_o[25] vdd BUFX2
XFILL_2_DFFPOSX1_455 gnd vdd FILL
XFILL_2_DFFPOSX1_444 gnd vdd FILL
XBUFX2_575 BUFX2_575/A gnd majID3_o[5] vdd BUFX2
XFILL_4_DFFPOSX1_84 gnd vdd FILL
XFILL_4_DFFPOSX1_62 gnd vdd FILL
XFILL_2_DFFPOSX1_477 gnd vdd FILL
XBUFX2_597 BUFX2_597/A gnd majID4_o[61] vdd BUFX2
XFILL_2_DFFPOSX1_499 gnd vdd FILL
XBUFX2_586 BUFX2_586/A gnd majID4_o[62] vdd BUFX2
XFILL_2_DFFPOSX1_466 gnd vdd FILL
XFILL_4_DFFPOSX1_73 gnd vdd FILL
XFILL_2_DFFPOSX1_488 gnd vdd FILL
XBUFX2_564 NOR2X1_89/A gnd majID3_o[15] vdd BUFX2
XFILL_4_DFFPOSX1_95 gnd vdd FILL
XFILL_5_DFFPOSX1_904 gnd vdd FILL
XFILL_5_DFFPOSX1_937 gnd vdd FILL
XFILL_5_DFFPOSX1_915 gnd vdd FILL
XFILL_5_DFFPOSX1_926 gnd vdd FILL
XFILL_5_DFFPOSX1_948 gnd vdd FILL
XFILL_5_DFFPOSX1_959 gnd vdd FILL
XFILL_0_BUFX2_271 gnd vdd FILL
XFILL_0_BUFX2_260 gnd vdd FILL
XFILL_0_AND2X2_6 gnd vdd FILL
XFILL_0_BUFX2_282 gnd vdd FILL
XFILL_0_BUFX2_293 gnd vdd FILL
XFILL_4_DFFPOSX1_516 gnd vdd FILL
XFILL_4_DFFPOSX1_527 gnd vdd FILL
XFILL_4_DFFPOSX1_505 gnd vdd FILL
XFILL_4_DFFPOSX1_538 gnd vdd FILL
XFILL_6_13_0 gnd vdd FILL
XFILL_4_DFFPOSX1_549 gnd vdd FILL
XFILL_10_11_1 gnd vdd FILL
XFILL_1_BUFX2_1007 gnd vdd FILL
XFILL_1_BUFX2_1029 gnd vdd FILL
XFILL_1_BUFX2_406 gnd vdd FILL
XFILL_0_NAND3X1_1 gnd vdd FILL
XFILL_1_BUFX2_439 gnd vdd FILL
XOAI21X1_423 NOR2X1_11/Y bundleStartMajId_i[47] BUFX4_245/Y gnd OAI21X1_424/B vdd
+ OAI21X1
XOAI21X1_412 XNOR2X1_1/Y BUFX4_215/Y OAI21X1_412/C gnd OAI21X1_412/Y vdd OAI21X1
XOAI21X1_401 INVX1_8/Y OAI21X1_401/B OAI21X1_401/C gnd OAI21X1_401/Y vdd OAI21X1
XFILL_3_DFFPOSX1_117 gnd vdd FILL
XOAI21X1_456 XNOR2X1_17/Y BUFX4_213/Y OAI21X1_456/C gnd OAI21X1_456/Y vdd OAI21X1
XOAI21X1_445 XNOR2X1_12/Y BUFX4_209/Y OAI21X1_445/C gnd OAI21X1_445/Y vdd OAI21X1
XFILL_1_CLKBUF1_19 gnd vdd FILL
XFILL_3_DFFPOSX1_106 gnd vdd FILL
XOAI21X1_434 XNOR2X1_9/Y BUFX4_194/Y OAI21X1_434/C gnd OAI21X1_434/Y vdd OAI21X1
XOAI21X1_478 XNOR2X1_21/Y BUFX4_200/Y OAI21X1_478/C gnd OAI21X1_478/Y vdd OAI21X1
XFILL_3_DFFPOSX1_139 gnd vdd FILL
XOAI21X1_489 OAI21X1_489/A BUFX4_213/Y OAI21X1_489/C gnd OAI21X1_489/Y vdd OAI21X1
XFILL_3_DFFPOSX1_128 gnd vdd FILL
XOAI21X1_467 XNOR2X1_20/Y BUFX4_199/Y OAI21X1_467/C gnd OAI21X1_467/Y vdd OAI21X1
XFILL_3_XNOR2X1_91 gnd vdd FILL
XDFFPOSX1_392 BUFX2_423/A CLKBUF1_19/Y OAI21X1_364/Y gnd vdd DFFPOSX1
XDFFPOSX1_381 BUFX2_411/A CLKBUF1_50/Y OAI21X1_353/Y gnd vdd DFFPOSX1
XDFFPOSX1_370 BUFX2_399/A CLKBUF1_6/Y OAI21X1_342/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_590 gnd vdd FILL
XNAND2X1_451 BUFX2_45/A BUFX4_342/Y gnd NAND2X1_451/Y vdd NAND2X1
XNAND2X1_462 BUFX2_58/A BUFX4_330/Y gnd NAND2X1_462/Y vdd NAND2X1
XNAND2X1_440 BUFX2_33/A BUFX4_384/Y gnd NAND2X1_440/Y vdd NAND2X1
XFILL_2_OAI21X1_155 gnd vdd FILL
XNAND2X1_473 BUFX2_110/A BUFX4_198/Y gnd NAND2X1_473/Y vdd NAND2X1
XNAND2X1_484 BUFX2_67/A BUFX4_231/Y gnd NAND2X1_484/Y vdd NAND2X1
XNAND2X1_495 NOR2X1_130/Y INVX1_186/Y gnd OR2X2_16/A vdd NAND2X1
XFILL_15_10_1 gnd vdd FILL
XFILL_2_OAI21X1_188 gnd vdd FILL
XFILL_0_INVX1_205 gnd vdd FILL
XFILL_0_INVX1_216 gnd vdd FILL
XFILL_0_INVX1_227 gnd vdd FILL
XFILL_0_DFFPOSX1_191 gnd vdd FILL
XFILL_0_DFFPOSX1_180 gnd vdd FILL
XFILL_0_OAI21X1_15 gnd vdd FILL
XFILL_1_BUFX2_973 gnd vdd FILL
XFILL_1_BUFX2_951 gnd vdd FILL
XFILL_0_OAI21X1_26 gnd vdd FILL
XFILL_0_OAI21X1_48 gnd vdd FILL
XFILL_1_BUFX2_962 gnd vdd FILL
XFILL_0_OAI21X1_37 gnd vdd FILL
XFILL_3_DFFPOSX1_640 gnd vdd FILL
XFILL_0_OAI21X1_59 gnd vdd FILL
XOAI21X1_1719 INVX2_121/Y BUFX4_302/Y OAI21X1_1719/C gnd DFFPOSX1_72/D vdd OAI21X1
XOAI21X1_1708 BUFX4_2/Y BUFX4_320/Y BUFX2_738/A gnd OAI21X1_1709/C vdd OAI21X1
XFILL_3_DFFPOSX1_662 gnd vdd FILL
XOAI21X1_990 BUFX4_136/Y BUFX4_81/Y BUFX2_388/A gnd OAI21X1_991/C vdd OAI21X1
XFILL_3_DFFPOSX1_651 gnd vdd FILL
XFILL_3_DFFPOSX1_673 gnd vdd FILL
XFILL_3_DFFPOSX1_695 gnd vdd FILL
XFILL_0_OAI21X1_708 gnd vdd FILL
XFILL_0_OAI21X1_719 gnd vdd FILL
XFILL_3_DFFPOSX1_684 gnd vdd FILL
XFILL_17_18_0 gnd vdd FILL
XFILL_33_11_1 gnd vdd FILL
XFILL_0_NAND2X1_736 gnd vdd FILL
XFILL_0_NAND2X1_703 gnd vdd FILL
XFILL_0_NAND2X1_714 gnd vdd FILL
XFILL_0_OAI21X1_1507 gnd vdd FILL
XFILL_2_DFFPOSX1_230 gnd vdd FILL
XFILL_0_NAND2X1_725 gnd vdd FILL
XBUFX2_350 BUFX2_350/A gnd instr3_o[0] vdd BUFX2
XFILL_35_2_1 gnd vdd FILL
XFILL_2_DFFPOSX1_252 gnd vdd FILL
XFILL_5_DFFPOSX1_30 gnd vdd FILL
XFILL_0_NAND2X1_769 gnd vdd FILL
XFILL_0_NAND2X1_758 gnd vdd FILL
XFILL_0_OAI21X1_1529 gnd vdd FILL
XFILL_0_OAI21X1_1518 gnd vdd FILL
XFILL_2_DFFPOSX1_263 gnd vdd FILL
XFILL_2_DFFPOSX1_274 gnd vdd FILL
XBUFX2_372 BUFX2_372/A gnd instr4_o[9] vdd BUFX2
XFILL_2_DFFPOSX1_241 gnd vdd FILL
XBUFX2_361 BUFX2_361/A gnd instr4_o[19] vdd BUFX2
XFILL_0_NAND2X1_747 gnd vdd FILL
XFILL_2_DFFPOSX1_296 gnd vdd FILL
XFILL_2_DFFPOSX1_285 gnd vdd FILL
XFILL_5_DFFPOSX1_52 gnd vdd FILL
XFILL_5_DFFPOSX1_63 gnd vdd FILL
XBUFX2_383 BUFX2_383/A gnd instr4_o[27] vdd BUFX2
XBUFX2_394 BUFX2_394/A gnd majID1_o[62] vdd BUFX2
XFILL_5_DFFPOSX1_41 gnd vdd FILL
XFILL_5_DFFPOSX1_701 gnd vdd FILL
XFILL_5_DFFPOSX1_85 gnd vdd FILL
XFILL_5_DFFPOSX1_96 gnd vdd FILL
XFILL_1_NOR3X1_11 gnd vdd FILL
XFILL_5_DFFPOSX1_712 gnd vdd FILL
XFILL_5_DFFPOSX1_74 gnd vdd FILL
XOAI21X1_61 INVX2_199/Y BUFX4_220/Y OAI21X1_61/C gnd OAI21X1_61/Y vdd OAI21X1
XOAI21X1_72 BUFX4_110/Y BUFX4_359/Y BUFX2_905/A gnd OAI21X1_73/C vdd OAI21X1
XFILL_5_DFFPOSX1_745 gnd vdd FILL
XFILL_5_DFFPOSX1_734 gnd vdd FILL
XFILL_5_DFFPOSX1_723 gnd vdd FILL
XOAI21X1_50 INVX2_188/Y BUFX4_228/Y OAI21X1_50/C gnd OAI21X1_50/Y vdd OAI21X1
XFILL_5_DFFPOSX1_756 gnd vdd FILL
XOAI21X1_94 BUFX4_11/A BUFX4_318/Y BUFX2_908/A gnd OAI21X1_95/C vdd OAI21X1
XFILL_5_DFFPOSX1_789 gnd vdd FILL
XFILL_5_DFFPOSX1_778 gnd vdd FILL
XFILL_5_DFFPOSX1_767 gnd vdd FILL
XOAI21X1_83 BUFX4_139/Y INVX2_151/Y OAI21X1_83/C gnd OAI21X1_83/Y vdd OAI21X1
XFILL_38_10_1 gnd vdd FILL
XFILL_4_DFFPOSX1_302 gnd vdd FILL
XFILL_0_DFFPOSX1_70 gnd vdd FILL
XFILL_4_DFFPOSX1_335 gnd vdd FILL
XFILL_4_DFFPOSX1_313 gnd vdd FILL
XFILL_4_DFFPOSX1_324 gnd vdd FILL
XFILL_2_DFFPOSX1_1005 gnd vdd FILL
XFILL_4_DFFPOSX1_346 gnd vdd FILL
XFILL_0_DFFPOSX1_92 gnd vdd FILL
XFILL_0_DFFPOSX1_81 gnd vdd FILL
XFILL_4_DFFPOSX1_357 gnd vdd FILL
XFILL_4_DFFPOSX1_368 gnd vdd FILL
XFILL_4_DFFPOSX1_379 gnd vdd FILL
XFILL_2_DFFPOSX1_1027 gnd vdd FILL
XFILL_2_DFFPOSX1_1016 gnd vdd FILL
XFILL_26_2_1 gnd vdd FILL
XFILL_1_2_1 gnd vdd FILL
XFILL_1_BUFX2_203 gnd vdd FILL
XFILL_1_BUFX2_214 gnd vdd FILL
XFILL_1_BUFX2_236 gnd vdd FILL
XOAI21X1_231 INVX2_161/Y BUFX4_290/Y OAI21X1_231/C gnd OAI21X1_231/Y vdd OAI21X1
XFILL_1_BUFX2_258 gnd vdd FILL
XFILL_1_BUFX2_247 gnd vdd FILL
XOAI21X1_220 BUFX4_124/Y BUFX4_40/Y BUFX2_971/A gnd OAI21X1_221/C vdd OAI21X1
XOAI21X1_253 INVX2_172/Y BUFX4_292/Y OAI21X1_253/C gnd OAI21X1_253/Y vdd OAI21X1
XOAI21X1_242 BUFX4_179/Y BUFX4_57/Y BUFX2_983/A gnd OAI21X1_243/C vdd OAI21X1
XOAI21X1_264 BUFX4_173/Y BUFX4_72/Y BUFX2_995/A gnd OAI21X1_265/C vdd OAI21X1
XOAI21X1_297 INVX2_194/Y BUFX4_292/Y OAI21X1_297/C gnd OAI21X1_297/Y vdd OAI21X1
XOAI21X1_275 INVX2_183/Y BUFX4_289/Y OAI21X1_275/C gnd OAI21X1_275/Y vdd OAI21X1
XOAI21X1_286 OR2X2_20/B BUFX4_27/Y BUFX2_1007/A gnd OAI21X1_287/C vdd OAI21X1
XAND2X2_31 INVX2_106/A AND2X2_31/B gnd AND2X2_31/Y vdd AND2X2
XAND2X2_20 AND2X2_20/A bundleStartMajId_i[50] gnd AND2X2_20/Y vdd AND2X2
XFILL_6_DFFPOSX1_429 gnd vdd FILL
XFILL_9_3_1 gnd vdd FILL
XNAND2X1_270 bundleStartMajId_i[56] bundleStartMajId_i[55] gnd NOR2X1_60/B vdd NAND2X1
XNAND2X1_292 bundleStartMajId_i[26] bundleStartMajId_i[25] gnd NOR3X1_5/B vdd NAND2X1
XNAND2X1_281 bundleStartMajId_i[40] bundleStartMajId_i[39] gnd NOR2X1_69/B vdd NAND2X1
XFILL_4_DFFPOSX1_880 gnd vdd FILL
XFILL_4_DFFPOSX1_891 gnd vdd FILL
XFILL_17_2_1 gnd vdd FILL
XFILL_0_INVX8_5 gnd vdd FILL
XFILL_0_BUFX4_300 gnd vdd FILL
XFILL_5_DFFPOSX1_1009 gnd vdd FILL
XFILL_0_BUFX4_322 gnd vdd FILL
XFILL_0_BUFX4_311 gnd vdd FILL
XFILL_1_BUFX2_770 gnd vdd FILL
XFILL_0_BUFX4_333 gnd vdd FILL
XOAI21X1_1505 OAI21X1_1505/A BUFX4_294/Y OAI21X1_1505/C gnd OAI21X1_1505/Y vdd OAI21X1
XFILL_1_OAI21X1_1725 gnd vdd FILL
XFILL_1_OAI21X1_1714 gnd vdd FILL
XFILL_0_BUFX4_366 gnd vdd FILL
XFILL_1_OAI21X1_1703 gnd vdd FILL
XOAI21X1_1527 NOR2X1_227/Y OAI21X1_1527/B OAI21X1_1527/C gnd OAI21X1_1527/Y vdd OAI21X1
XOAI21X1_1516 INVX2_110/Y NOR2X1_204/A BUFX4_284/Y gnd OAI21X1_1517/A vdd OAI21X1
XFILL_0_BUFX4_344 gnd vdd FILL
XOAI21X1_1538 BUFX4_160/Y BUFX4_66/A BUFX2_240/A gnd OAI21X1_1539/C vdd OAI21X1
XFILL_0_BUFX4_355 gnd vdd FILL
XFILL_0_BUFX4_377 gnd vdd FILL
XFILL_1_OAI21X1_1758 gnd vdd FILL
XFILL_1_OAI21X1_1736 gnd vdd FILL
XFILL_3_DFFPOSX1_470 gnd vdd FILL
XFILL_3_DFFPOSX1_481 gnd vdd FILL
XFILL_1_OAI21X1_1747 gnd vdd FILL
XFILL_0_BUFX4_388 gnd vdd FILL
XFILL_3_DFFPOSX1_492 gnd vdd FILL
XOAI21X1_1549 NAND2X1_644/Y BUFX4_303/Y OAI21X1_1549/C gnd OAI21X1_1549/Y vdd OAI21X1
XFILL_0_BUFX2_1015 gnd vdd FILL
XFILL_1_OAI21X1_1769 gnd vdd FILL
XFILL_1_OAI21X1_709 gnd vdd FILL
XFILL_0_OAI21X1_505 gnd vdd FILL
XFILL_0_OAI21X1_538 gnd vdd FILL
XFILL_0_OAI21X1_527 gnd vdd FILL
XFILL_0_OAI21X1_516 gnd vdd FILL
XFILL_0_BUFX2_1004 gnd vdd FILL
XFILL_0_OAI21X1_549 gnd vdd FILL
XFILL_6_DFFPOSX1_930 gnd vdd FILL
XFILL_0_BUFX2_1026 gnd vdd FILL
XFILL_6_DFFPOSX1_952 gnd vdd FILL
XFILL_6_DFFPOSX1_941 gnd vdd FILL
XFILL_0_CLKBUF1_16 gnd vdd FILL
XFILL_0_CLKBUF1_27 gnd vdd FILL
XFILL_0_NAND2X1_500 gnd vdd FILL
XFILL_0_CLKBUF1_49 gnd vdd FILL
XFILL_0_NAND2X1_511 gnd vdd FILL
XFILL_0_CLKBUF1_38 gnd vdd FILL
XFILL_0_NAND2X1_522 gnd vdd FILL
XFILL_1_NAND2X1_704 gnd vdd FILL
XFILL_1_NAND2X1_715 gnd vdd FILL
XFILL_0_NAND2X1_533 gnd vdd FILL
XFILL_0_NAND2X1_544 gnd vdd FILL
XFILL_0_OAI21X1_1315 gnd vdd FILL
XFILL_0_OAI21X1_1304 gnd vdd FILL
XFILL_1_NAND2X1_748 gnd vdd FILL
XFILL_1_NAND2X1_737 gnd vdd FILL
XFILL_0_NAND2X1_555 gnd vdd FILL
XFILL_0_OAI21X1_1337 gnd vdd FILL
XFILL_0_DFFPOSX1_905 gnd vdd FILL
XFILL_0_DFFPOSX1_916 gnd vdd FILL
XFILL_0_OAI21X1_1326 gnd vdd FILL
XFILL_0_NAND2X1_566 gnd vdd FILL
XFILL_0_OAI21X1_1348 gnd vdd FILL
XBUFX2_180 BUFX2_180/A gnd addr3_o[8] vdd BUFX2
XFILL_0_NAND2X1_577 gnd vdd FILL
XBUFX2_191 BUFX2_191/A gnd addr3_o[55] vdd BUFX2
XFILL_6_DFFPOSX1_20 gnd vdd FILL
XFILL_0_DFFPOSX1_949 gnd vdd FILL
XFILL_0_DFFPOSX1_938 gnd vdd FILL
XFILL_0_NAND2X1_588 gnd vdd FILL
XFILL_0_NAND2X1_599 gnd vdd FILL
XFILL_0_DFFPOSX1_927 gnd vdd FILL
XFILL_0_OAI21X1_1359 gnd vdd FILL
XFILL_6_DFFPOSX1_31 gnd vdd FILL
XFILL_6_DFFPOSX1_42 gnd vdd FILL
XFILL_5_DFFPOSX1_520 gnd vdd FILL
XFILL_5_DFFPOSX1_542 gnd vdd FILL
XFILL_20_9_0 gnd vdd FILL
XFILL_5_DFFPOSX1_531 gnd vdd FILL
XFILL_5_DFFPOSX1_553 gnd vdd FILL
XFILL_24_16_1 gnd vdd FILL
XFILL_5_DFFPOSX1_575 gnd vdd FILL
XFILL_5_DFFPOSX1_586 gnd vdd FILL
XFILL_5_DFFPOSX1_597 gnd vdd FILL
XFILL_5_DFFPOSX1_564 gnd vdd FILL
XFILL_1_BUFX4_8 gnd vdd FILL
XFILL_1_AOI21X1_4 gnd vdd FILL
XCLKBUF1_40 BUFX4_89/Y gnd CLKBUF1_40/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_110 gnd vdd FILL
XCLKBUF1_51 BUFX4_88/Y gnd CLKBUF1_51/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_121 gnd vdd FILL
XFILL_4_DFFPOSX1_154 gnd vdd FILL
XFILL_4_DFFPOSX1_143 gnd vdd FILL
XFILL_1_DFFPOSX1_60 gnd vdd FILL
XCLKBUF1_73 BUFX4_83/Y gnd CLKBUF1_73/Y vdd CLKBUF1
XCLKBUF1_84 BUFX4_83/Y gnd CLKBUF1_84/Y vdd CLKBUF1
XCLKBUF1_62 BUFX4_88/Y gnd CLKBUF1_62/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_132 gnd vdd FILL
XFILL_4_DFFPOSX1_176 gnd vdd FILL
XFILL_1_DFFPOSX1_82 gnd vdd FILL
XFILL_4_DFFPOSX1_187 gnd vdd FILL
XCLKBUF1_95 BUFX4_92/Y gnd CLKBUF1_95/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_93 gnd vdd FILL
XFILL_1_DFFPOSX1_71 gnd vdd FILL
XFILL_4_DFFPOSX1_165 gnd vdd FILL
XFILL_4_DFFPOSX1_198 gnd vdd FILL
XFILL_29_15_1 gnd vdd FILL
XFILL_11_9_0 gnd vdd FILL
XFILL_0_BUFX2_804 gnd vdd FILL
XFILL_0_BUFX2_815 gnd vdd FILL
XFILL_23_11_0 gnd vdd FILL
XFILL_0_BUFX2_826 gnd vdd FILL
XFILL_0_BUFX2_848 gnd vdd FILL
XINVX1_125 bundle_i[79] gnd INVX1_125/Y vdd INVX1
XINVX1_103 bundle_i[37] gnd INVX1_103/Y vdd INVX1
XINVX1_114 bundle_i[90] gnd INVX1_114/Y vdd INVX1
XFILL_0_BUFX2_837 gnd vdd FILL
XINVX1_147 bundle_i[121] gnd INVX1_147/Y vdd INVX1
XFILL_0_BUFX2_859 gnd vdd FILL
XINVX1_158 bundle_i[110] gnd INVX1_158/Y vdd INVX1
XINVX1_136 bundle_i[68] gnd INVX1_136/Y vdd INVX1
XFILL_3_XNOR2X1_2 gnd vdd FILL
XINVX1_169 bundle_i[99] gnd INVX1_169/Y vdd INVX1
XFILL_6_DFFPOSX1_215 gnd vdd FILL
XFILL_6_DFFPOSX1_226 gnd vdd FILL
XFILL_6_DFFPOSX1_204 gnd vdd FILL
XFILL_6_DFFPOSX1_237 gnd vdd FILL
XFILL_0_INVX2_35 gnd vdd FILL
XFILL_0_INVX2_46 gnd vdd FILL
XFILL_0_INVX2_24 gnd vdd FILL
XFILL_0_INVX2_13 gnd vdd FILL
XFILL_0_INVX2_68 gnd vdd FILL
XFILL_0_INVX2_57 gnd vdd FILL
XFILL_0_INVX2_79 gnd vdd FILL
XFILL_4_16_1 gnd vdd FILL
XFILL_0_CLKBUF1_3 gnd vdd FILL
XFILL_32_0_1 gnd vdd FILL
XFILL_28_10_0 gnd vdd FILL
XFILL_4_CLKBUF1_2 gnd vdd FILL
XOAI21X1_1302 BUFX4_11/Y BUFX4_381/Y BUFX2_157/A gnd OAI21X1_1303/C vdd OAI21X1
XFILL_0_BUFX4_141 gnd vdd FILL
XFILL_0_BUFX4_130 gnd vdd FILL
XOAI21X1_1313 NOR2X1_199/Y NAND2X1_611/Y OAI21X1_1313/C gnd OAI21X1_1313/Y vdd OAI21X1
XFILL_1_OAI21X1_1500 gnd vdd FILL
XFILL_1_OAI21X1_1533 gnd vdd FILL
XDFFPOSX1_903 BUFX2_154/A CLKBUF1_21/Y OAI21X1_1294/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1522 gnd vdd FILL
XOAI21X1_1335 AOI21X1_52/Y OAI21X1_1335/B OAI21X1_1335/C gnd OAI21X1_1335/Y vdd OAI21X1
XFILL_0_BUFX4_174 gnd vdd FILL
XDFFPOSX1_914 INVX1_209/A CLKBUF1_85/Y OAI21X1_1324/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1511 gnd vdd FILL
XOAI21X1_1346 INVX2_106/Y NOR3X1_18/B MUX2X1_2/S gnd OAI21X1_1347/B vdd OAI21X1
XOAI21X1_1324 INVX1_209/Y BUFX4_308/Y OAI21X1_1324/C gnd OAI21X1_1324/Y vdd OAI21X1
XFILL_0_BUFX4_185 gnd vdd FILL
XFILL_0_BUFX4_152 gnd vdd FILL
XFILL_0_BUFX4_163 gnd vdd FILL
XFILL_1_BUFX2_63 gnd vdd FILL
XFILL_0_OAI21X1_313 gnd vdd FILL
XDFFPOSX1_936 BUFX2_193/A CLKBUF1_57/Y OAI21X1_1385/Y gnd vdd DFFPOSX1
XDFFPOSX1_947 BUFX2_196/A CLKBUF1_70/Y OAI21X1_1417/Y gnd vdd DFFPOSX1
XFILL_1_BUFX2_41 gnd vdd FILL
XOAI21X1_1379 BUFX4_103/Y BUFX4_360/Y BUFX2_188/A gnd OAI21X1_1381/C vdd OAI21X1
XFILL_1_OAI21X1_1566 gnd vdd FILL
XOAI21X1_1368 INVX1_215/A INVX1_197/A INVX2_89/Y gnd OAI21X1_1369/C vdd OAI21X1
XDFFPOSX1_925 BUFX2_178/A CLKBUF1_36/Y OAI21X1_1354/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_302 gnd vdd FILL
XFILL_1_BUFX2_52 gnd vdd FILL
XOAI21X1_1357 AOI21X1_56/Y OAI21X1_1357/B OAI21X1_1357/C gnd OAI21X1_1357/Y vdd OAI21X1
XFILL_1_OAI21X1_1544 gnd vdd FILL
XFILL_1_OAI21X1_1555 gnd vdd FILL
XFILL_0_BUFX4_196 gnd vdd FILL
XFILL_1_OAI21X1_1588 gnd vdd FILL
XFILL_0_OAI21X1_346 gnd vdd FILL
XDFFPOSX1_969 BUFX2_220/A CLKBUF1_68/Y OAI21X1_1482/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1599 gnd vdd FILL
XFILL_1_OAI21X1_1577 gnd vdd FILL
XDFFPOSX1_958 BUFX2_208/A CLKBUF1_34/Y OAI21X1_1451/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_324 gnd vdd FILL
XFILL_1_OAI21X1_506 gnd vdd FILL
XFILL_1_BUFX2_96 gnd vdd FILL
XFILL_0_OAI21X1_335 gnd vdd FILL
XFILL_1_OAI21X1_517 gnd vdd FILL
XFILL_0_OAI21X1_379 gnd vdd FILL
XFILL_0_OAI21X1_368 gnd vdd FILL
XFILL_0_OAI21X1_357 gnd vdd FILL
XFILL_1_OAI21X1_539 gnd vdd FILL
XFILL_1_OAI21X1_528 gnd vdd FILL
XFILL_9_15_1 gnd vdd FILL
XFILL_6_DFFPOSX1_793 gnd vdd FILL
XFILL_1_OAI21X1_7 gnd vdd FILL
XFILL_3_11_0 gnd vdd FILL
XFILL_0_NAND2X1_352 gnd vdd FILL
XFILL_0_OAI21X1_1123 gnd vdd FILL
XFILL_0_OAI21X1_1112 gnd vdd FILL
XFILL_1_NAND2X1_501 gnd vdd FILL
XFILL_0_OAI21X1_1101 gnd vdd FILL
XFILL_1_NAND2X1_523 gnd vdd FILL
XFILL_0_NAND2X1_330 gnd vdd FILL
XFILL_0_NAND2X1_341 gnd vdd FILL
XFILL_0_DFFPOSX1_713 gnd vdd FILL
XFILL_0_OAI21X1_1156 gnd vdd FILL
XFILL_0_OAI21X1_1145 gnd vdd FILL
XFILL_1_NAND2X1_556 gnd vdd FILL
XFILL_1_BUFX4_309 gnd vdd FILL
XFILL_0_DFFPOSX1_702 gnd vdd FILL
XFILL_1_NAND2X1_534 gnd vdd FILL
XFILL_0_NAND2X1_374 gnd vdd FILL
XFILL_0_NAND2X1_385 gnd vdd FILL
XFILL_0_NAND2X1_363 gnd vdd FILL
XFILL_0_DFFPOSX1_724 gnd vdd FILL
XFILL_1_NAND2X1_545 gnd vdd FILL
XFILL_0_OAI21X1_1134 gnd vdd FILL
XFILL_0_DFFPOSX1_746 gnd vdd FILL
XFILL_0_DFFPOSX1_757 gnd vdd FILL
XFILL_0_OAI21X1_1178 gnd vdd FILL
XFILL_23_0_1 gnd vdd FILL
XFILL_0_DFFPOSX1_735 gnd vdd FILL
XFILL_1_NAND2X1_589 gnd vdd FILL
XFILL_1_NAND2X1_578 gnd vdd FILL
XFILL_0_NAND2X1_396 gnd vdd FILL
XFILL_0_OAI21X1_1167 gnd vdd FILL
XFILL_0_OAI21X1_1189 gnd vdd FILL
XFILL_0_DFFPOSX1_779 gnd vdd FILL
XFILL_0_DFFPOSX1_768 gnd vdd FILL
XFILL_5_DFFPOSX1_350 gnd vdd FILL
XFILL_5_DFFPOSX1_361 gnd vdd FILL
XFILL_5_DFFPOSX1_372 gnd vdd FILL
XFILL_5_DFFPOSX1_394 gnd vdd FILL
XFILL_5_DFFPOSX1_383 gnd vdd FILL
XINVX4_11 bundleStartMajId_i[38] gnd INVX4_11/Y vdd INVX4
XFILL_1_NAND2X1_10 gnd vdd FILL
XFILL_1_NAND2X1_21 gnd vdd FILL
XINVX4_33 bundleAddress_i[52] gnd INVX4_33/Y vdd INVX4
XFILL_1_NAND2X1_65 gnd vdd FILL
XINVX4_22 bundleStartMajId_i[15] gnd INVX4_22/Y vdd INVX4
XFILL_1_NAND2X1_43 gnd vdd FILL
XINVX4_44 bundleAddress_i[13] gnd INVX4_44/Y vdd INVX4
XFILL_1_NAND2X1_98 gnd vdd FILL
XFILL_1_NAND2X1_76 gnd vdd FILL
XFILL_1_NAND2X1_87 gnd vdd FILL
XFILL_1_BUFX2_5 gnd vdd FILL
XFILL_0_OAI21X1_880 gnd vdd FILL
XFILL_0_OAI21X1_891 gnd vdd FILL
XFILL_8_10_0 gnd vdd FILL
XFILL_6_1_1 gnd vdd FILL
XFILL_2_DFFPOSX1_50 gnd vdd FILL
XBUFX2_916 BUFX2_916/A gnd tid3_o[44] vdd BUFX2
XBUFX2_905 BUFX2_905/A gnd tid3_o[63] vdd BUFX2
XFILL_2_DFFPOSX1_818 gnd vdd FILL
XFILL_2_DFFPOSX1_61 gnd vdd FILL
XFILL_2_DFFPOSX1_807 gnd vdd FILL
XFILL_2_DFFPOSX1_72 gnd vdd FILL
XBUFX2_938 BUFX2_938/A gnd tid3_o[24] vdd BUFX2
XBUFX2_927 BUFX2_927/A gnd tid3_o[34] vdd BUFX2
XFILL_2_DFFPOSX1_829 gnd vdd FILL
XFILL_2_DFFPOSX1_94 gnd vdd FILL
XFILL_2_DFFPOSX1_83 gnd vdd FILL
XBUFX2_949 BUFX2_949/A gnd tid3_o[14] vdd BUFX2
XFILL_14_0_1 gnd vdd FILL
XFILL_0_OAI21X1_1690 gnd vdd FILL
XFILL_0_BUFX2_623 gnd vdd FILL
XFILL_0_BUFX2_612 gnd vdd FILL
XFILL_0_BUFX2_601 gnd vdd FILL
XFILL_0_BUFX2_656 gnd vdd FILL
XFILL_1_DFFPOSX1_408 gnd vdd FILL
XFILL_1_DFFPOSX1_419 gnd vdd FILL
XFILL_0_BUFX2_634 gnd vdd FILL
XFILL_0_BUFX2_645 gnd vdd FILL
XFILL_0_BUFX2_667 gnd vdd FILL
XFILL_0_BUFX2_678 gnd vdd FILL
XFILL_0_BUFX2_689 gnd vdd FILL
XBUFX4_220 BUFX4_26/Y gnd BUFX4_220/Y vdd BUFX4
XFILL_14_16_0 gnd vdd FILL
XBUFX4_231 BUFX4_25/Y gnd BUFX4_231/Y vdd BUFX4
XBUFX4_253 INVX8_5/Y gnd BUFX4_95/A vdd BUFX4
XBUFX4_242 INVX8_1/Y gnd BUFX4_242/Y vdd BUFX4
XBUFX4_264 enable_i gnd BUFX4_264/Y vdd BUFX4
XFILL_0_INVX2_130 gnd vdd FILL
XFILL_2_OAI21X1_1762 gnd vdd FILL
XFILL_0_INVX2_152 gnd vdd FILL
XBUFX4_297 BUFX4_303/A gnd BUFX4_297/Y vdd BUFX4
XBUFX4_286 INVX8_2/Y gnd BUFX4_286/Y vdd BUFX4
XBUFX4_275 INVX8_7/Y gnd BUFX4_79/A vdd BUFX4
XFILL_0_INVX2_141 gnd vdd FILL
XFILL_2_OAI21X1_1784 gnd vdd FILL
XFILL_0_INVX2_163 gnd vdd FILL
XFILL_34_8_0 gnd vdd FILL
XFILL_0_INVX2_185 gnd vdd FILL
XFILL_0_INVX2_174 gnd vdd FILL
XFILL_0_INVX2_196 gnd vdd FILL
XFILL_25_1 gnd vdd FILL
XOAI21X1_808 BUFX4_156/Y BUFX4_48/Y BUFX2_632/A gnd OAI21X1_809/C vdd OAI21X1
XOAI21X1_819 BUFX4_133/Y BUFX4_31/Y BUFX2_636/A gnd OAI21X1_821/C vdd OAI21X1
XOAI21X1_1110 INVX4_47/Y INVX4_32/Y OAI21X1_1110/C gnd OAI21X1_1111/A vdd OAI21X1
XOAI21X1_1121 OAI21X1_1121/A INVX2_95/A NAND2X1_484/Y gnd OAI21X1_1121/Y vdd OAI21X1
XDFFPOSX1_700 BUFX2_338/A CLKBUF1_25/Y OAI21X1_949/Y gnd vdd DFFPOSX1
XDFFPOSX1_711 BUFX2_350/A CLKBUF1_95/Y OAI21X1_971/Y gnd vdd DFFPOSX1
XOAI21X1_1143 XNOR2X1_62/Y BUFX4_202/Y NAND2X1_515/Y gnd OAI21X1_1143/Y vdd OAI21X1
XDFFPOSX1_722 BUFX2_359/A CLKBUF1_61/Y OAI21X1_993/Y gnd vdd DFFPOSX1
XOAI21X1_1154 NOR2X1_149/Y OAI21X1_1154/B NAND2X1_531/Y gnd OAI21X1_1154/Y vdd OAI21X1
XFILL_1_OAI21X1_1341 gnd vdd FILL
XFILL_1_OAI21X1_1330 gnd vdd FILL
XOAI21X1_1132 INVX1_188/A bundleAddress_i[45] BUFX4_239/Y gnd OAI21X1_1133/B vdd OAI21X1
XOAI21X1_1165 INVX1_193/A INVX8_3/Y INVX2_79/Y gnd NAND2X1_547/B vdd OAI21X1
XFILL_0_OAI21X1_121 gnd vdd FILL
XDFFPOSX1_755 BUFX2_4/A CLKBUF1_65/Y OAI21X1_1047/Y gnd vdd DFFPOSX1
XDFFPOSX1_744 BUFX2_1/A CLKBUF1_17/Y OAI21X1_1036/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_942 gnd vdd FILL
XFILL_0_OAI21X1_110 gnd vdd FILL
XFILL_1_DFFPOSX1_920 gnd vdd FILL
XOAI21X1_1176 NOR2X1_164/Y OAI21X1_1176/B NAND2X1_559/Y gnd OAI21X1_1176/Y vdd OAI21X1
XFILL_1_OAI21X1_1374 gnd vdd FILL
XFILL_1_DFFPOSX1_931 gnd vdd FILL
XOAI21X1_1198 NAND3X1_51/Y INVX2_90/Y BUFX4_243/Y gnd OAI21X1_1199/A vdd OAI21X1
XFILL_1_OAI21X1_1352 gnd vdd FILL
XDFFPOSX1_733 BUFX2_371/A CLKBUF1_77/Y OAI21X1_1015/Y gnd vdd DFFPOSX1
XOAI21X1_1187 NOR3X1_13/Y OAI21X1_1187/B NAND2X1_573/Y gnd OAI21X1_1187/Y vdd OAI21X1
XDFFPOSX1_766 BUFX2_16/A CLKBUF1_51/Y OAI21X1_1058/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1363 gnd vdd FILL
XFILL_1_OAI21X1_1385 gnd vdd FILL
XFILL_0_OAI21X1_132 gnd vdd FILL
XFILL_1_OAI21X1_1396 gnd vdd FILL
XFILL_1_DFFPOSX1_953 gnd vdd FILL
XFILL_1_DFFPOSX1_964 gnd vdd FILL
XDFFPOSX1_788 BUFX2_40/A CLKBUF1_21/Y OAI21X1_1080/Y gnd vdd DFFPOSX1
XDFFPOSX1_777 BUFX2_28/A CLKBUF1_89/Y OAI21X1_1069/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_314 gnd vdd FILL
XFILL_0_OAI21X1_143 gnd vdd FILL
XFILL_1_OAI21X1_303 gnd vdd FILL
XFILL_1_OAI21X1_325 gnd vdd FILL
XDFFPOSX1_799 BUFX2_52/A CLKBUF1_20/Y OAI21X1_1091/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_154 gnd vdd FILL
XFILL_1_DFFPOSX1_975 gnd vdd FILL
XFILL_0_OAI21X1_187 gnd vdd FILL
XFILL_1_OAI21X1_347 gnd vdd FILL
XFILL_1_DFFPOSX1_997 gnd vdd FILL
XFILL_19_15_0 gnd vdd FILL
XFILL_1_OAI21X1_369 gnd vdd FILL
XFILL_0_OAI21X1_165 gnd vdd FILL
XFILL_1_OAI21X1_358 gnd vdd FILL
XFILL_1_OAI21X1_336 gnd vdd FILL
XFILL_1_DFFPOSX1_986 gnd vdd FILL
XFILL_0_OAI21X1_176 gnd vdd FILL
XFILL_6_DFFPOSX1_590 gnd vdd FILL
XFILL_0_OAI21X1_198 gnd vdd FILL
XFILL_32_17_0 gnd vdd FILL
XFILL_0_NAND3X1_18 gnd vdd FILL
XFILL_0_NAND3X1_29 gnd vdd FILL
XFILL_0_BUFX4_20 gnd vdd FILL
XFILL_0_BUFX4_42 gnd vdd FILL
XFILL_0_BUFX4_53 gnd vdd FILL
XFILL_0_BUFX4_31 gnd vdd FILL
XFILL_0_BUFX4_75 gnd vdd FILL
XFILL_0_BUFX4_64 gnd vdd FILL
XFILL_25_8_0 gnd vdd FILL
XFILL_1_NAND2X1_331 gnd vdd FILL
XFILL_0_BUFX4_86 gnd vdd FILL
XFILL_1_NAND2X1_320 gnd vdd FILL
XFILL_0_8_0 gnd vdd FILL
XFILL_0_NAND2X1_160 gnd vdd FILL
XFILL_0_BUFX4_97 gnd vdd FILL
XFILL_1_BUFX4_128 gnd vdd FILL
XFILL_1_BUFX4_106 gnd vdd FILL
XFILL_0_DFFPOSX1_510 gnd vdd FILL
XFILL_1_BUFX4_117 gnd vdd FILL
XFILL_1_NAND2X1_364 gnd vdd FILL
XFILL_0_DFFPOSX1_521 gnd vdd FILL
XFILL_0_DFFPOSX1_532 gnd vdd FILL
XFILL_0_NAND2X1_171 gnd vdd FILL
XFILL_0_NAND2X1_182 gnd vdd FILL
XFILL_1_NAND2X1_353 gnd vdd FILL
XFILL_0_NAND2X1_193 gnd vdd FILL
XFILL_1_NAND2X1_386 gnd vdd FILL
XFILL_0_DFFPOSX1_543 gnd vdd FILL
XFILL_0_DFFPOSX1_576 gnd vdd FILL
XFILL_0_DFFPOSX1_565 gnd vdd FILL
XFILL_1_NAND2X1_397 gnd vdd FILL
XFILL_1_BUFX4_139 gnd vdd FILL
XFILL_0_DFFPOSX1_554 gnd vdd FILL
XFILL_0_DFFPOSX1_598 gnd vdd FILL
XFILL_0_DFFPOSX1_587 gnd vdd FILL
XFILL_5_DFFPOSX1_180 gnd vdd FILL
XFILL_5_DFFPOSX1_191 gnd vdd FILL
XFILL_0_OR2X2_12 gnd vdd FILL
XFILL_37_16_0 gnd vdd FILL
XFILL_8_9_0 gnd vdd FILL
XFILL_1_OAI21X1_881 gnd vdd FILL
XFILL_1_OAI21X1_870 gnd vdd FILL
XNAND3X1_20 bundleStartMajId_i[24] INVX1_30/Y NOR2X1_80/Y gnd NAND3X1_20/Y vdd NAND3X1
XNAND3X1_31 bundleStartMajId_i[18] INVX2_49/A INVX4_31/A gnd AND2X2_22/A vdd NAND3X1
XFILL_1_OAI21X1_892 gnd vdd FILL
XNAND3X1_64 INVX2_98/Y AND2X2_28/A INVX2_109/A gnd XNOR2X1_99/A vdd NAND3X1
XNAND3X1_42 AND2X2_28/A INVX2_98/Y INVX1_192/Y gnd NOR2X1_152/B vdd NAND3X1
XNAND3X1_53 bundleAddress_i[39] INVX1_202/Y NOR2X1_187/B gnd AND2X2_27/A vdd NAND3X1
XBUFX2_702 BUFX2_702/A gnd pid2_o[3] vdd BUFX2
XFILL_2_DFFPOSX1_604 gnd vdd FILL
XNOR2X1_20 INVX4_13/Y INVX4_14/Y gnd INVX1_13/A vdd NOR2X1
XBUFX2_746 BUFX2_746/A gnd pid4_o[30] vdd BUFX2
XBUFX2_713 BUFX2_713/A gnd pid3_o[31] vdd BUFX2
XFILL_3_DFFPOSX1_51 gnd vdd FILL
XFILL_3_DFFPOSX1_62 gnd vdd FILL
XFILL_2_DFFPOSX1_615 gnd vdd FILL
XNOR2X1_53 INVX2_37/Y INVX4_25/Y gnd NOR2X1_53/Y vdd NOR2X1
XFILL_3_DFFPOSX1_40 gnd vdd FILL
XNOR2X1_42 NOR2X1_42/A NOR2X1_42/B gnd NOR2X1_42/Y vdd NOR2X1
XBUFX2_724 BUFX2_724/A gnd pid3_o[12] vdd BUFX2
XNOR2X1_64 bundleStartMajId_i[43] NOR2X1_64/B gnd NOR2X1_64/Y vdd NOR2X1
XFILL_2_DFFPOSX1_648 gnd vdd FILL
XNOR2X1_31 OR2X2_8/A NOR2X1_31/B gnd AND2X2_7/A vdd NOR2X1
XBUFX2_735 BUFX2_735/A gnd pid3_o[2] vdd BUFX2
XFILL_2_DFFPOSX1_626 gnd vdd FILL
XFILL_2_DFFPOSX1_637 gnd vdd FILL
XFILL_3_DFFPOSX1_84 gnd vdd FILL
XBUFX2_757 BUFX2_757/A gnd pid4_o[29] vdd BUFX2
XFILL_3_DFFPOSX1_95 gnd vdd FILL
XBUFX2_768 BUFX2_768/A gnd pid4_o[28] vdd BUFX2
XNOR2X1_97 OR2X2_13/Y NOR2X1_97/B gnd NOR2X1_97/Y vdd NOR2X1
XFILL_16_8_0 gnd vdd FILL
XNOR2X1_86 INVX1_32/A NOR3X1_3/B gnd INVX2_49/A vdd NOR2X1
XNOR2X1_75 OR2X2_10/B OR2X2_10/A gnd NOR2X1_75/Y vdd NOR2X1
XFILL_2_DFFPOSX1_659 gnd vdd FILL
XBUFX2_779 BUFX2_779/A gnd tid1_o[53] vdd BUFX2
XFILL_3_DFFPOSX1_73 gnd vdd FILL
XFILL_0_NOR2X1_119 gnd vdd FILL
XFILL_0_NOR2X1_108 gnd vdd FILL
XFILL_0_BUFX2_431 gnd vdd FILL
XFILL_1_DFFPOSX1_205 gnd vdd FILL
XFILL_0_BUFX2_420 gnd vdd FILL
XFILL_0_BUFX2_475 gnd vdd FILL
XFILL_1_DFFPOSX1_238 gnd vdd FILL
XFILL_0_BUFX2_442 gnd vdd FILL
XFILL_0_BUFX2_453 gnd vdd FILL
XFILL_1_DFFPOSX1_216 gnd vdd FILL
XFILL_0_BUFX2_464 gnd vdd FILL
XFILL_1_DFFPOSX1_227 gnd vdd FILL
XFILL_1_DFFPOSX1_249 gnd vdd FILL
XFILL_0_BUFX2_486 gnd vdd FILL
XFILL_0_BUFX2_497 gnd vdd FILL
XFILL_4_DFFPOSX1_709 gnd vdd FILL
XFILL_1_OAI21X1_19 gnd vdd FILL
XNAND2X1_8 NAND2X1_8/A OAI21X1_8/B gnd OAI21X1_8/C vdd NAND2X1
XFILL_0_NAND2X1_40 gnd vdd FILL
XFILL_0_NAND2X1_62 gnd vdd FILL
XFILL_2_OAI21X1_1581 gnd vdd FILL
XFILL_0_NAND2X1_51 gnd vdd FILL
XNOR2X1_121 INVX4_32/Y INVX2_56/Y gnd INVX1_184/A vdd NOR2X1
XNOR2X1_132 INVX4_34/Y OR2X2_16/Y gnd XNOR2X1_59/A vdd NOR2X1
XFILL_2_OAI21X1_1570 gnd vdd FILL
XFILL_0_NAND2X1_73 gnd vdd FILL
XNOR2X1_110 INVX2_43/Y OR2X2_15/A gnd NOR2X1_110/Y vdd NOR2X1
XNOR2X1_143 INVX2_71/Y INVX1_190/A gnd XNOR2X1_64/A vdd NOR2X1
XNOR2X1_165 INVX1_195/A NOR2X1_165/B gnd NOR2X1_165/Y vdd NOR2X1
XNOR2X1_176 INVX2_91/Y NOR2X1_176/B gnd INVX4_49/A vdd NOR2X1
XNOR2X1_154 NOR2X1_154/A NOR2X1_160/B gnd XNOR2X1_68/A vdd NOR2X1
XFILL_0_NAND2X1_84 gnd vdd FILL
XFILL_0_NAND2X1_95 gnd vdd FILL
XNOR2X1_187 bundleAddress_i[41] NOR2X1_187/B gnd NOR2X1_187/Y vdd NOR2X1
XNOR2X1_198 INVX4_41/Y XNOR2X1_83/A gnd NOR2X1_199/B vdd NOR2X1
XOAI21X1_605 BUFX4_2/A BUFX4_323/Y BUFX2_557/A gnd OAI21X1_606/C vdd OAI21X1
XOAI21X1_627 NOR2X1_97/B INVX2_51/Y NOR2X1_96/B gnd OAI21X1_628/B vdd OAI21X1
XOAI21X1_638 BUFX4_2/A BUFX4_325/Y BUFX2_572/A gnd OAI21X1_640/C vdd OAI21X1
XOAI21X1_616 INVX2_50/Y INVX2_30/Y NOR2X1_89/B gnd OAI21X1_617/A vdd OAI21X1
XOAI21X1_649 NOR2X1_98/Y OAI21X1_649/B OAI21X1_649/C gnd OAI21X1_649/Y vdd OAI21X1
XFILL_21_14_1 gnd vdd FILL
XDFFPOSX1_541 BUFX2_574/A CLKBUF1_72/Y OAI21X1_643/Y gnd vdd DFFPOSX1
XDFFPOSX1_530 BUFX2_562/A CLKBUF1_90/Y OAI21X1_620/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_100 gnd vdd FILL
XFILL_1_DFFPOSX1_750 gnd vdd FILL
XFILL_1_OAI21X1_1171 gnd vdd FILL
XDFFPOSX1_563 BUFX2_592/A CLKBUF1_91/Y OAI21X1_703/Y gnd vdd DFFPOSX1
XDFFPOSX1_574 BUFX2_604/A CLKBUF1_63/Y OAI21X1_736/Y gnd vdd DFFPOSX1
XDFFPOSX1_552 BUFX2_619/A CLKBUF1_94/Y OAI21X1_671/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1182 gnd vdd FILL
XFILL_1_OAI21X1_1193 gnd vdd FILL
XFILL_1_OAI21X1_1160 gnd vdd FILL
XFILL_1_OAI21X1_133 gnd vdd FILL
XFILL_1_DFFPOSX1_761 gnd vdd FILL
XFILL_1_OAI21X1_111 gnd vdd FILL
XDFFPOSX1_585 BUFX2_616/A CLKBUF1_23/Y OAI21X1_765/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_772 gnd vdd FILL
XDFFPOSX1_596 BUFX2_628/A CLKBUF1_100/Y OAI21X1_799/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_122 gnd vdd FILL
XNAND2X1_600 INVX1_203/Y AND2X2_26/Y gnd NOR2X1_193/B vdd NAND2X1
XFILL_1_OAI21X1_144 gnd vdd FILL
XNAND2X1_611 MUX2X1_2/S NOR3X1_16/C gnd NAND2X1_611/Y vdd NAND2X1
XFILL_1_DFFPOSX1_783 gnd vdd FILL
XFILL_1_DFFPOSX1_794 gnd vdd FILL
XFILL_1_OAI21X1_166 gnd vdd FILL
XNAND2X1_633 NAND2X1_633/A XNOR2X1_98/A gnd NAND2X1_633/Y vdd NAND2X1
XINVX1_23 NOR3X1_4/B gnd INVX1_23/Y vdd INVX1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XNAND2X1_622 INVX1_214/Y NOR3X1_18/Y gnd INVX1_215/A vdd NAND2X1
XNAND2X1_644 NAND2X1_644/A INVX1_226/A gnd NAND2X1_644/Y vdd NAND2X1
XFILL_2_OAI21X1_348 gnd vdd FILL
XFILL_1_OAI21X1_155 gnd vdd FILL
XNAND2X1_655 BUFX2_676/A OAI21X1_7/A gnd NAND2X1_655/Y vdd NAND2X1
XFILL_1_OAI21X1_177 gnd vdd FILL
XNAND2X1_666 BUFX2_657/A BUFX4_312/Y gnd NAND2X1_666/Y vdd NAND2X1
XNAND2X1_677 BUFX2_669/A OAI21X1_1/A gnd NAND2X1_677/Y vdd NAND2X1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XFILL_1_OAI21X1_199 gnd vdd FILL
XINVX1_67 INVX1_67/A gnd INVX1_67/Y vdd INVX1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XFILL_1_OAI21X1_188 gnd vdd FILL
XFILL_2_OAI21X1_359 gnd vdd FILL
XNAND2X1_688 BUFX2_709/A BUFX4_217/Y gnd NAND2X1_688/Y vdd NAND2X1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XNAND2X1_699 BUFX2_690/A BUFX4_220/Y gnd NAND2X1_699/Y vdd NAND2X1
XINVX1_78 bundle_i[62] gnd INVX1_78/Y vdd INVX1
XINVX1_89 bundle_i[51] gnd INVX1_89/Y vdd INVX1
XDFFPOSX1_8 BUFX2_707/A CLKBUF1_87/Y DFFPOSX1_8/D gnd vdd DFFPOSX1
XFILL_1_NAND2X1_150 gnd vdd FILL
XFILL_0_DFFPOSX1_340 gnd vdd FILL
XFILL_1_NAND2X1_172 gnd vdd FILL
XFILL_0_DFFPOSX1_351 gnd vdd FILL
XFILL_1_NAND2X1_194 gnd vdd FILL
XFILL_0_DFFPOSX1_384 gnd vdd FILL
XFILL_0_DFFPOSX1_373 gnd vdd FILL
XFILL_0_DFFPOSX1_362 gnd vdd FILL
XFILL_26_13_1 gnd vdd FILL
XFILL_0_DFFPOSX1_395 gnd vdd FILL
XFILL_3_DFFPOSX1_822 gnd vdd FILL
XFILL_3_DFFPOSX1_811 gnd vdd FILL
XFILL_3_DFFPOSX1_800 gnd vdd FILL
XFILL_3_DFFPOSX1_855 gnd vdd FILL
XFILL_3_DFFPOSX1_833 gnd vdd FILL
XFILL_3_DFFPOSX1_866 gnd vdd FILL
XFILL_3_DFFPOSX1_844 gnd vdd FILL
XFILL_3_DFFPOSX1_888 gnd vdd FILL
XFILL_3_DFFPOSX1_877 gnd vdd FILL
XFILL_3_DFFPOSX1_899 gnd vdd FILL
XFILL_2_DFFPOSX1_412 gnd vdd FILL
XBUFX2_521 BUFX2_521/A gnd majID3_o[63] vdd BUFX2
XFILL_2_DFFPOSX1_423 gnd vdd FILL
XFILL_2_DFFPOSX1_401 gnd vdd FILL
XBUFX2_510 BUFX2_510/A gnd majID2_o[6] vdd BUFX2
XFILL_4_DFFPOSX1_30 gnd vdd FILL
XFILL_2_DFFPOSX1_456 gnd vdd FILL
XBUFX2_532 BUFX2_532/A gnd majID3_o[44] vdd BUFX2
XFILL_2_DFFPOSX1_445 gnd vdd FILL
XBUFX2_543 BUFX2_543/A gnd majID3_o[34] vdd BUFX2
XFILL_1_14_1 gnd vdd FILL
XFILL_2_DFFPOSX1_434 gnd vdd FILL
XBUFX2_554 INVX1_29/A gnd majID3_o[24] vdd BUFX2
XFILL_4_DFFPOSX1_41 gnd vdd FILL
XBUFX2_576 BUFX2_576/A gnd majID3_o[4] vdd BUFX2
XFILL_2_DFFPOSX1_478 gnd vdd FILL
XFILL_4_DFFPOSX1_52 gnd vdd FILL
XFILL_4_DFFPOSX1_63 gnd vdd FILL
XBUFX2_565 BUFX2_565/A gnd majID3_o[14] vdd BUFX2
XFILL_2_DFFPOSX1_489 gnd vdd FILL
XBUFX2_587 BUFX2_587/A gnd majID4_o[53] vdd BUFX2
XFILL_2_DFFPOSX1_467 gnd vdd FILL
XFILL_4_DFFPOSX1_74 gnd vdd FILL
XFILL_4_DFFPOSX1_85 gnd vdd FILL
XFILL_4_DFFPOSX1_96 gnd vdd FILL
XBUFX2_598 BUFX2_598/A gnd majID4_o[43] vdd BUFX2
XFILL_31_6_0 gnd vdd FILL
XFILL_5_DFFPOSX1_938 gnd vdd FILL
XFILL_5_DFFPOSX1_905 gnd vdd FILL
XFILL_5_DFFPOSX1_916 gnd vdd FILL
XFILL_5_DFFPOSX1_927 gnd vdd FILL
XFILL_5_DFFPOSX1_949 gnd vdd FILL
XFILL_0_BUFX2_250 gnd vdd FILL
XFILL_0_BUFX2_283 gnd vdd FILL
XFILL_0_AND2X2_7 gnd vdd FILL
XFILL_0_BUFX2_272 gnd vdd FILL
XFILL_0_BUFX2_261 gnd vdd FILL
XFILL_0_BUFX2_294 gnd vdd FILL
XFILL_4_DFFPOSX1_528 gnd vdd FILL
XFILL_4_DFFPOSX1_506 gnd vdd FILL
XFILL_4_DFFPOSX1_517 gnd vdd FILL
XFILL_4_DFFPOSX1_539 gnd vdd FILL
XFILL_6_13_1 gnd vdd FILL
XFILL_1_BUFX2_1019 gnd vdd FILL
XFILL_2_DFFPOSX1_990 gnd vdd FILL
XFILL_22_6_0 gnd vdd FILL
XFILL_1_BUFX2_418 gnd vdd FILL
XFILL_1_BUFX2_429 gnd vdd FILL
XFILL_0_NAND3X1_2 gnd vdd FILL
XOAI21X1_413 NOR2X1_6/B INVX4_3/Y INVX2_15/Y gnd OAI21X1_414/C vdd OAI21X1
XOAI21X1_402 INVX2_40/Y INVX2_11/Y INVX2_12/Y gnd OAI21X1_403/C vdd OAI21X1
XFILL_3_DFFPOSX1_118 gnd vdd FILL
XFILL_3_DFFPOSX1_107 gnd vdd FILL
XOAI21X1_457 XNOR2X1_18/Y BUFX4_213/Y OAI21X1_457/C gnd OAI21X1_457/Y vdd OAI21X1
XOAI21X1_446 NOR2X1_21/Y AOI21X1_2/Y BUFX4_245/Y gnd OAI21X1_447/C vdd OAI21X1
XOAI21X1_424 INVX1_10/Y OAI21X1_424/B OAI21X1_424/C gnd OAI21X1_424/Y vdd OAI21X1
XOAI21X1_435 INVX1_11/Y bundleStartMajId_i[39] BUFX4_245/Y gnd OAI21X1_436/A vdd OAI21X1
XOAI21X1_479 NOR2X1_47/Y bundleStartMajId_i[11] BUFX4_240/Y gnd OAI21X1_480/B vdd
+ OAI21X1
XFILL_3_DFFPOSX1_129 gnd vdd FILL
XOAI21X1_468 AND2X2_9/Y bundleStartMajId_i[17] BUFX4_244/Y gnd OAI21X1_469/A vdd OAI21X1
XFILL_3_XNOR2X1_92 gnd vdd FILL
XDFFPOSX1_382 BUFX2_412/A CLKBUF1_50/Y OAI21X1_354/Y gnd vdd DFFPOSX1
XDFFPOSX1_360 BUFX2_427/A CLKBUF1_41/Y OAI21X1_332/Y gnd vdd DFFPOSX1
XDFFPOSX1_371 BUFX2_400/A CLKBUF1_13/Y OAI21X1_343/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_591 gnd vdd FILL
XFILL_2_OAI21X1_123 gnd vdd FILL
XFILL_1_DFFPOSX1_580 gnd vdd FILL
XDFFPOSX1_393 BUFX2_424/A CLKBUF1_24/Y OAI21X1_365/Y gnd vdd DFFPOSX1
XNAND2X1_430 BUFX2_22/A BUFX4_311/Y gnd NAND2X1_430/Y vdd NAND2X1
XNAND2X1_463 BUFX2_59/A BUFX4_357/Y gnd NAND2X1_463/Y vdd NAND2X1
XNAND2X1_441 BUFX2_34/A BUFX4_350/Y gnd NAND2X1_441/Y vdd NAND2X1
XNAND2X1_452 BUFX2_47/A BUFX4_364/Y gnd NAND2X1_452/Y vdd NAND2X1
XNAND2X1_474 bundleAddress_i[58] bundleAddress_i[57] gnd NOR2X1_124/B vdd NAND2X1
XNAND2X1_485 BUFX2_68/A BUFX4_231/Y gnd NAND2X1_485/Y vdd NAND2X1
XNAND2X1_496 BUFX2_72/A OAI21X1_8/B gnd NAND2X1_496/Y vdd NAND2X1
XFILL_5_7_0 gnd vdd FILL
XFILL_0_INVX1_206 gnd vdd FILL
XFILL_0_INVX1_217 gnd vdd FILL
XFILL_13_6_0 gnd vdd FILL
XFILL_0_DFFPOSX1_181 gnd vdd FILL
XFILL_0_DFFPOSX1_170 gnd vdd FILL
XFILL_0_DFFPOSX1_192 gnd vdd FILL
XFILL_0_OAI21X1_38 gnd vdd FILL
XFILL_0_OAI21X1_27 gnd vdd FILL
XFILL_1_BUFX2_952 gnd vdd FILL
XFILL_0_OAI21X1_16 gnd vdd FILL
XFILL_1_BUFX2_941 gnd vdd FILL
XFILL_1_BUFX2_996 gnd vdd FILL
XFILL_1_BUFX2_985 gnd vdd FILL
XFILL_3_DFFPOSX1_630 gnd vdd FILL
XFILL_0_OAI21X1_49 gnd vdd FILL
XFILL_3_DFFPOSX1_641 gnd vdd FILL
XOAI21X1_1709 BUFX4_173/Y INVX2_116/Y OAI21X1_1709/C gnd DFFPOSX1_67/D vdd OAI21X1
XOAI21X1_991 BUFX4_296/Y INVX1_150/Y OAI21X1_991/C gnd OAI21X1_991/Y vdd OAI21X1
XOAI21X1_980 BUFX4_140/Y BUFX4_39/Y BUFX2_383/A gnd OAI21X1_981/C vdd OAI21X1
XFILL_3_DFFPOSX1_652 gnd vdd FILL
XFILL_3_DFFPOSX1_663 gnd vdd FILL
XFILL_3_DFFPOSX1_674 gnd vdd FILL
XFILL_0_OAI21X1_709 gnd vdd FILL
XFILL_3_DFFPOSX1_696 gnd vdd FILL
XFILL_3_DFFPOSX1_685 gnd vdd FILL
XFILL_17_18_1 gnd vdd FILL
XFILL_2_DFFPOSX1_220 gnd vdd FILL
XFILL_0_NAND2X1_726 gnd vdd FILL
XFILL_0_NAND2X1_704 gnd vdd FILL
XFILL_0_NAND2X1_715 gnd vdd FILL
XFILL_2_DFFPOSX1_231 gnd vdd FILL
XFILL_11_14_0 gnd vdd FILL
XFILL_2_DFFPOSX1_242 gnd vdd FILL
XBUFX2_362 BUFX2_362/A gnd instr4_o[18] vdd BUFX2
XFILL_0_NAND2X1_748 gnd vdd FILL
XFILL_5_DFFPOSX1_20 gnd vdd FILL
XFILL_0_NAND2X1_759 gnd vdd FILL
XFILL_0_NAND2X1_737 gnd vdd FILL
XFILL_0_OAI21X1_1519 gnd vdd FILL
XFILL_2_DFFPOSX1_253 gnd vdd FILL
XFILL_2_DFFPOSX1_264 gnd vdd FILL
XBUFX2_340 BUFX2_340/A gnd instr3_o[9] vdd BUFX2
XFILL_0_OAI21X1_1508 gnd vdd FILL
XBUFX2_351 BUFX2_351/A gnd instr3_o[27] vdd BUFX2
XFILL_2_DFFPOSX1_275 gnd vdd FILL
XFILL_5_DFFPOSX1_53 gnd vdd FILL
XFILL_5_DFFPOSX1_64 gnd vdd FILL
XBUFX2_373 BUFX2_373/A gnd instr4_o[8] vdd BUFX2
XBUFX2_384 BUFX2_384/A gnd instr4_o[26] vdd BUFX2
XBUFX2_395 BUFX2_395/A gnd majID1_o[53] vdd BUFX2
XFILL_5_DFFPOSX1_31 gnd vdd FILL
XFILL_2_DFFPOSX1_297 gnd vdd FILL
XFILL_2_DFFPOSX1_286 gnd vdd FILL
XFILL_5_DFFPOSX1_42 gnd vdd FILL
XFILL_5_DFFPOSX1_75 gnd vdd FILL
XFILL_5_DFFPOSX1_86 gnd vdd FILL
XFILL_5_DFFPOSX1_97 gnd vdd FILL
XFILL_5_DFFPOSX1_702 gnd vdd FILL
XFILL_1_NOR3X1_12 gnd vdd FILL
XFILL_5_DFFPOSX1_713 gnd vdd FILL
XFILL_5_DFFPOSX1_746 gnd vdd FILL
XOAI21X1_62 INVX2_200/Y BUFX4_208/Y OAI21X1_62/C gnd OAI21X1_62/Y vdd OAI21X1
XOAI21X1_51 INVX2_189/Y BUFX4_193/Y OAI21X1_51/C gnd OAI21X1_51/Y vdd OAI21X1
XFILL_5_DFFPOSX1_735 gnd vdd FILL
XOAI21X1_40 INVX2_178/Y BUFX4_215/Y OAI21X1_40/C gnd OAI21X1_40/Y vdd OAI21X1
XFILL_5_DFFPOSX1_724 gnd vdd FILL
XOAI21X1_84 BUFX4_5/Y BUFX4_341/Y BUFX2_961/A gnd OAI21X1_85/C vdd OAI21X1
XOAI21X1_95 BUFX4_178/Y INVX2_157/Y OAI21X1_95/C gnd OAI21X1_95/Y vdd OAI21X1
XOAI21X1_73 BUFX4_149/Y OAI21X1_8/A OAI21X1_73/C gnd OAI21X1_73/Y vdd OAI21X1
XFILL_5_DFFPOSX1_757 gnd vdd FILL
XFILL_5_DFFPOSX1_779 gnd vdd FILL
XFILL_5_DFFPOSX1_768 gnd vdd FILL
XFILL_4_DFFPOSX1_303 gnd vdd FILL
XFILL_4_DFFPOSX1_336 gnd vdd FILL
XFILL_4_DFFPOSX1_325 gnd vdd FILL
XFILL_0_DFFPOSX1_60 gnd vdd FILL
XFILL_4_DFFPOSX1_314 gnd vdd FILL
XFILL_0_DFFPOSX1_71 gnd vdd FILL
XFILL_16_13_0 gnd vdd FILL
XFILL_0_DFFPOSX1_82 gnd vdd FILL
XFILL_0_DFFPOSX1_93 gnd vdd FILL
XFILL_4_DFFPOSX1_358 gnd vdd FILL
XFILL_4_DFFPOSX1_347 gnd vdd FILL
XFILL_4_DFFPOSX1_369 gnd vdd FILL
XFILL_2_DFFPOSX1_1017 gnd vdd FILL
XFILL_2_DFFPOSX1_1006 gnd vdd FILL
XFILL_2_DFFPOSX1_1028 gnd vdd FILL
XFILL_1_BUFX2_226 gnd vdd FILL
XFILL_1_BUFX2_237 gnd vdd FILL
XOAI21X1_221 INVX2_156/Y INVX8_2/A OAI21X1_221/C gnd OAI21X1_221/Y vdd OAI21X1
XOAI21X1_210 BUFX4_158/Y BUFX4_59/Y BUFX2_1014/A gnd OAI21X1_211/C vdd OAI21X1
XOAI21X1_254 BUFX4_165/Y BUFX4_34/Y BUFX2_989/A gnd OAI21X1_255/C vdd OAI21X1
XOAI21X1_232 BUFX4_147/Y BUFX4_77/Y BUFX2_977/A gnd OAI21X1_233/C vdd OAI21X1
XOAI21X1_243 INVX2_167/Y BUFX4_296/Y OAI21X1_243/C gnd OAI21X1_243/Y vdd OAI21X1
XOAI21X1_265 INVX2_178/Y BUFX4_302/Y OAI21X1_265/C gnd OAI21X1_265/Y vdd OAI21X1
XOAI21X1_276 BUFX4_137/Y BUFX4_47/Y BUFX2_1001/A gnd OAI21X1_277/C vdd OAI21X1
XOAI21X1_298 BUFX4_137/Y BUFX4_66/Y BUFX2_1013/A gnd OAI21X1_299/C vdd OAI21X1
XOAI21X1_287 INVX2_189/Y BUFX4_301/Y OAI21X1_287/C gnd OAI21X1_287/Y vdd OAI21X1
XAND2X2_32 INVX1_211/A AND2X2_32/B gnd AND2X2_33/B vdd AND2X2
XAND2X2_21 AND2X2_21/A NOR3X1_6/A gnd AND2X2_21/Y vdd AND2X2
XAND2X2_10 NOR2X1_47/Y NOR2X1_50/Y gnd AND2X2_10/Y vdd AND2X2
XFILL_6_DFFPOSX1_408 gnd vdd FILL
XDFFPOSX1_190 BUFX2_860/A CLKBUF1_3/Y OAI21X1_34/Y gnd vdd DFFPOSX1
XFILL_6_DFFPOSX1_419 gnd vdd FILL
XFILL_34_14_0 gnd vdd FILL
XNAND2X1_260 bundleStartMajId_i[3] INVX1_44/A gnd NOR3X1_4/B vdd NAND2X1
XNAND2X1_271 INVX4_30/Y OAI21X1_522/Y gnd OAI21X1_524/A vdd NAND2X1
XNAND2X1_282 NOR2X1_69/Y INVX1_27/Y gnd NOR2X1_70/B vdd NAND2X1
XNAND2X1_293 bundleStartMajId_i[24] bundleStartMajId_i[23] gnd NOR2X1_83/B vdd NAND2X1
XFILL_4_DFFPOSX1_881 gnd vdd FILL
XFILL_4_DFFPOSX1_870 gnd vdd FILL
XFILL_4_DFFPOSX1_892 gnd vdd FILL
XFILL_0_INVX8_6 gnd vdd FILL
XFILL_0_BUFX4_312 gnd vdd FILL
XFILL_1_BUFX2_760 gnd vdd FILL
XFILL_0_BUFX4_301 gnd vdd FILL
XFILL_0_BUFX4_323 gnd vdd FILL
XFILL_0_BUFX4_334 gnd vdd FILL
XFILL_1_BUFX2_782 gnd vdd FILL
XFILL_1_OAI21X1_1715 gnd vdd FILL
XFILL_1_BUFX2_793 gnd vdd FILL
XFILL_0_BUFX4_356 gnd vdd FILL
XOAI21X1_1528 BUFX4_121/Y BUFX4_38/Y BUFX2_236/A gnd OAI21X1_1530/C vdd OAI21X1
XOAI21X1_1517 OAI21X1_1517/A AOI21X1_61/Y OAI21X1_1517/C gnd OAI21X1_1517/Y vdd OAI21X1
XFILL_0_BUFX4_367 gnd vdd FILL
XOAI21X1_1506 NAND3X1_65/Y NOR3X1_16/B INVX4_42/Y gnd OAI21X1_1507/C vdd OAI21X1
XFILL_1_OAI21X1_1704 gnd vdd FILL
XOAI21X1_1539 OAI21X1_1539/A BUFX4_294/Y OAI21X1_1539/C gnd OAI21X1_1539/Y vdd OAI21X1
XFILL_0_BUFX4_345 gnd vdd FILL
XFILL_1_OAI21X1_1726 gnd vdd FILL
XFILL_1_OAI21X1_1737 gnd vdd FILL
XFILL_3_DFFPOSX1_471 gnd vdd FILL
XFILL_3_DFFPOSX1_482 gnd vdd FILL
XFILL_1_OAI21X1_1748 gnd vdd FILL
XFILL_0_BUFX4_378 gnd vdd FILL
XFILL_3_DFFPOSX1_460 gnd vdd FILL
XFILL_0_BUFX2_1005 gnd vdd FILL
XFILL_1_OAI21X1_1759 gnd vdd FILL
XFILL_3_DFFPOSX1_493 gnd vdd FILL
XFILL_0_BUFX2_1016 gnd vdd FILL
XFILL_0_OAI21X1_506 gnd vdd FILL
XFILL_0_OAI21X1_528 gnd vdd FILL
XFILL_0_OAI21X1_517 gnd vdd FILL
XFILL_0_BUFX2_1027 gnd vdd FILL
XFILL_0_OAI21X1_539 gnd vdd FILL
XFILL_6_DFFPOSX1_997 gnd vdd FILL
XFILL_6_DFFPOSX1_986 gnd vdd FILL
XFILL_6_DFFPOSX1_975 gnd vdd FILL
XFILL_0_CLKBUF1_17 gnd vdd FILL
XFILL_0_CLKBUF1_39 gnd vdd FILL
XFILL_0_NAND2X1_501 gnd vdd FILL
XFILL_0_CLKBUF1_28 gnd vdd FILL
XFILL_1_NAND2X1_705 gnd vdd FILL
XFILL_36_5_0 gnd vdd FILL
XFILL_0_NAND2X1_523 gnd vdd FILL
XFILL_0_NAND2X1_534 gnd vdd FILL
XFILL_0_NAND2X1_512 gnd vdd FILL
XFILL_1_NAND2X1_716 gnd vdd FILL
XFILL_0_OAI21X1_1305 gnd vdd FILL
XFILL_1_NAND2X1_749 gnd vdd FILL
XFILL_0_OAI21X1_1338 gnd vdd FILL
XFILL_0_DFFPOSX1_906 gnd vdd FILL
XBUFX2_170 BUFX2_170/A gnd addr3_o[17] vdd BUFX2
XFILL_0_NAND2X1_556 gnd vdd FILL
XFILL_0_OAI21X1_1327 gnd vdd FILL
XFILL_0_NAND2X1_567 gnd vdd FILL
XFILL_0_OAI21X1_1349 gnd vdd FILL
XFILL_0_NAND2X1_578 gnd vdd FILL
XFILL_0_NAND2X1_545 gnd vdd FILL
XFILL_0_OAI21X1_1316 gnd vdd FILL
XBUFX2_192 BUFX2_192/A gnd addr3_o[54] vdd BUFX2
XFILL_0_DFFPOSX1_939 gnd vdd FILL
XFILL_0_NAND2X1_589 gnd vdd FILL
XFILL_0_DFFPOSX1_917 gnd vdd FILL
XBUFX2_181 BUFX2_181/A gnd addr3_o[7] vdd BUFX2
XFILL_0_DFFPOSX1_928 gnd vdd FILL
XFILL_6_DFFPOSX1_76 gnd vdd FILL
XFILL_5_DFFPOSX1_510 gnd vdd FILL
XFILL_6_DFFPOSX1_87 gnd vdd FILL
XFILL_6_DFFPOSX1_65 gnd vdd FILL
XFILL_5_DFFPOSX1_521 gnd vdd FILL
XFILL_5_DFFPOSX1_543 gnd vdd FILL
XFILL_20_9_1 gnd vdd FILL
XFILL_5_DFFPOSX1_532 gnd vdd FILL
XFILL_6_DFFPOSX1_98 gnd vdd FILL
XFILL_5_DFFPOSX1_554 gnd vdd FILL
XFILL_5_DFFPOSX1_587 gnd vdd FILL
XFILL_5_DFFPOSX1_576 gnd vdd FILL
XFILL_5_DFFPOSX1_565 gnd vdd FILL
XFILL_5_DFFPOSX1_598 gnd vdd FILL
XFILL_1_AOI21X1_5 gnd vdd FILL
XFILL_1_BUFX4_9 gnd vdd FILL
XFILL_4_DFFPOSX1_111 gnd vdd FILL
XFILL_4_DFFPOSX1_100 gnd vdd FILL
XCLKBUF1_30 BUFX4_87/Y gnd CLKBUF1_30/Y vdd CLKBUF1
XCLKBUF1_41 BUFX4_90/Y gnd CLKBUF1_41/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_133 gnd vdd FILL
XFILL_1_DFFPOSX1_50 gnd vdd FILL
XFILL_4_DFFPOSX1_144 gnd vdd FILL
XCLKBUF1_74 BUFX4_85/Y gnd CLKBUF1_74/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_122 gnd vdd FILL
XCLKBUF1_63 BUFX4_91/Y gnd CLKBUF1_63/Y vdd CLKBUF1
XCLKBUF1_52 BUFX4_88/Y gnd CLKBUF1_52/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_83 gnd vdd FILL
XCLKBUF1_96 BUFX4_85/Y gnd CLKBUF1_96/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_61 gnd vdd FILL
XFILL_4_DFFPOSX1_155 gnd vdd FILL
XFILL_1_DFFPOSX1_72 gnd vdd FILL
XCLKBUF1_85 BUFX4_88/Y gnd CLKBUF1_85/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_166 gnd vdd FILL
XFILL_4_DFFPOSX1_177 gnd vdd FILL
XFILL_4_DFFPOSX1_188 gnd vdd FILL
XFILL_1_DFFPOSX1_94 gnd vdd FILL
XFILL_27_5_0 gnd vdd FILL
XFILL_4_DFFPOSX1_199 gnd vdd FILL
XFILL_2_5_0 gnd vdd FILL
XFILL_2_BUFX4_254 gnd vdd FILL
XFILL_2_BUFX4_298 gnd vdd FILL
XFILL_11_9_1 gnd vdd FILL
XFILL_10_4_0 gnd vdd FILL
XFILL_0_BUFX2_805 gnd vdd FILL
XFILL_0_BUFX2_816 gnd vdd FILL
XFILL_23_11_1 gnd vdd FILL
XFILL_0_BUFX2_849 gnd vdd FILL
XFILL_0_BUFX2_827 gnd vdd FILL
XFILL_0_BUFX2_838 gnd vdd FILL
XINVX1_115 bundle_i[89] gnd INVX1_115/Y vdd INVX1
XINVX1_104 bundle_i[36] gnd INVX1_104/Y vdd INVX1
XINVX1_148 bundle_i[120] gnd INVX1_148/Y vdd INVX1
XINVX1_126 bundle_i[78] gnd INVX1_126/Y vdd INVX1
XINVX1_137 bundle_i[67] gnd INVX1_137/Y vdd INVX1
XFILL_3_XNOR2X1_3 gnd vdd FILL
XINVX1_159 bundle_i[109] gnd INVX1_159/Y vdd INVX1
XFILL_0_INVX2_25 gnd vdd FILL
XFILL_0_INVX2_36 gnd vdd FILL
XFILL_0_INVX2_14 gnd vdd FILL
XFILL_0_INVX2_58 gnd vdd FILL
XFILL_0_INVX2_47 gnd vdd FILL
XFILL_0_INVX2_69 gnd vdd FILL
XFILL_18_5_0 gnd vdd FILL
XFILL_0_CLKBUF1_4 gnd vdd FILL
XFILL_28_10_1 gnd vdd FILL
XFILL_4_CLKBUF1_3 gnd vdd FILL
XFILL_3_XNOR2X1_100 gnd vdd FILL
XOAI21X1_1303 OAI21X1_1303/A BUFX4_170/Y OAI21X1_1303/C gnd OAI21X1_1303/Y vdd OAI21X1
XFILL_0_BUFX4_142 gnd vdd FILL
XFILL_0_BUFX4_120 gnd vdd FILL
XFILL_1_BUFX2_590 gnd vdd FILL
XFILL_0_BUFX4_131 gnd vdd FILL
XOAI21X1_1314 BUFX4_6/A BUFX4_370/Y BUFX2_162/A gnd OAI21X1_1315/C vdd OAI21X1
XFILL_0_BUFX4_164 gnd vdd FILL
XOAI21X1_1336 BUFX4_103/Y BUFX4_339/Y BUFX2_171/A gnd OAI21X1_1338/C vdd OAI21X1
XDFFPOSX1_904 BUFX2_155/A CLKBUF1_68/Y OAI21X1_1296/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1523 gnd vdd FILL
XDFFPOSX1_915 BUFX2_167/A CLKBUF1_49/Y OAI21X1_1327/Y gnd vdd DFFPOSX1
XFILL_0_BUFX4_175 gnd vdd FILL
XFILL_1_OAI21X1_1512 gnd vdd FILL
XOAI21X1_1325 INVX2_106/Y NOR3X1_17/B INVX4_43/Y gnd NAND2X1_616/B vdd OAI21X1
XOAI21X1_1347 AOI21X1_54/Y OAI21X1_1347/B OAI21X1_1347/C gnd OAI21X1_1347/Y vdd OAI21X1
XFILL_0_BUFX4_153 gnd vdd FILL
XFILL_1_OAI21X1_1501 gnd vdd FILL
XFILL_0_BUFX4_197 gnd vdd FILL
XDFFPOSX1_948 BUFX2_197/A CLKBUF1_29/Y OAI21X1_1420/Y gnd vdd DFFPOSX1
XFILL_1_BUFX2_42 gnd vdd FILL
XDFFPOSX1_937 BUFX2_194/A CLKBUF1_73/Y OAI21X1_1387/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1567 gnd vdd FILL
XOAI21X1_1369 NOR2X1_211/B INVX1_216/Y OAI21X1_1369/C gnd OAI21X1_1371/A vdd OAI21X1
XFILL_3_DFFPOSX1_290 gnd vdd FILL
XFILL_0_OAI21X1_303 gnd vdd FILL
XOAI21X1_1358 BUFX4_1/A BUFX4_357/Y BUFX2_180/A gnd OAI21X1_1360/C vdd OAI21X1
XFILL_1_OAI21X1_1556 gnd vdd FILL
XFILL_1_OAI21X1_1534 gnd vdd FILL
XFILL_0_BUFX4_186 gnd vdd FILL
XFILL_1_BUFX2_31 gnd vdd FILL
XDFFPOSX1_926 BUFX2_179/A CLKBUF1_76/Y OAI21X1_1357/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1545 gnd vdd FILL
XFILL_1_OAI21X1_1589 gnd vdd FILL
XFILL_0_OAI21X1_314 gnd vdd FILL
XFILL_1_OAI21X1_1578 gnd vdd FILL
XFILL_0_OAI21X1_325 gnd vdd FILL
XDFFPOSX1_959 BUFX2_209/A CLKBUF1_34/Y OAI21X1_1453/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_507 gnd vdd FILL
XFILL_1_BUFX2_97 gnd vdd FILL
XFILL_0_OAI21X1_336 gnd vdd FILL
XFILL_1_BUFX2_86 gnd vdd FILL
XFILL_1_BUFX2_75 gnd vdd FILL
XFILL_1_OAI21X1_518 gnd vdd FILL
XFILL_0_OAI21X1_347 gnd vdd FILL
XFILL_0_OAI21X1_369 gnd vdd FILL
XFILL_0_OAI21X1_358 gnd vdd FILL
XFILL_1_OAI21X1_529 gnd vdd FILL
XFILL_6_DFFPOSX1_761 gnd vdd FILL
XFILL_6_DFFPOSX1_750 gnd vdd FILL
XFILL_6_DFFPOSX1_772 gnd vdd FILL
XFILL_6_DFFPOSX1_783 gnd vdd FILL
XFILL_1_OAI21X1_8 gnd vdd FILL
XFILL_3_11_1 gnd vdd FILL
XFILL_0_OAI21X1_1102 gnd vdd FILL
XFILL_0_OAI21X1_1124 gnd vdd FILL
XFILL_0_OAI21X1_1113 gnd vdd FILL
XFILL_1_NAND2X1_524 gnd vdd FILL
XFILL_0_NAND2X1_331 gnd vdd FILL
XFILL_0_NAND2X1_320 gnd vdd FILL
XFILL_0_NAND2X1_342 gnd vdd FILL
XFILL_0_NAND2X1_353 gnd vdd FILL
XFILL_0_NAND2X1_386 gnd vdd FILL
XFILL_0_NAND2X1_375 gnd vdd FILL
XFILL_0_DFFPOSX1_725 gnd vdd FILL
XFILL_0_OAI21X1_1146 gnd vdd FILL
XFILL_0_NAND2X1_364 gnd vdd FILL
XFILL_1_NAND2X1_557 gnd vdd FILL
XFILL_0_DFFPOSX1_714 gnd vdd FILL
XFILL_0_OAI21X1_1157 gnd vdd FILL
XFILL_0_DFFPOSX1_703 gnd vdd FILL
XFILL_0_OAI21X1_1135 gnd vdd FILL
XFILL_0_DFFPOSX1_747 gnd vdd FILL
XFILL_0_DFFPOSX1_758 gnd vdd FILL
XFILL_0_DFFPOSX1_736 gnd vdd FILL
XFILL_0_OAI21X1_1168 gnd vdd FILL
XFILL_0_OAI21X1_1179 gnd vdd FILL
XFILL_0_NAND2X1_397 gnd vdd FILL
XFILL_0_DFFPOSX1_769 gnd vdd FILL
XFILL_5_DFFPOSX1_340 gnd vdd FILL
XFILL_5_DFFPOSX1_362 gnd vdd FILL
XFILL_5_DFFPOSX1_351 gnd vdd FILL
XFILL_5_DFFPOSX1_395 gnd vdd FILL
XFILL_5_DFFPOSX1_384 gnd vdd FILL
XFILL_5_DFFPOSX1_373 gnd vdd FILL
XFILL_1_NAND2X1_22 gnd vdd FILL
XFILL_1_NAND2X1_44 gnd vdd FILL
XINVX4_34 bundleAddress_i[47] gnd INVX4_34/Y vdd INVX4
XINVX4_23 bundleStartMajId_i[14] gnd INVX4_23/Y vdd INVX4
XINVX4_12 bundleStartMajId_i[36] gnd INVX4_12/Y vdd INVX4
XINVX4_45 bundleAddress_i[8] gnd INVX4_45/Y vdd INVX4
XFILL_1_NAND2X1_66 gnd vdd FILL
XFILL_1_NAND2X1_99 gnd vdd FILL
XFILL_0_OAI21X1_892 gnd vdd FILL
XFILL_1_BUFX2_6 gnd vdd FILL
XFILL_0_OAI21X1_881 gnd vdd FILL
XFILL_0_OAI21X1_870 gnd vdd FILL
XFILL_8_10_1 gnd vdd FILL
XFILL_2_OAI21X1_1218 gnd vdd FILL
XFILL_2_DFFPOSX1_808 gnd vdd FILL
XBUFX2_906 BUFX2_906/A gnd tid3_o[62] vdd BUFX2
XFILL_2_DFFPOSX1_51 gnd vdd FILL
XFILL_2_DFFPOSX1_819 gnd vdd FILL
XFILL_2_DFFPOSX1_62 gnd vdd FILL
XFILL_2_DFFPOSX1_40 gnd vdd FILL
XBUFX2_928 BUFX2_928/A gnd tid3_o[60] vdd BUFX2
XBUFX2_917 BUFX2_917/A gnd tid3_o[61] vdd BUFX2
XFILL_2_DFFPOSX1_73 gnd vdd FILL
XBUFX2_939 BUFX2_939/A gnd tid3_o[59] vdd BUFX2
XFILL_2_DFFPOSX1_84 gnd vdd FILL
XFILL_2_DFFPOSX1_95 gnd vdd FILL
XFILL_0_OAI21X1_1691 gnd vdd FILL
XFILL_0_OAI21X1_1680 gnd vdd FILL
XFILL_0_BUFX2_613 gnd vdd FILL
XFILL_0_BUFX2_624 gnd vdd FILL
XFILL_0_BUFX2_602 gnd vdd FILL
XFILL_0_BUFX2_657 gnd vdd FILL
XFILL_0_BUFX2_646 gnd vdd FILL
XFILL_1_DFFPOSX1_409 gnd vdd FILL
XFILL_0_BUFX2_635 gnd vdd FILL
XFILL_4_DFFPOSX1_1030 gnd vdd FILL
XFILL_0_BUFX2_679 gnd vdd FILL
XFILL_0_BUFX2_668 gnd vdd FILL
XBUFX4_210 BUFX4_25/Y gnd OAI21X1_8/B vdd BUFX4
XBUFX4_221 BUFX4_25/Y gnd BUFX4_221/Y vdd BUFX4
XFILL_14_16_1 gnd vdd FILL
XBUFX4_243 INVX8_1/Y gnd BUFX4_243/Y vdd BUFX4
XBUFX4_254 INVX8_5/Y gnd BUFX4_7/A vdd BUFX4
XBUFX4_232 BUFX4_20/Y gnd BUFX4_232/Y vdd BUFX4
XFILL_0_INVX2_131 gnd vdd FILL
XFILL_0_INVX2_153 gnd vdd FILL
XBUFX4_265 enable_i gnd BUFX4_265/Y vdd BUFX4
XBUFX4_298 BUFX4_303/A gnd INVX8_2/A vdd BUFX4
XBUFX4_287 INVX8_2/Y gnd BUFX4_287/Y vdd BUFX4
XBUFX4_276 INVX8_7/Y gnd BUFX4_66/A vdd BUFX4
XFILL_0_INVX2_120 gnd vdd FILL
XFILL_0_INVX2_142 gnd vdd FILL
XFILL_34_8_1 gnd vdd FILL
XFILL_0_INVX2_164 gnd vdd FILL
XFILL_0_INVX2_175 gnd vdd FILL
XFILL_0_INVX2_186 gnd vdd FILL
XFILL_33_3_0 gnd vdd FILL
XFILL_25_2 gnd vdd FILL
XFILL_0_INVX2_197 gnd vdd FILL
XFILL_18_1 gnd vdd FILL
XOAI21X1_809 OAI21X1_809/A BUFX4_289/Y OAI21X1_809/C gnd OAI21X1_809/Y vdd OAI21X1
XOAI21X1_1111 OAI21X1_1111/A BUFX4_198/Y NAND2X1_475/Y gnd OAI21X1_1111/Y vdd OAI21X1
XOAI21X1_1100 INVX2_54/Y BUFX4_234/Y NAND2X1_466/Y gnd OAI21X1_1100/Y vdd OAI21X1
XOAI21X1_1122 XNOR2X1_56/Y BUFX4_231/Y NAND2X1_485/Y gnd OAI21X1_1122/Y vdd OAI21X1
XDFFPOSX1_701 BUFX2_339/A CLKBUF1_31/Y OAI21X1_951/Y gnd vdd DFFPOSX1
XOAI21X1_1155 NOR2X1_148/B INVX1_192/A BUFX4_238/Y gnd OAI21X1_1156/B vdd OAI21X1
XOAI21X1_1144 XNOR2X1_63/Y BUFX4_229/Y NAND2X1_516/Y gnd OAI21X1_1144/Y vdd OAI21X1
XFILL_1_OAI21X1_1342 gnd vdd FILL
XFILL_1_OAI21X1_1331 gnd vdd FILL
XFILL_1_OAI21X1_1320 gnd vdd FILL
XDFFPOSX1_712 BUFX2_357/A CLKBUF1_2/Y OAI21X1_973/Y gnd vdd DFFPOSX1
XDFFPOSX1_723 BUFX2_360/A CLKBUF1_92/Y OAI21X1_995/Y gnd vdd DFFPOSX1
XOAI21X1_1133 INVX1_187/Y OAI21X1_1133/B NAND2X1_503/Y gnd OAI21X1_1133/Y vdd OAI21X1
XFILL_0_OAI21X1_100 gnd vdd FILL
XDFFPOSX1_756 BUFX2_5/A CLKBUF1_65/Y OAI21X1_1048/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_111 gnd vdd FILL
XFILL_1_DFFPOSX1_943 gnd vdd FILL
XOAI21X1_1177 INVX2_102/A INVX1_195/A BUFX4_243/Y gnd OAI21X1_1178/B vdd OAI21X1
XFILL_1_OAI21X1_1375 gnd vdd FILL
XFILL_1_DFFPOSX1_932 gnd vdd FILL
XDFFPOSX1_745 BUFX2_2/A CLKBUF1_73/Y OAI21X1_1037/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_921 gnd vdd FILL
XFILL_1_OAI21X1_1353 gnd vdd FILL
XDFFPOSX1_734 BUFX2_372/A CLKBUF1_83/Y OAI21X1_1017/Y gnd vdd DFFPOSX1
XOAI21X1_1188 NOR3X1_14/C INVX4_48/Y INVX2_87/Y gnd NAND2X1_575/B vdd OAI21X1
XFILL_1_DFFPOSX1_910 gnd vdd FILL
XOAI21X1_1166 NAND2X1_547/Y NOR2X1_157/Y NAND2X1_545/Y gnd OAI21X1_1166/Y vdd OAI21X1
XFILL_1_OAI21X1_1364 gnd vdd FILL
XFILL_0_OAI21X1_133 gnd vdd FILL
XFILL_1_OAI21X1_1397 gnd vdd FILL
XFILL_1_DFFPOSX1_954 gnd vdd FILL
XDFFPOSX1_789 BUFX2_41/A CLKBUF1_68/Y OAI21X1_1081/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_315 gnd vdd FILL
XFILL_0_OAI21X1_122 gnd vdd FILL
XFILL_1_OAI21X1_1386 gnd vdd FILL
XFILL_0_OAI21X1_144 gnd vdd FILL
XFILL_1_DFFPOSX1_965 gnd vdd FILL
XDFFPOSX1_778 BUFX2_29/A CLKBUF1_49/Y OAI21X1_1070/Y gnd vdd DFFPOSX1
XOAI21X1_1199 OAI21X1_1199/A NOR2X1_174/Y NAND2X1_583/Y gnd OAI21X1_1199/Y vdd OAI21X1
XFILL_1_OAI21X1_326 gnd vdd FILL
XDFFPOSX1_767 BUFX2_17/A CLKBUF1_52/Y OAI21X1_1059/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_976 gnd vdd FILL
XFILL_0_OAI21X1_155 gnd vdd FILL
XFILL_1_OAI21X1_304 gnd vdd FILL
XFILL_0_OAI21X1_166 gnd vdd FILL
XFILL_1_DFFPOSX1_998 gnd vdd FILL
XFILL_19_15_1 gnd vdd FILL
XFILL_1_DFFPOSX1_987 gnd vdd FILL
XFILL_1_OAI21X1_337 gnd vdd FILL
XFILL_1_OAI21X1_348 gnd vdd FILL
XFILL_0_OAI21X1_188 gnd vdd FILL
XFILL_0_OAI21X1_177 gnd vdd FILL
XFILL_1_OAI21X1_359 gnd vdd FILL
XFILL_0_OAI21X1_199 gnd vdd FILL
XFILL_0_BUFX4_10 gnd vdd FILL
XFILL_32_17_1 gnd vdd FILL
XFILL_0_NAND3X1_19 gnd vdd FILL
XFILL_13_11_0 gnd vdd FILL
XFILL_0_BUFX4_43 gnd vdd FILL
XFILL_0_BUFX4_32 gnd vdd FILL
XFILL_0_BUFX4_54 gnd vdd FILL
XFILL_0_BUFX4_21 gnd vdd FILL
XFILL_0_BUFX4_65 gnd vdd FILL
XFILL_25_8_1 gnd vdd FILL
XFILL_0_BUFX4_87 gnd vdd FILL
XFILL_1_NAND2X1_332 gnd vdd FILL
XFILL_0_BUFX4_76 gnd vdd FILL
XFILL_0_NAND2X1_150 gnd vdd FILL
XFILL_0_8_1 gnd vdd FILL
XFILL_0_NAND2X1_161 gnd vdd FILL
XFILL_0_DFFPOSX1_500 gnd vdd FILL
XFILL_1_NAND2X1_354 gnd vdd FILL
XFILL_1_BUFX4_118 gnd vdd FILL
XFILL_1_BUFX4_107 gnd vdd FILL
XFILL_24_3_0 gnd vdd FILL
XFILL_0_BUFX4_98 gnd vdd FILL
XFILL_0_DFFPOSX1_533 gnd vdd FILL
XFILL_0_NAND2X1_172 gnd vdd FILL
XFILL_0_NAND2X1_194 gnd vdd FILL
XFILL_1_NAND2X1_365 gnd vdd FILL
XFILL_0_NAND2X1_183 gnd vdd FILL
XFILL_0_DFFPOSX1_522 gnd vdd FILL
XFILL_0_DFFPOSX1_511 gnd vdd FILL
XFILL_0_DFFPOSX1_544 gnd vdd FILL
XFILL_0_DFFPOSX1_555 gnd vdd FILL
XFILL_0_DFFPOSX1_566 gnd vdd FILL
XFILL_1_BUFX4_129 gnd vdd FILL
XFILL_1_NAND2X1_398 gnd vdd FILL
XFILL_1_NAND2X1_387 gnd vdd FILL
XFILL_0_DFFPOSX1_599 gnd vdd FILL
XFILL_0_DFFPOSX1_588 gnd vdd FILL
XFILL_0_DFFPOSX1_577 gnd vdd FILL
XFILL_5_DFFPOSX1_170 gnd vdd FILL
XFILL_5_DFFPOSX1_181 gnd vdd FILL
XFILL_5_DFFPOSX1_192 gnd vdd FILL
XFILL_0_OR2X2_13 gnd vdd FILL
XFILL_37_16_1 gnd vdd FILL
XFILL_8_9_1 gnd vdd FILL
XFILL_1_OAI21X1_882 gnd vdd FILL
XFILL_1_OAI21X1_860 gnd vdd FILL
XFILL_18_10_0 gnd vdd FILL
XNAND3X1_10 NOR2X1_11/Y NOR2X1_42/Y NOR2X1_30/Y gnd NOR3X1_4/C vdd NAND3X1
XNAND3X1_32 NOR2X1_105/Y NOR2X1_42/Y NOR2X1_30/Y gnd NOR3X1_8/C vdd NAND3X1
XNAND3X1_21 NOR2X1_19/Y NOR2X1_69/Y NOR2X1_74/Y gnd NOR2X1_82/B vdd NAND3X1
XFILL_1_OAI21X1_871 gnd vdd FILL
XFILL_7_4_0 gnd vdd FILL
XNAND3X1_54 bundleAddress_i[38] INVX1_204/Y NOR2X1_190/Y gnd XNOR2X1_79/A vdd NAND3X1
XNAND3X1_65 bundleAddress_i[29] AND2X2_31/B INVX1_223/Y gnd NAND3X1_65/Y vdd NAND3X1
XFILL_1_OAI21X1_893 gnd vdd FILL
XNAND3X1_43 bundleAddress_i[23] NOR2X1_158/Y NOR2X1_156/Y gnd XNOR2X1_71/A vdd NAND3X1
XFILL_31_12_0 gnd vdd FILL
XFILL_2_DFFPOSX1_605 gnd vdd FILL
XNOR2X1_21 bundleStartMajId_i[32] NOR2X1_21/B gnd NOR2X1_21/Y vdd NOR2X1
XBUFX2_703 BUFX2_703/A gnd pid2_o[2] vdd BUFX2
XNOR2X1_10 NOR2X1_10/A NOR2X1_10/B gnd AND2X2_2/B vdd NOR2X1
XBUFX2_736 BUFX2_736/A gnd pid3_o[28] vdd BUFX2
XBUFX2_714 BUFX2_714/A gnd pid3_o[30] vdd BUFX2
XBUFX2_725 BUFX2_725/A gnd pid3_o[29] vdd BUFX2
XFILL_3_DFFPOSX1_30 gnd vdd FILL
XFILL_3_DFFPOSX1_52 gnd vdd FILL
XNOR2X1_54 INVX4_25/Y INVX4_26/Y gnd INVX1_43/A vdd NOR2X1
XFILL_2_DFFPOSX1_627 gnd vdd FILL
XNOR2X1_43 INVX4_22/Y NOR3X1_4/C gnd NOR2X1_43/Y vdd NOR2X1
XNOR2X1_32 INVX4_17/Y NOR2X1_33/B gnd NOR2X1_32/Y vdd NOR2X1
XFILL_2_DFFPOSX1_616 gnd vdd FILL
XFILL_2_DFFPOSX1_638 gnd vdd FILL
XFILL_3_DFFPOSX1_41 gnd vdd FILL
XBUFX2_747 BUFX2_747/A gnd pid4_o[21] vdd BUFX2
XFILL_3_DFFPOSX1_85 gnd vdd FILL
XFILL_3_DFFPOSX1_63 gnd vdd FILL
XFILL_2_DFFPOSX1_649 gnd vdd FILL
XNOR2X1_76 OR2X2_6/B NOR2X1_76/B gnd NOR2X1_76/Y vdd NOR2X1
XFILL_16_8_1 gnd vdd FILL
XNOR2X1_87 INVX2_49/Y NOR2X1_87/B gnd INVX2_50/A vdd NOR2X1
XBUFX2_769 BUFX2_769/A gnd pid4_o[1] vdd BUFX2
XFILL_3_DFFPOSX1_74 gnd vdd FILL
XNOR2X1_65 bundleStartMajId_i[42] NOR2X1_65/B gnd NOR2X1_66/A vdd NOR2X1
XBUFX2_758 BUFX2_758/A gnd pid4_o[11] vdd BUFX2
XNOR2X1_98 bundleStartMajId_i[4] NOR2X1_98/B gnd NOR2X1_98/Y vdd NOR2X1
XFILL_3_DFFPOSX1_96 gnd vdd FILL
XFILL_15_3_0 gnd vdd FILL
XFILL_0_NOR2X1_109 gnd vdd FILL
XFILL_0_BUFX2_432 gnd vdd FILL
XFILL_0_BUFX2_421 gnd vdd FILL
XFILL_0_BUFX2_410 gnd vdd FILL
XFILL_1_DFFPOSX1_217 gnd vdd FILL
XFILL_1_DFFPOSX1_228 gnd vdd FILL
XFILL_0_BUFX2_443 gnd vdd FILL
XFILL_1_DFFPOSX1_206 gnd vdd FILL
XFILL_0_BUFX2_454 gnd vdd FILL
XFILL_0_BUFX2_465 gnd vdd FILL
XFILL_1_DFFPOSX1_239 gnd vdd FILL
XFILL_0_BUFX2_487 gnd vdd FILL
XFILL_0_BUFX2_498 gnd vdd FILL
XFILL_0_BUFX2_476 gnd vdd FILL
XFILL_36_11_0 gnd vdd FILL
XNAND2X1_9 NAND2X1_9/A OAI21X1_9/B gnd OAI21X1_9/C vdd NAND2X1
XNOR2X1_100 bundleStartMajId_i[2] AND2X2_17/Y gnd NOR2X1_100/Y vdd NOR2X1
XFILL_0_NAND2X1_30 gnd vdd FILL
XFILL_0_NAND2X1_52 gnd vdd FILL
XFILL_0_NAND2X1_41 gnd vdd FILL
XNOR2X1_122 bundleAddress_i[61] bundleAddress_i[60] gnd NOR2X1_215/B vdd NOR2X1
XNOR2X1_133 OR2X2_16/B NOR2X1_133/B gnd NOR2X1_133/Y vdd NOR2X1
XNOR2X1_111 INVX4_17/Y NOR2X1_112/B gnd XNOR2X1_50/A vdd NOR2X1
XFILL_0_NAND2X1_63 gnd vdd FILL
XFILL_0_NAND2X1_74 gnd vdd FILL
XNOR2X1_144 NOR2X1_144/A INVX1_190/A gnd XNOR2X1_65/A vdd NOR2X1
XNOR2X1_166 NOR2X1_166/A INVX1_224/A gnd AND2X2_24/B vdd NOR2X1
XNOR2X1_155 INVX1_208/A NOR2X1_155/B gnd INVX2_100/A vdd NOR2X1
XFILL_0_NAND2X1_85 gnd vdd FILL
XFILL_0_NAND2X1_96 gnd vdd FILL
XNOR2X1_177 bundleAddress_i[58] INVX1_183/Y gnd NOR2X1_177/Y vdd NOR2X1
XNOR2X1_188 bundleAddress_i[40] NOR2X1_188/B gnd NOR2X1_189/A vdd NOR2X1
XNOR2X1_199 bundleAddress_i[25] NOR2X1_199/B gnd NOR2X1_199/Y vdd NOR2X1
XOAI21X1_606 XNOR2X1_36/Y BUFX4_161/Y OAI21X1_606/C gnd OAI21X1_606/Y vdd OAI21X1
XOAI21X1_628 NOR2X1_93/Y OAI21X1_628/B OAI21X1_628/C gnd OAI21X1_628/Y vdd OAI21X1
XOAI21X1_639 OAI21X1_639/A INVX2_36/Y NOR2X1_96/B gnd OAI21X1_640/A vdd OAI21X1
XOAI21X1_617 OAI21X1_617/A NOR2X1_88/Y OAI21X1_617/C gnd OAI21X1_617/Y vdd OAI21X1
XFILL_1_OAI21X1_1150 gnd vdd FILL
XDFFPOSX1_520 BUFX2_551/A CLKBUF1_9/Y OAI21X1_596/Y gnd vdd DFFPOSX1
XDFFPOSX1_531 BUFX2_563/A CLKBUF1_90/Y OAI21X1_623/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_101 gnd vdd FILL
XFILL_1_DFFPOSX1_751 gnd vdd FILL
XFILL_1_DFFPOSX1_740 gnd vdd FILL
XDFFPOSX1_542 BUFX2_575/A CLKBUF1_72/Y OAI21X1_646/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1172 gnd vdd FILL
XFILL_1_OAI21X1_1161 gnd vdd FILL
XDFFPOSX1_564 BUFX2_593/A CLKBUF1_79/Y OAI21X1_706/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1183 gnd vdd FILL
XDFFPOSX1_553 BUFX2_630/A CLKBUF1_41/Y OAI21X1_675/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_112 gnd vdd FILL
XFILL_1_DFFPOSX1_773 gnd vdd FILL
XFILL_1_OAI21X1_123 gnd vdd FILL
XFILL_1_DFFPOSX1_762 gnd vdd FILL
XFILL_1_OAI21X1_134 gnd vdd FILL
XDFFPOSX1_575 BUFX2_605/A CLKBUF1_1/Y OAI21X1_738/Y gnd vdd DFFPOSX1
XDFFPOSX1_586 INVX1_42/A CLKBUF1_88/Y OAI21X1_767/Y gnd vdd DFFPOSX1
XNAND2X1_601 AND2X2_27/A NAND2X1_601/B gnd NAND2X1_601/Y vdd NAND2X1
XDFFPOSX1_597 BUFX2_629/A CLKBUF1_79/Y OAI21X1_801/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1194 gnd vdd FILL
XNAND2X1_612 INVX2_101/Y AND2X2_31/Y gnd NAND2X1_612/Y vdd NAND2X1
XFILL_1_DFFPOSX1_784 gnd vdd FILL
XFILL_2_OAI21X1_305 gnd vdd FILL
XFILL_1_OAI21X1_167 gnd vdd FILL
XNAND2X1_634 XNOR2X1_99/A NAND2X1_634/B gnd NAND2X1_634/Y vdd NAND2X1
XNAND2X1_623 BUFX4_310/Y INVX1_217/A gnd NAND2X1_623/Y vdd NAND2X1
XFILL_1_OAI21X1_145 gnd vdd FILL
XNAND2X1_645 bundleAddress_i[5] NOR2X1_231/Y gnd INVX2_112/A vdd NAND2X1
XINVX1_13 INVX1_13/A gnd NOR3X1_1/B vdd INVX1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XFILL_1_OAI21X1_156 gnd vdd FILL
XFILL_1_DFFPOSX1_795 gnd vdd FILL
XNAND2X1_667 BUFX2_658/A BUFX4_380/Y gnd NAND2X1_667/Y vdd NAND2X1
XNAND2X1_678 BUFX2_670/A BUFX4_368/Y gnd NAND2X1_678/Y vdd NAND2X1
XFILL_1_OAI21X1_178 gnd vdd FILL
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XINVX1_57 INVX1_57/A gnd INVX1_57/Y vdd INVX1
XFILL_1_OAI21X1_189 gnd vdd FILL
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XNAND2X1_656 BUFX2_677/A OAI21X1_6/A gnd NAND2X1_656/Y vdd NAND2X1
XNAND2X1_689 BUFX2_710/A BUFX4_207/Y gnd NAND2X1_689/Y vdd NAND2X1
XINVX1_68 INVX1_68/A gnd INVX1_68/Y vdd INVX1
XINVX1_79 bundle_i[61] gnd INVX1_79/Y vdd INVX1
XDFFPOSX1_9 BUFX2_708/A CLKBUF1_58/Y DFFPOSX1_9/D gnd vdd DFFPOSX1
XFILL_0_DFFPOSX1_330 gnd vdd FILL
XFILL_0_DFFPOSX1_341 gnd vdd FILL
XFILL_1_NAND2X1_151 gnd vdd FILL
XFILL_0_DFFPOSX1_374 gnd vdd FILL
XFILL_0_DFFPOSX1_352 gnd vdd FILL
XFILL_1_NAND2X1_195 gnd vdd FILL
XFILL_1_NAND2X1_184 gnd vdd FILL
XFILL_0_DFFPOSX1_363 gnd vdd FILL
XFILL_0_DFFPOSX1_396 gnd vdd FILL
XFILL_0_DFFPOSX1_385 gnd vdd FILL
XFILL_3_DFFPOSX1_812 gnd vdd FILL
XFILL_3_DFFPOSX1_823 gnd vdd FILL
XFILL_3_DFFPOSX1_801 gnd vdd FILL
XFILL_3_DFFPOSX1_856 gnd vdd FILL
XFILL_3_DFFPOSX1_834 gnd vdd FILL
XFILL_3_DFFPOSX1_845 gnd vdd FILL
XFILL_3_DFFPOSX1_889 gnd vdd FILL
XFILL_3_DFFPOSX1_878 gnd vdd FILL
XFILL_3_DFFPOSX1_867 gnd vdd FILL
XFILL_2_OAI21X1_861 gnd vdd FILL
XFILL_1_OAI21X1_690 gnd vdd FILL
XFILL_1_INVX1_140 gnd vdd FILL
XFILL_2_OAI21X1_894 gnd vdd FILL
XBUFX2_511 BUFX2_511/A gnd majID2_o[5] vdd BUFX2
XFILL_2_DFFPOSX1_413 gnd vdd FILL
XBUFX2_500 BUFX2_500/A gnd majID2_o[15] vdd BUFX2
XFILL_2_DFFPOSX1_402 gnd vdd FILL
XFILL_4_DFFPOSX1_20 gnd vdd FILL
XBUFX2_533 BUFX2_533/A gnd majID3_o[61] vdd BUFX2
XFILL_4_DFFPOSX1_31 gnd vdd FILL
XFILL_2_DFFPOSX1_424 gnd vdd FILL
XFILL_2_DFFPOSX1_435 gnd vdd FILL
XFILL_2_DFFPOSX1_446 gnd vdd FILL
XBUFX2_544 BUFX2_544/A gnd majID3_o[60] vdd BUFX2
XBUFX2_522 BUFX2_522/A gnd majID3_o[62] vdd BUFX2
XFILL_4_DFFPOSX1_42 gnd vdd FILL
XFILL_4_DFFPOSX1_75 gnd vdd FILL
XFILL_4_DFFPOSX1_53 gnd vdd FILL
XFILL_2_DFFPOSX1_479 gnd vdd FILL
XFILL_4_DFFPOSX1_64 gnd vdd FILL
XFILL_2_DFFPOSX1_468 gnd vdd FILL
XFILL_2_DFFPOSX1_457 gnd vdd FILL
XBUFX2_588 BUFX2_588/A gnd majID4_o[52] vdd BUFX2
XBUFX2_555 BUFX2_555/A gnd majID3_o[59] vdd BUFX2
XBUFX2_577 BUFX2_577/A gnd majID3_o[57] vdd BUFX2
XBUFX2_566 BUFX2_566/A gnd majID3_o[58] vdd BUFX2
XFILL_4_DFFPOSX1_86 gnd vdd FILL
XFILL_4_DFFPOSX1_97 gnd vdd FILL
XBUFX2_599 BUFX2_599/A gnd majID4_o[42] vdd BUFX2
XFILL_31_6_1 gnd vdd FILL
XFILL_5_DFFPOSX1_906 gnd vdd FILL
XFILL_5_DFFPOSX1_917 gnd vdd FILL
XFILL_5_DFFPOSX1_928 gnd vdd FILL
XFILL_5_DFFPOSX1_939 gnd vdd FILL
XFILL_30_1_0 gnd vdd FILL
XFILL_22_17_0 gnd vdd FILL
XFILL_0_BUFX2_240 gnd vdd FILL
XFILL_0_BUFX2_251 gnd vdd FILL
XFILL_0_BUFX2_262 gnd vdd FILL
XFILL_0_AND2X2_8 gnd vdd FILL
XFILL_0_BUFX2_273 gnd vdd FILL
XFILL_2_AND2X2_22 gnd vdd FILL
XFILL_0_BUFX2_295 gnd vdd FILL
XFILL_0_BUFX2_284 gnd vdd FILL
XFILL_4_DFFPOSX1_507 gnd vdd FILL
XFILL_4_DFFPOSX1_518 gnd vdd FILL
XFILL_4_DFFPOSX1_529 gnd vdd FILL
XFILL_38_2_0 gnd vdd FILL
XFILL_1_BUFX2_1009 gnd vdd FILL
XFILL_2_DFFPOSX1_980 gnd vdd FILL
XFILL_2_DFFPOSX1_991 gnd vdd FILL
XFILL_22_6_1 gnd vdd FILL
XFILL_1_BUFX2_408 gnd vdd FILL
XFILL_27_16_0 gnd vdd FILL
XFILL_21_1_0 gnd vdd FILL
XFILL_0_NAND3X1_3 gnd vdd FILL
XOAI21X1_414 NOR2X1_6/B OR2X2_1/A OAI21X1_414/C gnd OAI21X1_415/A vdd OAI21X1
XOAI21X1_403 INVX2_40/Y NOR2X1_4/A OAI21X1_403/C gnd OAI21X1_404/A vdd OAI21X1
XFILL_1_BUFX2_419 gnd vdd FILL
XOAI21X1_447 INVX1_14/Y BUFX4_245/Y OAI21X1_447/C gnd OAI21X1_447/Y vdd OAI21X1
XFILL_3_DFFPOSX1_108 gnd vdd FILL
XOAI21X1_436 OAI21X1_436/A NOR2X1_17/Y OAI21X1_436/C gnd OAI21X1_436/Y vdd OAI21X1
XOAI21X1_425 XNOR2X1_6/Y BUFX4_221/Y OAI21X1_425/C gnd OAI21X1_425/Y vdd OAI21X1
XFILL_3_DFFPOSX1_119 gnd vdd FILL
XOAI21X1_458 INVX1_17/Y bundleStartMajId_i[23] BUFX4_241/Y gnd OAI21X1_459/A vdd OAI21X1
XOAI21X1_469 OAI21X1_469/A AND2X2_8/Y OAI21X1_469/C gnd OAI21X1_469/Y vdd OAI21X1
XFILL_3_XNOR2X1_60 gnd vdd FILL
XFILL_3_XNOR2X1_93 gnd vdd FILL
XFILL_3_XNOR2X1_71 gnd vdd FILL
XDFFPOSX1_350 BUFX2_1023/A CLKBUF1_92/Y OAI21X1_317/Y gnd vdd DFFPOSX1
XDFFPOSX1_361 BUFX2_438/A CLKBUF1_66/Y OAI21X1_333/Y gnd vdd DFFPOSX1
XDFFPOSX1_372 BUFX2_401/A CLKBUF1_75/Y OAI21X1_344/Y gnd vdd DFFPOSX1
XDFFPOSX1_383 BUFX2_413/A CLKBUF1_33/Y OAI21X1_355/Y gnd vdd DFFPOSX1
XDFFPOSX1_394 BUFX2_425/A CLKBUF1_19/Y OAI21X1_366/Y gnd vdd DFFPOSX1
XNAND2X1_420 BUFX2_11/A BUFX4_311/Y gnd NAND2X1_420/Y vdd NAND2X1
XFILL_1_DFFPOSX1_592 gnd vdd FILL
XFILL_1_DFFPOSX1_570 gnd vdd FILL
XFILL_1_DFFPOSX1_581 gnd vdd FILL
XNAND2X1_431 BUFX2_23/A BUFX4_377/Y gnd NAND2X1_431/Y vdd NAND2X1
XNAND2X1_442 BUFX2_36/A BUFX4_350/Y gnd NAND2X1_442/Y vdd NAND2X1
XNAND2X1_453 BUFX2_48/A BUFX4_364/Y gnd NAND2X1_453/Y vdd NAND2X1
XNAND2X1_475 BUFX2_121/A BUFX4_198/Y gnd NAND2X1_475/Y vdd NAND2X1
XFILL_2_OAI21X1_168 gnd vdd FILL
XNAND2X1_486 BUFX2_69/A BUFX4_231/Y gnd NAND2X1_486/Y vdd NAND2X1
XNAND2X1_497 bundleAddress_i[49] bundleAddress_i[48] gnd OR2X2_16/B vdd NAND2X1
XNAND2X1_464 BUFX2_60/A BUFX4_339/Y gnd NAND2X1_464/Y vdd NAND2X1
XFILL_5_7_1 gnd vdd FILL
XFILL_29_2_0 gnd vdd FILL
XFILL_4_2_0 gnd vdd FILL
XFILL_0_INVX1_207 gnd vdd FILL
XFILL_0_INVX1_218 gnd vdd FILL
XFILL_2_17_0 gnd vdd FILL
XFILL_13_6_1 gnd vdd FILL
XFILL_0_DFFPOSX1_171 gnd vdd FILL
XFILL_0_DFFPOSX1_182 gnd vdd FILL
XFILL_1_BUFX2_920 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XFILL_0_DFFPOSX1_160 gnd vdd FILL
XFILL_1_BUFX2_931 gnd vdd FILL
XFILL_0_DFFPOSX1_193 gnd vdd FILL
XFILL_0_OAI21X1_39 gnd vdd FILL
XFILL_0_OAI21X1_17 gnd vdd FILL
XFILL_1_BUFX2_964 gnd vdd FILL
XFILL_1_BUFX2_942 gnd vdd FILL
XFILL_0_OAI21X1_28 gnd vdd FILL
XFILL_1_BUFX2_975 gnd vdd FILL
XFILL_1_BUFX2_986 gnd vdd FILL
XOAI21X1_970 BUFX4_106/Y BUFX4_318/Y BUFX2_350/A gnd OAI21X1_971/C vdd OAI21X1
XFILL_3_DFFPOSX1_620 gnd vdd FILL
XFILL_3_DFFPOSX1_631 gnd vdd FILL
XFILL_3_DFFPOSX1_664 gnd vdd FILL
XOAI21X1_992 BUFX4_136/Y BUFX4_75/Y BUFX2_359/A gnd OAI21X1_993/C vdd OAI21X1
XOAI21X1_981 BUFX4_293/Y INVX1_145/Y OAI21X1_981/C gnd OAI21X1_981/Y vdd OAI21X1
XFILL_3_DFFPOSX1_642 gnd vdd FILL
XFILL_3_DFFPOSX1_653 gnd vdd FILL
XFILL_3_DFFPOSX1_675 gnd vdd FILL
XFILL_3_DFFPOSX1_697 gnd vdd FILL
XFILL_3_DFFPOSX1_686 gnd vdd FILL
XFILL_7_16_0 gnd vdd FILL
XFILL_2_OAI21X1_680 gnd vdd FILL
XFILL_0_NAND2X1_705 gnd vdd FILL
XFILL_0_NAND2X1_727 gnd vdd FILL
XFILL_2_DFFPOSX1_221 gnd vdd FILL
XFILL_2_DFFPOSX1_210 gnd vdd FILL
XFILL_0_NAND2X1_716 gnd vdd FILL
XFILL_0_NAND2X1_749 gnd vdd FILL
XFILL_5_DFFPOSX1_21 gnd vdd FILL
XFILL_2_DFFPOSX1_232 gnd vdd FILL
XFILL_2_DFFPOSX1_254 gnd vdd FILL
XFILL_2_DFFPOSX1_243 gnd vdd FILL
XFILL_2_DFFPOSX1_265 gnd vdd FILL
XFILL_0_NAND2X1_738 gnd vdd FILL
XFILL_0_OAI21X1_1509 gnd vdd FILL
XFILL_11_14_1 gnd vdd FILL
XBUFX2_330 BUFX2_330/A gnd instr3_o[18] vdd BUFX2
XBUFX2_363 BUFX2_363/A gnd instr4_o[17] vdd BUFX2
XBUFX2_341 BUFX2_341/A gnd instr3_o[8] vdd BUFX2
XBUFX2_352 BUFX2_352/A gnd instr3_o[26] vdd BUFX2
XFILL_5_DFFPOSX1_10 gnd vdd FILL
XBUFX2_385 BUFX2_385/A gnd instr4_o[25] vdd BUFX2
XFILL_5_DFFPOSX1_32 gnd vdd FILL
XFILL_5_DFFPOSX1_43 gnd vdd FILL
XBUFX2_374 BUFX2_374/A gnd instr4_o[7] vdd BUFX2
XFILL_2_DFFPOSX1_276 gnd vdd FILL
XFILL_5_DFFPOSX1_54 gnd vdd FILL
XFILL_2_DFFPOSX1_298 gnd vdd FILL
XBUFX2_396 BUFX2_396/A gnd majID1_o[52] vdd BUFX2
XFILL_2_DFFPOSX1_287 gnd vdd FILL
XFILL_5_DFFPOSX1_76 gnd vdd FILL
XFILL_5_DFFPOSX1_87 gnd vdd FILL
XFILL_5_DFFPOSX1_65 gnd vdd FILL
XFILL_1_NOR3X1_13 gnd vdd FILL
XFILL_5_DFFPOSX1_703 gnd vdd FILL
XFILL_5_DFFPOSX1_98 gnd vdd FILL
XOAI21X1_52 INVX2_190/Y BUFX4_191/Y OAI21X1_52/C gnd OAI21X1_52/Y vdd OAI21X1
XFILL_5_DFFPOSX1_725 gnd vdd FILL
XOAI21X1_41 INVX2_179/Y BUFX4_208/Y OAI21X1_41/C gnd OAI21X1_41/Y vdd OAI21X1
XFILL_5_DFFPOSX1_736 gnd vdd FILL
XOAI21X1_30 INVX2_168/Y BUFX4_195/Y OAI21X1_30/C gnd OAI21X1_30/Y vdd OAI21X1
XFILL_5_DFFPOSX1_714 gnd vdd FILL
XOAI21X1_63 INVX2_201/Y BUFX4_180/Y OAI21X1_63/C gnd OAI21X1_63/Y vdd OAI21X1
XOAI21X1_96 BUFX4_11/A BUFX4_322/Y BUFX2_909/A gnd OAI21X1_97/C vdd OAI21X1
XFILL_5_DFFPOSX1_747 gnd vdd FILL
XFILL_5_DFFPOSX1_758 gnd vdd FILL
XOAI21X1_85 BUFX4_170/Y INVX2_152/Y OAI21X1_85/C gnd OAI21X1_85/Y vdd OAI21X1
XOAI21X1_74 BUFX4_106/Y BUFX4_318/Y BUFX2_906/A gnd OAI21X1_75/C vdd OAI21X1
XFILL_1_BUFX4_290 gnd vdd FILL
XFILL_5_DFFPOSX1_769 gnd vdd FILL
XFILL_4_DFFPOSX1_304 gnd vdd FILL
XFILL_0_DFFPOSX1_50 gnd vdd FILL
XFILL_4_DFFPOSX1_326 gnd vdd FILL
XFILL_4_DFFPOSX1_315 gnd vdd FILL
XFILL_0_DFFPOSX1_61 gnd vdd FILL
XFILL_16_13_1 gnd vdd FILL
XFILL_4_DFFPOSX1_337 gnd vdd FILL
XFILL_0_DFFPOSX1_94 gnd vdd FILL
XFILL_4_DFFPOSX1_348 gnd vdd FILL
XFILL_0_DFFPOSX1_83 gnd vdd FILL
XFILL_0_DFFPOSX1_72 gnd vdd FILL
XFILL_4_DFFPOSX1_359 gnd vdd FILL
XFILL_2_DFFPOSX1_1018 gnd vdd FILL
XFILL_2_DFFPOSX1_1007 gnd vdd FILL
XFILL_2_DFFPOSX1_1029 gnd vdd FILL
XFILL_1_BUFX2_216 gnd vdd FILL
XFILL_1_BUFX2_205 gnd vdd FILL
XFILL_1_BUFX2_227 gnd vdd FILL
XFILL_1_BUFX2_249 gnd vdd FILL
XOAI21X1_222 BUFX4_148/Y BUFX4_35/Y BUFX2_972/A gnd OAI21X1_223/C vdd OAI21X1
XOAI21X1_200 BUFX4_149/Y BUFX4_79/Y BUFX2_969/A gnd OAI21X1_201/C vdd OAI21X1
XOAI21X1_211 INVX2_151/Y BUFX4_303/Y OAI21X1_211/C gnd OAI21X1_211/Y vdd OAI21X1
XOAI21X1_255 INVX2_173/Y BUFX4_293/Y OAI21X1_255/C gnd OAI21X1_255/Y vdd OAI21X1
XOAI21X1_233 INVX2_162/Y BUFX4_295/Y OAI21X1_233/C gnd OAI21X1_233/Y vdd OAI21X1
XOAI21X1_244 BUFX4_162/Y BUFX4_51/Y BUFX2_984/A gnd OAI21X1_245/C vdd OAI21X1
XOAI21X1_277 INVX2_184/Y BUFX4_293/Y OAI21X1_277/C gnd OAI21X1_277/Y vdd OAI21X1
XOAI21X1_299 INVX2_195/Y BUFX4_293/Y OAI21X1_299/C gnd OAI21X1_299/Y vdd OAI21X1
XOAI21X1_288 BUFX4_159/Y BUFX4_67/A BUFX2_1008/A gnd OAI21X1_289/C vdd OAI21X1
XOAI21X1_266 BUFX4_151/Y BUFX4_70/Y BUFX2_996/A gnd OAI21X1_267/C vdd OAI21X1
XAND2X2_22 AND2X2_22/A INVX2_31/Y gnd AND2X2_22/Y vdd AND2X2
XAND2X2_11 NOR2X1_59/Y NOR2X1_60/Y gnd INVX4_30/A vdd AND2X2
XAND2X2_33 INVX2_107/Y AND2X2_33/B gnd AND2X2_33/Y vdd AND2X2
XDFFPOSX1_191 BUFX2_861/A CLKBUF1_17/Y OAI21X1_35/Y gnd vdd DFFPOSX1
XDFFPOSX1_180 BUFX2_849/A CLKBUF1_43/Y OAI21X1_24/Y gnd vdd DFFPOSX1
XFILL_0_NOR3X1_1 gnd vdd FILL
XFILL_34_14_1 gnd vdd FILL
XNAND2X1_261 BUFX2_515/A BUFX4_221/Y gnd OAI21X1_496/C vdd NAND2X1
XNAND2X1_250 bundleStartMajId_i[7] NOR2X1_52/Y gnd INVX1_22/A vdd NAND2X1
XNAND2X1_294 INVX2_48/A NOR2X1_83/Y gnd INVX1_31/A vdd NAND2X1
XNAND2X1_283 bundleStartMajId_i[36] INVX2_42/Y gnd OAI21X1_575/B vdd NAND2X1
XNAND2X1_272 bundleStartMajId_i[52] INVX1_9/Y gnd NOR2X1_104/A vdd NAND2X1
XFILL_4_DFFPOSX1_882 gnd vdd FILL
XFILL_4_DFFPOSX1_871 gnd vdd FILL
XFILL_4_DFFPOSX1_860 gnd vdd FILL
XFILL_4_DFFPOSX1_893 gnd vdd FILL
XFILL_0_INVX8_7 gnd vdd FILL
XFILL_2_XNOR2X1_100 gnd vdd FILL
XFILL_0_BUFX4_313 gnd vdd FILL
XFILL_0_BUFX4_302 gnd vdd FILL
XFILL_0_BUFX4_324 gnd vdd FILL
XFILL_1_NOR2X1_90 gnd vdd FILL
XFILL_1_BUFX2_772 gnd vdd FILL
XFILL_1_BUFX2_783 gnd vdd FILL
XOAI21X1_1529 INVX1_225/A INVX1_195/A BUFX4_284/Y gnd OAI21X1_1530/B vdd OAI21X1
XOAI21X1_1518 INVX2_110/Y NOR2X1_204/A INVX2_81/Y gnd OAI21X1_1519/C vdd OAI21X1
XFILL_1_OAI21X1_1716 gnd vdd FILL
XFILL_0_BUFX4_346 gnd vdd FILL
XFILL_0_BUFX4_357 gnd vdd FILL
XOAI21X1_1507 INVX1_224/A INVX1_223/A OAI21X1_1507/C gnd OAI21X1_1509/A vdd OAI21X1
XFILL_1_OAI21X1_1705 gnd vdd FILL
XFILL_0_BUFX4_335 gnd vdd FILL
XFILL_1_OAI21X1_1727 gnd vdd FILL
XFILL_3_DFFPOSX1_483 gnd vdd FILL
XFILL_0_BUFX4_368 gnd vdd FILL
XFILL_1_OAI21X1_1738 gnd vdd FILL
XFILL_0_BUFX4_379 gnd vdd FILL
XFILL_3_DFFPOSX1_450 gnd vdd FILL
XFILL_1_OAI21X1_1749 gnd vdd FILL
XFILL_3_DFFPOSX1_461 gnd vdd FILL
XFILL_3_DFFPOSX1_472 gnd vdd FILL
XFILL_0_OAI21X1_507 gnd vdd FILL
XFILL_3_DFFPOSX1_494 gnd vdd FILL
XFILL_0_OAI21X1_529 gnd vdd FILL
XFILL_0_BUFX2_1006 gnd vdd FILL
XFILL_0_OAI21X1_518 gnd vdd FILL
XFILL_6_DFFPOSX1_921 gnd vdd FILL
XFILL_6_DFFPOSX1_910 gnd vdd FILL
XFILL_0_BUFX2_1017 gnd vdd FILL
XFILL_0_BUFX2_1028 gnd vdd FILL
XFILL_6_DFFPOSX1_954 gnd vdd FILL
XFILL_6_DFFPOSX1_943 gnd vdd FILL
XFILL_6_DFFPOSX1_932 gnd vdd FILL
XFILL_6_1 gnd vdd FILL
XFILL_6_DFFPOSX1_965 gnd vdd FILL
XFILL_0_CLKBUF1_18 gnd vdd FILL
XFILL_0_CLKBUF1_29 gnd vdd FILL
XFILL_0_NAND2X1_502 gnd vdd FILL
XFILL_36_5_1 gnd vdd FILL
XFILL_0_NAND2X1_524 gnd vdd FILL
XFILL_0_NAND2X1_513 gnd vdd FILL
XFILL_0_OAI21X1_1306 gnd vdd FILL
XFILL_0_NAND2X1_535 gnd vdd FILL
XFILL_35_0_0 gnd vdd FILL
XBUFX2_171 BUFX2_171/A gnd addr3_o[16] vdd BUFX2
XFILL_2_XNOR2X1_90 gnd vdd FILL
XFILL_0_OAI21X1_1339 gnd vdd FILL
XFILL_0_NAND2X1_557 gnd vdd FILL
XFILL_0_OAI21X1_1328 gnd vdd FILL
XFILL_0_NAND2X1_568 gnd vdd FILL
XFILL_1_NAND2X1_717 gnd vdd FILL
XFILL_1_NAND2X1_728 gnd vdd FILL
XFILL_0_NAND2X1_546 gnd vdd FILL
XFILL_0_OAI21X1_1317 gnd vdd FILL
XFILL_0_DFFPOSX1_907 gnd vdd FILL
XBUFX2_160 BUFX2_160/A gnd addr3_o[26] vdd BUFX2
XFILL_6_DFFPOSX1_11 gnd vdd FILL
XBUFX2_193 BUFX2_193/A gnd addr4_o[63] vdd BUFX2
XFILL_6_DFFPOSX1_44 gnd vdd FILL
XFILL_6_DFFPOSX1_22 gnd vdd FILL
XFILL_0_DFFPOSX1_918 gnd vdd FILL
XFILL_0_DFFPOSX1_929 gnd vdd FILL
XBUFX2_182 BUFX2_182/A gnd addr3_o[6] vdd BUFX2
XFILL_6_DFFPOSX1_33 gnd vdd FILL
XFILL_0_NAND2X1_579 gnd vdd FILL
XFILL_6_DFFPOSX1_55 gnd vdd FILL
XFILL_5_DFFPOSX1_500 gnd vdd FILL
XFILL_5_DFFPOSX1_511 gnd vdd FILL
XFILL_5_DFFPOSX1_544 gnd vdd FILL
XFILL_5_DFFPOSX1_533 gnd vdd FILL
XFILL_5_DFFPOSX1_522 gnd vdd FILL
XFILL_5_DFFPOSX1_555 gnd vdd FILL
XFILL_5_DFFPOSX1_588 gnd vdd FILL
XFILL_5_DFFPOSX1_566 gnd vdd FILL
XFILL_5_DFFPOSX1_577 gnd vdd FILL
XFILL_5_DFFPOSX1_599 gnd vdd FILL
XBUFX2_1030 BUFX2_1030/A gnd tid4_o[56] vdd BUFX2
XFILL_1_AOI21X1_6 gnd vdd FILL
XCLKBUF1_42 BUFX4_87/Y gnd CLKBUF1_42/Y vdd CLKBUF1
XCLKBUF1_31 BUFX4_85/Y gnd CLKBUF1_31/Y vdd CLKBUF1
XCLKBUF1_20 BUFX4_89/Y gnd CLKBUF1_20/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_101 gnd vdd FILL
XFILL_4_DFFPOSX1_134 gnd vdd FILL
XFILL_4_DFFPOSX1_145 gnd vdd FILL
XFILL_4_DFFPOSX1_112 gnd vdd FILL
XFILL_1_DFFPOSX1_51 gnd vdd FILL
XFILL_4_DFFPOSX1_123 gnd vdd FILL
XCLKBUF1_64 BUFX4_83/Y gnd CLKBUF1_64/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_40 gnd vdd FILL
XCLKBUF1_75 BUFX4_90/Y gnd CLKBUF1_75/Y vdd CLKBUF1
XCLKBUF1_53 BUFX4_88/Y gnd CLKBUF1_53/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_178 gnd vdd FILL
XFILL_4_DFFPOSX1_156 gnd vdd FILL
XFILL_1_DFFPOSX1_84 gnd vdd FILL
XFILL_1_DFFPOSX1_62 gnd vdd FILL
XCLKBUF1_86 BUFX4_92/Y gnd CLKBUF1_86/Y vdd CLKBUF1
XCLKBUF1_97 BUFX4_87/Y gnd CLKBUF1_97/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_73 gnd vdd FILL
XFILL_4_DFFPOSX1_167 gnd vdd FILL
XFILL_4_DFFPOSX1_189 gnd vdd FILL
XFILL_1_DFFPOSX1_95 gnd vdd FILL
XFILL_27_5_1 gnd vdd FILL
XFILL_2_BUFX4_222 gnd vdd FILL
XFILL_2_5_1 gnd vdd FILL
XFILL_26_0_0 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XFILL_10_4_1 gnd vdd FILL
XFILL_0_BUFX2_806 gnd vdd FILL
XFILL_0_BUFX2_817 gnd vdd FILL
XFILL_0_BUFX2_828 gnd vdd FILL
XINVX1_116 bundle_i[88] gnd INVX1_116/Y vdd INVX1
XINVX1_105 bundle_i[35] gnd INVX1_105/Y vdd INVX1
XFILL_0_BUFX2_839 gnd vdd FILL
XINVX1_127 bundle_i[77] gnd INVX1_127/Y vdd INVX1
XINVX1_149 bundle_i[119] gnd INVX1_149/Y vdd INVX1
XINVX1_138 bundle_i[66] gnd INVX1_138/Y vdd INVX1
XFILL_6_DFFPOSX1_217 gnd vdd FILL
XFILL_6_DFFPOSX1_206 gnd vdd FILL
XFILL_6_DFFPOSX1_239 gnd vdd FILL
XFILL_6_DFFPOSX1_228 gnd vdd FILL
XFILL_9_1_0 gnd vdd FILL
XFILL_0_INVX2_37 gnd vdd FILL
XFILL_0_INVX2_26 gnd vdd FILL
XFILL_0_INVX2_15 gnd vdd FILL
XFILL_0_INVX2_59 gnd vdd FILL
XFILL_0_INVX2_48 gnd vdd FILL
XFILL_4_DFFPOSX1_690 gnd vdd FILL
XFILL_18_5_1 gnd vdd FILL
XFILL_0_CLKBUF1_5 gnd vdd FILL
XFILL_17_0_0 gnd vdd FILL
XFILL_3_XNOR2X1_101 gnd vdd FILL
XFILL_1_BUFX2_580 gnd vdd FILL
XFILL_0_BUFX4_110 gnd vdd FILL
XFILL_0_BUFX4_132 gnd vdd FILL
XFILL_0_BUFX4_121 gnd vdd FILL
XFILL_1_BUFX2_591 gnd vdd FILL
XOAI21X1_1304 BUFX4_6/Y BUFX4_350/Y BUFX2_158/A gnd OAI21X1_1305/C vdd OAI21X1
XFILL_0_BUFX4_165 gnd vdd FILL
XFILL_1_BUFX2_10 gnd vdd FILL
XFILL_0_BUFX4_143 gnd vdd FILL
XFILL_1_INVX1_90 gnd vdd FILL
XFILL_1_BUFX2_21 gnd vdd FILL
XOAI21X1_1337 INVX1_212/A INVX2_82/Y BUFX4_310/Y gnd OAI21X1_1338/B vdd OAI21X1
XFILL_1_OAI21X1_1524 gnd vdd FILL
XDFFPOSX1_905 BUFX2_156/A CLKBUF1_49/Y OAI21X1_1299/Y gnd vdd DFFPOSX1
XOAI21X1_1326 BUFX4_6/A BUFX4_344/Y BUFX2_167/A gnd OAI21X1_1327/C vdd OAI21X1
XFILL_1_OAI21X1_1513 gnd vdd FILL
XFILL_0_BUFX4_176 gnd vdd FILL
XOAI21X1_1315 XNOR2X1_84/Y BUFX4_169/Y OAI21X1_1315/C gnd OAI21X1_1315/Y vdd OAI21X1
XFILL_0_BUFX4_154 gnd vdd FILL
XFILL_1_OAI21X1_1502 gnd vdd FILL
XFILL_0_BUFX4_198 gnd vdd FILL
XDFFPOSX1_938 BUFX2_205/A CLKBUF1_91/Y OAI21X1_1389/Y gnd vdd DFFPOSX1
XDFFPOSX1_916 BUFX2_168/A CLKBUF1_68/Y OAI21X1_1330/Y gnd vdd DFFPOSX1
XFILL_0_BUFX4_187 gnd vdd FILL
XFILL_3_DFFPOSX1_291 gnd vdd FILL
XDFFPOSX1_927 BUFX2_180/A CLKBUF1_69/Y OAI21X1_1360/Y gnd vdd DFFPOSX1
XOAI21X1_1359 INVX1_215/A INVX4_45/Y BUFX4_308/Y gnd OAI21X1_1360/B vdd OAI21X1
XFILL_1_OAI21X1_1557 gnd vdd FILL
XOAI21X1_1348 BUFX4_6/Y NAND2X1_7/B BUFX2_176/A gnd OAI21X1_1349/C vdd OAI21X1
XFILL_1_OAI21X1_1546 gnd vdd FILL
XFILL_1_BUFX2_54 gnd vdd FILL
XFILL_1_OAI21X1_1535 gnd vdd FILL
XFILL_1_BUFX2_32 gnd vdd FILL
XFILL_3_DFFPOSX1_280 gnd vdd FILL
XFILL_0_OAI21X1_304 gnd vdd FILL
XFILL_1_BUFX2_65 gnd vdd FILL
XDFFPOSX1_949 BUFX2_198/A CLKBUF1_5/Y OAI21X1_1424/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_315 gnd vdd FILL
XFILL_1_OAI21X1_1568 gnd vdd FILL
XFILL_1_OAI21X1_1579 gnd vdd FILL
XFILL_1_OAI21X1_508 gnd vdd FILL
XFILL_0_OAI21X1_337 gnd vdd FILL
XFILL_1_BUFX2_76 gnd vdd FILL
XFILL_0_OAI21X1_326 gnd vdd FILL
XFILL_0_OAI21X1_348 gnd vdd FILL
XFILL_0_OAI21X1_359 gnd vdd FILL
XFILL_1_OAI21X1_519 gnd vdd FILL
XFILL_1_OAI21X1_9 gnd vdd FILL
XFILL_0_NAND2X1_310 gnd vdd FILL
XFILL_0_OAI21X1_1114 gnd vdd FILL
XFILL_0_NAND2X1_343 gnd vdd FILL
XFILL_0_OAI21X1_1103 gnd vdd FILL
XFILL_0_NAND2X1_332 gnd vdd FILL
XFILL_1_NAND2X1_514 gnd vdd FILL
XFILL_0_NAND2X1_321 gnd vdd FILL
XFILL_0_DFFPOSX1_715 gnd vdd FILL
XFILL_0_DFFPOSX1_704 gnd vdd FILL
XFILL_0_OAI21X1_1125 gnd vdd FILL
XFILL_0_OAI21X1_1147 gnd vdd FILL
XFILL_0_NAND2X1_354 gnd vdd FILL
XFILL_0_NAND2X1_376 gnd vdd FILL
XFILL_1_NAND2X1_558 gnd vdd FILL
XFILL_1_NOR2X1_1 gnd vdd FILL
XFILL_0_NAND2X1_365 gnd vdd FILL
XFILL_1_NAND2X1_547 gnd vdd FILL
XFILL_0_OAI21X1_1136 gnd vdd FILL
XFILL_0_DFFPOSX1_737 gnd vdd FILL
XFILL_0_DFFPOSX1_748 gnd vdd FILL
XFILL_0_OAI21X1_1169 gnd vdd FILL
XFILL_0_OAI21X1_1158 gnd vdd FILL
XFILL_0_DFFPOSX1_726 gnd vdd FILL
XFILL_0_NAND2X1_398 gnd vdd FILL
XFILL_0_NAND2X1_387 gnd vdd FILL
XFILL_1_NAND2X1_569 gnd vdd FILL
XFILL_0_DFFPOSX1_759 gnd vdd FILL
XFILL_5_DFFPOSX1_330 gnd vdd FILL
XFILL_5_DFFPOSX1_341 gnd vdd FILL
XFILL_5_DFFPOSX1_352 gnd vdd FILL
XFILL_5_DFFPOSX1_363 gnd vdd FILL
XFILL_5_DFFPOSX1_374 gnd vdd FILL
XFILL_24_14_0 gnd vdd FILL
XFILL_5_DFFPOSX1_396 gnd vdd FILL
XFILL_5_DFFPOSX1_385 gnd vdd FILL
XFILL_1_NAND2X1_23 gnd vdd FILL
XFILL_1_NAND2X1_12 gnd vdd FILL
XFILL_1_NAND2X1_34 gnd vdd FILL
XFILL_1_NAND2X1_56 gnd vdd FILL
XINVX4_24 bundleStartMajId_i[10] gnd INVX4_24/Y vdd INVX4
XINVX4_13 bundleStartMajId_i[35] gnd INVX4_13/Y vdd INVX4
XINVX4_35 bundleAddress_i[44] gnd INVX4_35/Y vdd INVX4
XINVX4_46 bundleAddress_i[0] gnd INVX4_46/Y vdd INVX4
XFILL_1_NAND2X1_89 gnd vdd FILL
XFILL_1_NAND2X1_78 gnd vdd FILL
XFILL_0_OAI21X1_882 gnd vdd FILL
XFILL_0_OAI21X1_860 gnd vdd FILL
XFILL_0_OAI21X1_871 gnd vdd FILL
XFILL_0_OAI21X1_893 gnd vdd FILL
XFILL_2_DFFPOSX1_30 gnd vdd FILL
XBUFX2_929 BUFX2_929/A gnd tid3_o[33] vdd BUFX2
XBUFX2_918 BUFX2_918/A gnd tid3_o[43] vdd BUFX2
XFILL_2_DFFPOSX1_52 gnd vdd FILL
XFILL_2_DFFPOSX1_63 gnd vdd FILL
XFILL_2_DFFPOSX1_809 gnd vdd FILL
XBUFX2_907 BUFX2_907/A gnd tid3_o[53] vdd BUFX2
XFILL_2_DFFPOSX1_41 gnd vdd FILL
XFILL_2_DFFPOSX1_85 gnd vdd FILL
XFILL_2_DFFPOSX1_96 gnd vdd FILL
XFILL_2_DFFPOSX1_74 gnd vdd FILL
XFILL_29_13_0 gnd vdd FILL
XFILL_0_OAI21X1_1670 gnd vdd FILL
XFILL_0_OAI21X1_1692 gnd vdd FILL
XFILL_0_OAI21X1_1681 gnd vdd FILL
XFILL_0_BUFX4_1 gnd vdd FILL
XFILL_0_BUFX2_614 gnd vdd FILL
XFILL_0_BUFX2_603 gnd vdd FILL
XFILL_0_BUFX2_658 gnd vdd FILL
XFILL_0_BUFX2_636 gnd vdd FILL
XFILL_0_BUFX2_625 gnd vdd FILL
XFILL_0_BUFX2_647 gnd vdd FILL
XFILL_4_DFFPOSX1_1020 gnd vdd FILL
XFILL_0_BUFX2_669 gnd vdd FILL
XFILL_4_DFFPOSX1_1031 gnd vdd FILL
XBUFX4_211 BUFX4_24/Y gnd BUFX4_211/Y vdd BUFX4
XBUFX4_200 BUFX4_25/Y gnd BUFX4_200/Y vdd BUFX4
XFILL_2_OAI21X1_1742 gnd vdd FILL
XBUFX4_255 INVX8_5/Y gnd BUFX4_4/A vdd BUFX4
XFILL_0_INVX2_110 gnd vdd FILL
XBUFX4_244 INVX8_1/Y gnd BUFX4_244/Y vdd BUFX4
XBUFX4_222 BUFX4_20/Y gnd BUFX4_222/Y vdd BUFX4
XBUFX4_233 BUFX4_22/Y gnd BUFX4_233/Y vdd BUFX4
XFILL_4_14_0 gnd vdd FILL
XFILL_0_INVX2_143 gnd vdd FILL
XFILL_0_INVX2_132 gnd vdd FILL
XBUFX4_266 enable_i gnd INVX8_4/A vdd BUFX4
XBUFX4_288 INVX8_2/Y gnd BUFX4_288/Y vdd BUFX4
XFILL_0_INVX2_121 gnd vdd FILL
XBUFX4_277 INVX8_7/Y gnd BUFX4_73/A vdd BUFX4
XFILL_0_INVX2_165 gnd vdd FILL
XFILL_0_INVX2_176 gnd vdd FILL
XFILL_2_OAI21X1_1797 gnd vdd FILL
XBUFX4_299 BUFX4_303/A gnd BUFX4_299/Y vdd BUFX4
XFILL_0_INVX4_1 gnd vdd FILL
XFILL_0_INVX2_154 gnd vdd FILL
XFILL_33_3_1 gnd vdd FILL
XFILL_0_INVX2_187 gnd vdd FILL
XFILL_0_INVX2_198 gnd vdd FILL
XFILL_18_2 gnd vdd FILL
XOAI21X1_1112 NAND2X1_476/Y INVX2_59/Y INVX2_60/Y gnd OAI21X1_1113/C vdd OAI21X1
XOAI21X1_1101 INVX2_55/Y BUFX4_230/Y NAND2X1_467/Y gnd OAI21X1_1101/Y vdd OAI21X1
XDFFPOSX1_713 BUFX2_358/A CLKBUF1_17/Y OAI21X1_975/Y gnd vdd DFFPOSX1
XOAI21X1_1123 INVX2_95/Y INVX4_33/Y INVX2_64/Y gnd NAND2X1_488/B vdd OAI21X1
XOAI21X1_1156 AOI21X1_38/Y OAI21X1_1156/B NAND2X1_532/Y gnd OAI21X1_1156/Y vdd OAI21X1
XOAI21X1_1145 INVX1_190/Y bundleAddress_i[37] BUFX4_238/Y gnd OAI21X1_1146/A vdd OAI21X1
XFILL_1_DFFPOSX1_900 gnd vdd FILL
XFILL_1_OAI21X1_1332 gnd vdd FILL
XDFFPOSX1_702 BUFX2_340/A CLKBUF1_40/Y OAI21X1_953/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1310 gnd vdd FILL
XFILL_1_OAI21X1_1321 gnd vdd FILL
XOAI21X1_1134 XNOR2X1_60/Y BUFX4_186/Y NAND2X1_504/Y gnd OAI21X1_1134/Y vdd OAI21X1
XFILL_0_OAI21X1_101 gnd vdd FILL
XDFFPOSX1_746 BUFX2_13/A CLKBUF1_12/Y OAI21X1_1038/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_112 gnd vdd FILL
XDFFPOSX1_757 BUFX2_6/A CLKBUF1_70/Y OAI21X1_1049/Y gnd vdd DFFPOSX1
XOAI21X1_1178 AOI21X1_40/Y OAI21X1_1178/B NAND2X1_560/Y gnd OAI21X1_1178/Y vdd OAI21X1
XDFFPOSX1_735 BUFX2_373/A CLKBUF1_73/Y OAI21X1_1019/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1343 gnd vdd FILL
XFILL_1_DFFPOSX1_922 gnd vdd FILL
XFILL_1_DFFPOSX1_933 gnd vdd FILL
XFILL_1_OAI21X1_1354 gnd vdd FILL
XFILL_1_OAI21X1_1365 gnd vdd FILL
XDFFPOSX1_724 BUFX2_361/A CLKBUF1_58/Y OAI21X1_997/Y gnd vdd DFFPOSX1
XOAI21X1_1167 XNOR2X1_71/Y BUFX4_226/Y NAND2X1_548/Y gnd OAI21X1_1167/Y vdd OAI21X1
XFILL_1_DFFPOSX1_911 gnd vdd FILL
XOAI21X1_1189 NAND2X1_575/Y NOR3X1_14/Y NAND2X1_576/Y gnd OAI21X1_1189/Y vdd OAI21X1
XFILL_1_OAI21X1_1398 gnd vdd FILL
XFILL_1_DFFPOSX1_944 gnd vdd FILL
XFILL_1_DFFPOSX1_966 gnd vdd FILL
XFILL_0_OAI21X1_123 gnd vdd FILL
XFILL_0_OAI21X1_134 gnd vdd FILL
XFILL_1_OAI21X1_1387 gnd vdd FILL
XFILL_0_OAI21X1_145 gnd vdd FILL
XFILL_1_DFFPOSX1_955 gnd vdd FILL
XFILL_1_OAI21X1_1376 gnd vdd FILL
XDFFPOSX1_779 BUFX2_30/A CLKBUF1_62/Y OAI21X1_1071/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_316 gnd vdd FILL
XFILL_1_OAI21X1_305 gnd vdd FILL
XDFFPOSX1_768 BUFX2_18/A CLKBUF1_83/Y OAI21X1_1060/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_178 gnd vdd FILL
XFILL_0_OAI21X1_167 gnd vdd FILL
XFILL_1_DFFPOSX1_999 gnd vdd FILL
XFILL_1_DFFPOSX1_977 gnd vdd FILL
XFILL_1_DFFPOSX1_988 gnd vdd FILL
XFILL_1_OAI21X1_349 gnd vdd FILL
XFILL_0_OAI21X1_156 gnd vdd FILL
XFILL_1_OAI21X1_338 gnd vdd FILL
XFILL_1_OAI21X1_327 gnd vdd FILL
XFILL_9_13_0 gnd vdd FILL
XFILL_6_DFFPOSX1_570 gnd vdd FILL
XFILL_0_OAI21X1_189 gnd vdd FILL
XFILL_6_DFFPOSX1_581 gnd vdd FILL
XFILL_6_DFFPOSX1_592 gnd vdd FILL
XFILL_0_BUFX4_11 gnd vdd FILL
XFILL_13_11_1 gnd vdd FILL
XFILL_0_BUFX4_44 gnd vdd FILL
XFILL_0_BUFX4_22 gnd vdd FILL
XFILL_0_BUFX4_33 gnd vdd FILL
XFILL_0_BUFX4_55 gnd vdd FILL
XFILL_0_BUFX4_77 gnd vdd FILL
XFILL_0_NAND2X1_140 gnd vdd FILL
XFILL_0_BUFX4_66 gnd vdd FILL
XFILL_0_NAND2X1_151 gnd vdd FILL
XFILL_1_NAND2X1_311 gnd vdd FILL
XFILL_1_BUFX4_108 gnd vdd FILL
XFILL_24_3_1 gnd vdd FILL
XFILL_1_NAND2X1_333 gnd vdd FILL
XFILL_0_DFFPOSX1_512 gnd vdd FILL
XFILL_1_BUFX4_119 gnd vdd FILL
XFILL_0_BUFX4_99 gnd vdd FILL
XFILL_0_BUFX4_88 gnd vdd FILL
XFILL_0_DFFPOSX1_501 gnd vdd FILL
XFILL_0_DFFPOSX1_523 gnd vdd FILL
XFILL_0_NAND2X1_195 gnd vdd FILL
XFILL_1_NAND2X1_366 gnd vdd FILL
XFILL_0_NAND2X1_184 gnd vdd FILL
XFILL_0_NAND2X1_162 gnd vdd FILL
XFILL_0_NAND2X1_173 gnd vdd FILL
XFILL_1_NAND2X1_377 gnd vdd FILL
XFILL_0_DFFPOSX1_545 gnd vdd FILL
XFILL_0_DFFPOSX1_534 gnd vdd FILL
XFILL_0_DFFPOSX1_567 gnd vdd FILL
XFILL_1_NAND2X1_399 gnd vdd FILL
XFILL_0_DFFPOSX1_556 gnd vdd FILL
XFILL_0_DFFPOSX1_578 gnd vdd FILL
XFILL_0_DFFPOSX1_589 gnd vdd FILL
XFILL_5_DFFPOSX1_171 gnd vdd FILL
XFILL_5_DFFPOSX1_160 gnd vdd FILL
XFILL_5_DFFPOSX1_182 gnd vdd FILL
XFILL_5_DFFPOSX1_193 gnd vdd FILL
XOAI21X1_1690 BUFX4_248/Y BUFX4_361/Y BUFX2_728/A gnd OAI21X1_1691/C vdd OAI21X1
XFILL_0_OR2X2_14 gnd vdd FILL
XFILL_1_OAI21X1_861 gnd vdd FILL
XNAND3X1_11 NOR2X1_51/Y INVX2_45/Y INVX1_21/Y gnd NOR3X1_4/A vdd NAND3X1
XFILL_18_10_1 gnd vdd FILL
XNAND3X1_22 NOR2X1_82/Y INVX1_31/Y AND2X2_13/Y gnd NOR2X1_87/B vdd NAND3X1
XFILL_1_OAI21X1_850 gnd vdd FILL
XFILL_1_OAI21X1_872 gnd vdd FILL
XFILL_7_4_1 gnd vdd FILL
XFILL_0_OAI21X1_690 gnd vdd FILL
XFILL_1_OAI21X1_883 gnd vdd FILL
XNAND3X1_55 INVX2_99/A AND2X2_29/B AND2X2_29/A gnd AND2X2_30/A vdd NAND3X1
XNAND3X1_33 INVX2_45/Y NOR2X1_51/Y NOR3X1_9/Y gnd NAND3X1_33/Y vdd NAND3X1
XNAND3X1_66 INVX1_224/Y INVX4_51/A AND2X2_23/B gnd NOR2X1_226/B vdd NAND3X1
XNAND3X1_44 INVX2_101/Y NOR2X1_159/Y INVX2_100/A gnd INVX1_224/A vdd NAND3X1
XFILL_1_OAI21X1_894 gnd vdd FILL
XFILL_31_12_1 gnd vdd FILL
XNOR2X1_11 NOR2X1_5/B NOR2X1_11/B gnd NOR2X1_11/Y vdd NOR2X1
XFILL_2_OAI21X1_1016 gnd vdd FILL
XFILL_2_OAI21X1_1027 gnd vdd FILL
XFILL_2_DFFPOSX1_639 gnd vdd FILL
XFILL_3_DFFPOSX1_20 gnd vdd FILL
XFILL_3_DFFPOSX1_53 gnd vdd FILL
XBUFX2_726 BUFX2_726/A gnd pid3_o[11] vdd BUFX2
XBUFX2_715 BUFX2_715/A gnd pid3_o[21] vdd BUFX2
XFILL_2_DFFPOSX1_606 gnd vdd FILL
XNOR2X1_44 NOR2X1_44/A NOR3X1_4/C gnd NOR2X1_45/B vdd NOR2X1
XNOR2X1_55 INVX2_37/Y NOR2X1_99/B gnd INVX1_44/A vdd NOR2X1
XNOR2X1_33 NOR3X1_6/B NOR2X1_33/B gnd NOR2X1_33/Y vdd NOR2X1
XFILL_2_DFFPOSX1_617 gnd vdd FILL
XNOR2X1_22 OR2X2_4/Y NOR2X1_22/B gnd NOR2X1_22/Y vdd NOR2X1
XBUFX2_737 BUFX2_737/A gnd pid3_o[1] vdd BUFX2
XFILL_2_DFFPOSX1_628 gnd vdd FILL
XFILL_3_DFFPOSX1_31 gnd vdd FILL
XBUFX2_704 BUFX2_704/A gnd pid2_o[28] vdd BUFX2
XFILL_3_DFFPOSX1_42 gnd vdd FILL
XFILL_3_DFFPOSX1_75 gnd vdd FILL
XBUFX2_759 BUFX2_759/A gnd pid4_o[10] vdd BUFX2
XBUFX2_748 BUFX2_748/A gnd pid4_o[20] vdd BUFX2
XFILL_3_DFFPOSX1_64 gnd vdd FILL
XFILL_3_DFFPOSX1_86 gnd vdd FILL
XNOR2X1_77 OR2X2_8/A NOR2X1_77/B gnd INVX2_48/A vdd NOR2X1
XNOR2X1_88 bundleStartMajId_i[18] INVX2_50/A gnd NOR2X1_88/Y vdd NOR2X1
XNOR2X1_66 NOR2X1_66/A MUX2X1_1/Y gnd NOR2X1_66/Y vdd NOR2X1
XNOR2X1_99 INVX2_38/Y NOR2X1_99/B gnd NOR2X1_99/Y vdd NOR2X1
XFILL_3_DFFPOSX1_97 gnd vdd FILL
XFILL_15_3_1 gnd vdd FILL
XINVX2_200 bundleTid_i[9] gnd INVX2_200/Y vdd INVX2
XFILL_0_BUFX2_411 gnd vdd FILL
XFILL_0_BUFX2_422 gnd vdd FILL
XFILL_0_BUFX2_400 gnd vdd FILL
XFILL_1_DFFPOSX1_218 gnd vdd FILL
XFILL_1_DFFPOSX1_207 gnd vdd FILL
XFILL_1_DFFPOSX1_229 gnd vdd FILL
XFILL_0_BUFX2_433 gnd vdd FILL
XFILL_0_BUFX2_466 gnd vdd FILL
XFILL_0_BUFX2_444 gnd vdd FILL
XFILL_0_BUFX2_455 gnd vdd FILL
XFILL_0_BUFX2_488 gnd vdd FILL
XFILL_0_BUFX2_499 gnd vdd FILL
XFILL_0_BUFX2_477 gnd vdd FILL
XFILL_36_11_1 gnd vdd FILL
XFILL_0_NAND2X1_20 gnd vdd FILL
XFILL_0_NAND2X1_31 gnd vdd FILL
XFILL_0_NAND2X1_64 gnd vdd FILL
XFILL_0_NAND2X1_53 gnd vdd FILL
XFILL_0_NAND2X1_42 gnd vdd FILL
XNOR2X1_123 NOR2X1_215/B INVX1_184/A gnd NOR2X1_123/Y vdd NOR2X1
XNOR2X1_101 BUFX2_581/A NOR2X1_96/B gnd NOR2X1_101/Y vdd NOR2X1
XNOR2X1_112 NOR3X1_6/B NOR2X1_112/B gnd AND2X2_21/A vdd NOR2X1
XFILL_2_OAI21X1_1594 gnd vdd FILL
XFILL_30_1 gnd vdd FILL
XNOR2X1_134 NOR2X1_220/A INVX1_186/A gnd INVX1_188/A vdd NOR2X1
XNOR2X1_145 NOR2X1_145/A INVX1_190/A gnd NOR2X1_146/B vdd NOR2X1
XFILL_0_NAND2X1_97 gnd vdd FILL
XNOR2X1_167 bundleAddress_i[13] AND2X2_24/Y gnd NOR2X1_167/Y vdd NOR2X1
XFILL_0_NAND2X1_75 gnd vdd FILL
XNOR2X1_156 INVX2_100/Y NOR2X1_160/B gnd NOR2X1_156/Y vdd NOR2X1
XFILL_0_NAND2X1_86 gnd vdd FILL
XNOR2X1_178 bundleAddress_i[56] INVX4_47/A gnd NOR2X1_178/Y vdd NOR2X1
XNOR2X1_189 NOR2X1_189/A MUX2X1_2/Y gnd NOR2X1_189/Y vdd NOR2X1
XOAI21X1_629 BUFX4_93/Y BUFX4_323/Y BUFX2_568/A gnd OAI21X1_630/C vdd OAI21X1
XOAI21X1_607 BUFX4_9/A BUFX4_325/Y BUFX2_558/A gnd OAI21X1_608/C vdd OAI21X1
XOAI21X1_618 BUFX4_112/Y BUFX4_372/Y BUFX2_562/A gnd OAI21X1_620/C vdd OAI21X1
XDFFPOSX1_510 BUFX2_540/A CLKBUF1_50/Y OAI21X1_571/Y gnd vdd DFFPOSX1
XDFFPOSX1_521 BUFX2_552/A CLKBUF1_79/Y OAI21X1_600/Y gnd vdd DFFPOSX1
XDFFPOSX1_532 NOR2X1_89/A CLKBUF1_79/Y AOI21X1_18/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1140 gnd vdd FILL
XFILL_1_DFFPOSX1_741 gnd vdd FILL
XDFFPOSX1_543 BUFX2_576/A CLKBUF1_11/Y OAI21X1_649/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1151 gnd vdd FILL
XFILL_1_OAI21X1_1173 gnd vdd FILL
XDFFPOSX1_565 BUFX2_594/A CLKBUF1_88/Y OAI21X1_708/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1184 gnd vdd FILL
XFILL_1_DFFPOSX1_730 gnd vdd FILL
XFILL_1_OAI21X1_1162 gnd vdd FILL
XDFFPOSX1_554 BUFX2_641/A CLKBUF1_94/Y OAI21X1_678/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_752 gnd vdd FILL
XFILL_1_OAI21X1_102 gnd vdd FILL
XFILL_1_DFFPOSX1_774 gnd vdd FILL
XFILL_1_OAI21X1_124 gnd vdd FILL
XFILL_1_OAI21X1_113 gnd vdd FILL
XFILL_1_OAI21X1_135 gnd vdd FILL
XDFFPOSX1_598 BUFX2_631/A CLKBUF1_100/Y OAI21X1_805/Y gnd vdd DFFPOSX1
XDFFPOSX1_587 BUFX2_618/A CLKBUF1_9/Y OAI21X1_769/Y gnd vdd DFFPOSX1
XNAND2X1_602 bundleAddress_i[40] bundleAddress_i[39] gnd OR2X2_19/A vdd NAND2X1
XFILL_1_DFFPOSX1_763 gnd vdd FILL
XDFFPOSX1_576 BUFX2_606/A CLKBUF1_88/Y OAI21X1_741/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1195 gnd vdd FILL
XFILL_1_DFFPOSX1_785 gnd vdd FILL
XFILL_1_OAI21X1_168 gnd vdd FILL
XFILL_1_OAI21X1_146 gnd vdd FILL
XNAND2X1_624 INVX2_94/A INVX4_50/A gnd NOR2X1_220/B vdd NAND2X1
XNAND2X1_635 INVX4_51/A AND2X2_23/B gnd INVX1_223/A vdd NAND2X1
XNAND2X1_646 NAND2X1_646/A INVX2_112/A gnd NAND2X1_646/Y vdd NAND2X1
XNAND2X1_613 bundleAddress_i[22] bundleAddress_i[21] gnd NOR2X1_201/B vdd NAND2X1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XFILL_1_OAI21X1_157 gnd vdd FILL
XFILL_1_DFFPOSX1_796 gnd vdd FILL
XNAND2X1_657 BUFX2_678/A BUFX4_336/Y gnd NAND2X1_657/Y vdd NAND2X1
XFILL_1_OAI21X1_179 gnd vdd FILL
XNAND2X1_668 BUFX2_659/A BUFX4_366/Y gnd NAND2X1_668/Y vdd NAND2X1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XNAND2X1_679 BUFX2_671/A NAND2X1_7/B gnd NAND2X1_679/Y vdd NAND2X1
XINVX1_58 INVX1_58/A gnd INVX1_58/Y vdd INVX1
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XINVX1_69 INVX1_69/A gnd INVX1_69/Y vdd INVX1
XFILL_1_NAND2X1_130 gnd vdd FILL
XFILL_0_DFFPOSX1_342 gnd vdd FILL
XFILL_0_DFFPOSX1_331 gnd vdd FILL
XFILL_1_NAND2X1_174 gnd vdd FILL
XFILL_1_NAND2X1_163 gnd vdd FILL
XFILL_0_DFFPOSX1_320 gnd vdd FILL
XFILL_0_DFFPOSX1_353 gnd vdd FILL
XFILL_0_DFFPOSX1_375 gnd vdd FILL
XFILL_0_DFFPOSX1_364 gnd vdd FILL
XFILL_1_NAND2X1_185 gnd vdd FILL
XFILL_1_NAND2X1_196 gnd vdd FILL
XFILL_0_DFFPOSX1_397 gnd vdd FILL
XFILL_0_DFFPOSX1_386 gnd vdd FILL
XFILL_3_DFFPOSX1_813 gnd vdd FILL
XFILL_3_DFFPOSX1_802 gnd vdd FILL
XFILL_3_DFFPOSX1_835 gnd vdd FILL
XFILL_3_DFFPOSX1_824 gnd vdd FILL
XFILL_3_DFFPOSX1_857 gnd vdd FILL
XFILL_3_DFFPOSX1_846 gnd vdd FILL
XFILL_3_DFFPOSX1_879 gnd vdd FILL
XFILL_3_DFFPOSX1_868 gnd vdd FILL
XFILL_1_NOR2X1_230 gnd vdd FILL
XFILL_1_OAI21X1_680 gnd vdd FILL
XFILL_1_OAI21X1_691 gnd vdd FILL
XFILL_2_DFFPOSX1_414 gnd vdd FILL
XFILL_1_INVX1_185 gnd vdd FILL
XBUFX2_512 BUFX2_512/A gnd majID2_o[4] vdd BUFX2
XBUFX2_501 BUFX2_501/A gnd majID2_o[14] vdd BUFX2
XFILL_2_DFFPOSX1_403 gnd vdd FILL
XFILL_4_DFFPOSX1_21 gnd vdd FILL
XFILL_4_DFFPOSX1_32 gnd vdd FILL
XBUFX2_545 BUFX2_545/A gnd majID3_o[33] vdd BUFX2
XBUFX2_534 BUFX2_534/A gnd majID3_o[43] vdd BUFX2
XBUFX2_523 BUFX2_523/A gnd majID3_o[53] vdd BUFX2
XFILL_2_DFFPOSX1_447 gnd vdd FILL
XFILL_4_DFFPOSX1_10 gnd vdd FILL
XFILL_2_DFFPOSX1_425 gnd vdd FILL
XFILL_2_DFFPOSX1_436 gnd vdd FILL
XBUFX2_578 BUFX2_578/A gnd majID3_o[3] vdd BUFX2
XFILL_4_DFFPOSX1_43 gnd vdd FILL
XBUFX2_567 BUFX2_567/A gnd majID3_o[13] vdd BUFX2
XFILL_2_DFFPOSX1_458 gnd vdd FILL
XFILL_2_DFFPOSX1_469 gnd vdd FILL
XFILL_4_DFFPOSX1_54 gnd vdd FILL
XFILL_4_DFFPOSX1_65 gnd vdd FILL
XBUFX2_556 NOR2X1_81/A gnd majID3_o[23] vdd BUFX2
XFILL_4_DFFPOSX1_76 gnd vdd FILL
XFILL_4_DFFPOSX1_87 gnd vdd FILL
XBUFX2_589 BUFX2_589/A gnd majID4_o[51] vdd BUFX2
XFILL_4_DFFPOSX1_98 gnd vdd FILL
XFILL_5_DFFPOSX1_918 gnd vdd FILL
XFILL_5_DFFPOSX1_929 gnd vdd FILL
XFILL_5_DFFPOSX1_907 gnd vdd FILL
XFILL_30_1_1 gnd vdd FILL
XFILL_22_17_1 gnd vdd FILL
XFILL_0_BUFX2_230 gnd vdd FILL
XFILL_0_BUFX2_241 gnd vdd FILL
XFILL_0_BUFX2_274 gnd vdd FILL
XFILL_0_BUFX2_252 gnd vdd FILL
XFILL_0_BUFX2_263 gnd vdd FILL
XFILL_0_BUFX2_285 gnd vdd FILL
XFILL_0_BUFX2_296 gnd vdd FILL
XFILL_0_AND2X2_9 gnd vdd FILL
XFILL_4_DFFPOSX1_519 gnd vdd FILL
XFILL_4_DFFPOSX1_508 gnd vdd FILL
XFILL_38_2_1 gnd vdd FILL
XFILL_2_DFFPOSX1_981 gnd vdd FILL
XFILL_2_DFFPOSX1_970 gnd vdd FILL
XFILL_2_DFFPOSX1_992 gnd vdd FILL
XFILL_1_BUFX2_409 gnd vdd FILL
XFILL_27_16_1 gnd vdd FILL
XFILL_21_1_1 gnd vdd FILL
XFILL_0_NAND3X1_4 gnd vdd FILL
XOAI21X1_404 OAI21X1_404/A BUFX4_222/Y OAI21X1_404/C gnd OAI21X1_404/Y vdd OAI21X1
XFILL_3_DFFPOSX1_109 gnd vdd FILL
XOAI21X1_437 XNOR2X1_10/Y BUFX4_209/Y OAI21X1_437/C gnd OAI21X1_437/Y vdd OAI21X1
XOAI21X1_426 INVX1_10/A INVX4_7/Y INVX2_18/Y gnd OAI21X1_426/Y vdd OAI21X1
XOAI21X1_415 OAI21X1_415/A BUFX4_181/Y OAI21X1_415/C gnd OAI21X1_415/Y vdd OAI21X1
XOAI21X1_448 INVX1_16/A bundleStartMajId_i[31] BUFX4_245/Y gnd OAI21X1_449/B vdd OAI21X1
XOAI21X1_459 OAI21X1_459/A NOR2X1_35/Y OAI21X1_459/C gnd OAI21X1_459/Y vdd OAI21X1
XFILL_21_12_0 gnd vdd FILL
XFILL_3_XNOR2X1_50 gnd vdd FILL
XDFFPOSX1_340 BUFX2_1012/A CLKBUF1_3/Y OAI21X1_297/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_72 gnd vdd FILL
XFILL_3_XNOR2X1_83 gnd vdd FILL
XFILL_3_XNOR2X1_61 gnd vdd FILL
XFILL_1_DFFPOSX1_560 gnd vdd FILL
XDFFPOSX1_373 BUFX2_402/A CLKBUF1_48/Y OAI21X1_345/Y gnd vdd DFFPOSX1
XDFFPOSX1_362 BUFX2_449/A CLKBUF1_66/Y OAI21X1_334/Y gnd vdd DFFPOSX1
XDFFPOSX1_351 BUFX2_1024/A CLKBUF1_77/Y OAI21X1_319/Y gnd vdd DFFPOSX1
XFILL_2_OAI21X1_103 gnd vdd FILL
XNAND2X1_410 BUFX2_63/A BUFX4_382/Y gnd NAND2X1_410/Y vdd NAND2X1
XDFFPOSX1_395 BUFX2_426/A CLKBUF1_5/Y OAI21X1_367/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_582 gnd vdd FILL
XFILL_1_DFFPOSX1_593 gnd vdd FILL
XDFFPOSX1_384 BUFX2_414/A CLKBUF1_15/Y OAI21X1_356/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_571 gnd vdd FILL
XNAND2X1_432 BUFX2_25/A BUFX4_377/Y gnd NAND2X1_432/Y vdd NAND2X1
XNAND2X1_421 BUFX2_12/A OAI21X1_5/A gnd NAND2X1_421/Y vdd NAND2X1
XNAND2X1_443 BUFX2_37/A BUFX4_384/Y gnd NAND2X1_443/Y vdd NAND2X1
XFILL_2_OAI21X1_136 gnd vdd FILL
XNAND2X1_454 BUFX2_49/A BUFX4_364/Y gnd NAND2X1_454/Y vdd NAND2X1
XNAND2X1_487 bundleAddress_i[52] bundleAddress_i[51] gnd INVX2_96/A vdd NAND2X1
XNAND2X1_476 INVX1_185/Y INVX1_184/A gnd NAND2X1_476/Y vdd NAND2X1
XNAND2X1_465 BUFX2_61/A BUFX4_360/Y gnd NAND2X1_465/Y vdd NAND2X1
XFILL_29_2_1 gnd vdd FILL
XNAND2X1_498 BUFX2_73/A BUFX4_223/Y gnd NAND2X1_498/Y vdd NAND2X1
XFILL_4_2_1 gnd vdd FILL
XFILL_0_INVX1_219 gnd vdd FILL
XFILL_0_INVX1_208 gnd vdd FILL
XFILL_2_17_1 gnd vdd FILL
XFILL_1_XNOR2X1_100 gnd vdd FILL
XFILL_0_DFFPOSX1_150 gnd vdd FILL
XFILL_1_BUFX2_921 gnd vdd FILL
XFILL_0_DFFPOSX1_183 gnd vdd FILL
XFILL_26_11_0 gnd vdd FILL
XFILL_0_DFFPOSX1_161 gnd vdd FILL
XFILL_12_1_1 gnd vdd FILL
XFILL_0_DFFPOSX1_172 gnd vdd FILL
XFILL_1_BUFX2_910 gnd vdd FILL
XFILL_0_DFFPOSX1_194 gnd vdd FILL
XFILL_1_BUFX2_954 gnd vdd FILL
XFILL_0_OAI21X1_29 gnd vdd FILL
XFILL_1_BUFX2_965 gnd vdd FILL
XFILL_0_OAI21X1_18 gnd vdd FILL
XFILL_3_DFFPOSX1_632 gnd vdd FILL
XFILL_3_DFFPOSX1_621 gnd vdd FILL
XFILL_3_DFFPOSX1_610 gnd vdd FILL
XFILL_1_BUFX2_998 gnd vdd FILL
XOAI21X1_960 BUFX4_7/A BUFX4_315/Y BUFX2_344/A gnd OAI21X1_961/C vdd OAI21X1
XFILL_3_DFFPOSX1_654 gnd vdd FILL
XOAI21X1_971 BUFX4_178/Y INVX1_140/Y OAI21X1_971/C gnd OAI21X1_971/Y vdd OAI21X1
XOAI21X1_993 BUFX4_296/Y INVX1_151/Y OAI21X1_993/C gnd OAI21X1_993/Y vdd OAI21X1
XFILL_3_DFFPOSX1_643 gnd vdd FILL
XFILL_3_DFFPOSX1_665 gnd vdd FILL
XOAI21X1_982 BUFX4_152/Y BUFX4_35/Y BUFX2_384/A gnd OAI21X1_983/C vdd OAI21X1
XFILL_3_DFFPOSX1_698 gnd vdd FILL
XFILL_3_DFFPOSX1_687 gnd vdd FILL
XFILL_3_DFFPOSX1_676 gnd vdd FILL
XINVX2_90 bundleAddress_i[4] gnd INVX2_90/Y vdd INVX2
XFILL_7_16_1 gnd vdd FILL
XFILL_2_DFFPOSX1_211 gnd vdd FILL
XFILL_2_DFFPOSX1_200 gnd vdd FILL
XBUFX2_320 BUFX2_320/A gnd instr2_o[26] vdd BUFX2
XFILL_2_DFFPOSX1_222 gnd vdd FILL
XFILL_0_NAND2X1_717 gnd vdd FILL
XFILL_0_NAND2X1_706 gnd vdd FILL
XFILL_5_DFFPOSX1_11 gnd vdd FILL
XBUFX2_342 BUFX2_342/A gnd instr3_o[7] vdd BUFX2
XBUFX2_331 BUFX2_331/A gnd instr3_o[17] vdd BUFX2
XFILL_2_DFFPOSX1_255 gnd vdd FILL
XFILL_0_NAND2X1_739 gnd vdd FILL
XFILL_2_DFFPOSX1_244 gnd vdd FILL
XFILL_1_12_0 gnd vdd FILL
XFILL_0_NAND2X1_728 gnd vdd FILL
XFILL_2_DFFPOSX1_233 gnd vdd FILL
XBUFX2_353 BUFX2_353/A gnd instr3_o[25] vdd BUFX2
XFILL_2_DFFPOSX1_266 gnd vdd FILL
XFILL_5_DFFPOSX1_44 gnd vdd FILL
XBUFX2_375 BUFX2_375/A gnd instr4_o[6] vdd BUFX2
XFILL_5_DFFPOSX1_22 gnd vdd FILL
XBUFX2_364 BUFX2_364/A gnd instr4_o[16] vdd BUFX2
XFILL_5_DFFPOSX1_55 gnd vdd FILL
XFILL_2_DFFPOSX1_277 gnd vdd FILL
XFILL_5_DFFPOSX1_33 gnd vdd FILL
XBUFX2_386 BUFX2_386/A gnd instr4_o[24] vdd BUFX2
XFILL_2_DFFPOSX1_288 gnd vdd FILL
XOAI21X1_20 INVX2_158/Y BUFX4_227/Y OAI21X1_20/C gnd OAI21X1_20/Y vdd OAI21X1
XFILL_32_9_0 gnd vdd FILL
XFILL_5_DFFPOSX1_77 gnd vdd FILL
XFILL_2_DFFPOSX1_299 gnd vdd FILL
XFILL_5_DFFPOSX1_88 gnd vdd FILL
XFILL_1_NOR3X1_14 gnd vdd FILL
XFILL_5_DFFPOSX1_66 gnd vdd FILL
XBUFX2_397 BUFX2_397/A gnd majID1_o[51] vdd BUFX2
XFILL_5_DFFPOSX1_715 gnd vdd FILL
XOAI21X1_53 INVX2_191/Y BUFX4_198/Y OAI21X1_53/C gnd OAI21X1_53/Y vdd OAI21X1
XFILL_5_DFFPOSX1_704 gnd vdd FILL
XOAI21X1_42 INVX2_180/Y BUFX4_234/Y OAI21X1_42/C gnd OAI21X1_42/Y vdd OAI21X1
XFILL_5_DFFPOSX1_737 gnd vdd FILL
XOAI21X1_31 INVX2_169/Y BUFX4_195/Y OAI21X1_31/C gnd OAI21X1_31/Y vdd OAI21X1
XFILL_5_DFFPOSX1_726 gnd vdd FILL
XFILL_5_DFFPOSX1_99 gnd vdd FILL
XOAI21X1_64 INVX2_202/Y BUFX4_207/Y OAI21X1_64/C gnd OAI21X1_64/Y vdd OAI21X1
XFILL_5_DFFPOSX1_759 gnd vdd FILL
XFILL_5_DFFPOSX1_748 gnd vdd FILL
XOAI21X1_75 OR2X2_20/B OAI21X1_9/A OAI21X1_75/C gnd OAI21X1_75/Y vdd OAI21X1
XFILL_1_BUFX4_291 gnd vdd FILL
XOAI21X1_86 BUFX4_1/Y BUFX4_348/Y BUFX2_966/A gnd OAI21X1_87/C vdd OAI21X1
XFILL_1_BUFX4_280 gnd vdd FILL
XOAI21X1_97 BUFX4_165/Y INVX2_158/Y OAI21X1_97/C gnd OAI21X1_97/Y vdd OAI21X1
XFILL_4_DFFPOSX1_316 gnd vdd FILL
XFILL_0_DFFPOSX1_51 gnd vdd FILL
XFILL_0_DFFPOSX1_62 gnd vdd FILL
XFILL_4_DFFPOSX1_327 gnd vdd FILL
XFILL_0_DFFPOSX1_40 gnd vdd FILL
XFILL_4_DFFPOSX1_305 gnd vdd FILL
XFILL_0_DFFPOSX1_84 gnd vdd FILL
XFILL_0_DFFPOSX1_95 gnd vdd FILL
XFILL_4_DFFPOSX1_349 gnd vdd FILL
XFILL_4_DFFPOSX1_338 gnd vdd FILL
XFILL_0_DFFPOSX1_73 gnd vdd FILL
XFILL_6_11_0 gnd vdd FILL
XFILL_2_DFFPOSX1_1019 gnd vdd FILL
XFILL_2_DFFPOSX1_1008 gnd vdd FILL
XFILL_23_9_0 gnd vdd FILL
XFILL_1_BUFX2_206 gnd vdd FILL
XOAI21X1_201 OAI21X1_8/A BUFX4_291/Y OAI21X1_201/C gnd OAI21X1_201/Y vdd OAI21X1
XOAI21X1_212 BUFX4_174/Y BUFX4_56/Y BUFX2_1025/A gnd OAI21X1_213/C vdd OAI21X1
XFILL_1_BUFX2_239 gnd vdd FILL
XFILL_6_DFFPOSX1_3 gnd vdd FILL
XOAI21X1_234 BUFX4_150/Y BUFX4_71/Y BUFX2_978/A gnd OAI21X1_235/C vdd OAI21X1
XOAI21X1_223 INVX2_157/Y BUFX4_292/Y OAI21X1_223/C gnd OAI21X1_223/Y vdd OAI21X1
XOAI21X1_245 INVX2_168/Y BUFX4_297/Y OAI21X1_245/C gnd OAI21X1_245/Y vdd OAI21X1
XOAI21X1_256 BUFX4_158/Y BUFX4_28/Y BUFX2_990/A gnd OAI21X1_257/C vdd OAI21X1
XOAI21X1_289 INVX2_190/Y BUFX4_292/Y OAI21X1_289/C gnd OAI21X1_289/Y vdd OAI21X1
XOAI21X1_267 INVX2_179/Y BUFX4_296/Y OAI21X1_267/C gnd OAI21X1_267/Y vdd OAI21X1
XOAI21X1_278 BUFX4_140/Y BUFX4_45/Y BUFX2_1002/A gnd OAI21X1_279/C vdd OAI21X1
XAND2X2_12 bundleStartMajId_i[50] bundleStartMajId_i[49] gnd AND2X2_12/Y vdd AND2X2
XAND2X2_23 INVX1_188/A AND2X2_23/B gnd AND2X2_24/A vdd AND2X2
XDFFPOSX1_181 BUFX2_850/A CLKBUF1_74/Y OAI21X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_170 BUFX2_897/A CLKBUF1_26/Y OAI21X1_14/Y gnd vdd DFFPOSX1
XFILL_0_NOR3X1_2 gnd vdd FILL
XDFFPOSX1_192 BUFX2_862/A CLKBUF1_82/Y OAI21X1_36/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_390 gnd vdd FILL
XNAND2X1_240 BUFX2_504/A BUFX4_200/Y gnd OAI21X1_478/C vdd NAND2X1
XNAND2X1_262 INVX1_23/Y NOR2X1_52/Y gnd OAI21X1_499/A vdd NAND2X1
XNAND2X1_251 BUFX2_509/A BUFX4_221/Y gnd OAI21X1_487/C vdd NAND2X1
XFILL_4_DFFPOSX1_850 gnd vdd FILL
XNAND2X1_284 NOR2X1_19/Y NOR2X1_69/Y gnd OR2X2_6/B vdd NAND2X1
XNAND2X1_295 bundleStartMajId_i[22] bundleStartMajId_i[21] gnd INVX1_32/A vdd NAND2X1
XNAND2X1_273 AND2X2_12/Y OAI22X1_1/C gnd XNOR2X1_27/A vdd NAND2X1
XFILL_4_DFFPOSX1_883 gnd vdd FILL
XFILL_4_DFFPOSX1_872 gnd vdd FILL
XFILL_4_DFFPOSX1_861 gnd vdd FILL
XFILL_4_DFFPOSX1_894 gnd vdd FILL
XFILL_12_17_0 gnd vdd FILL
XFILL_0_OAI21X1_1 gnd vdd FILL
XFILL_14_9_0 gnd vdd FILL
XFILL_2_XNOR2X1_101 gnd vdd FILL
XFILL_1_BUFX2_762 gnd vdd FILL
XFILL_1_BUFX2_751 gnd vdd FILL
XFILL_0_BUFX4_325 gnd vdd FILL
XFILL_0_BUFX4_303 gnd vdd FILL
XFILL_1_NOR2X1_80 gnd vdd FILL
XFILL_1_NOR2X1_91 gnd vdd FILL
XFILL_1_BUFX2_773 gnd vdd FILL
XFILL_0_BUFX4_314 gnd vdd FILL
XFILL_1_BUFX2_795 gnd vdd FILL
XFILL_0_BUFX4_336 gnd vdd FILL
XFILL_0_BUFX4_347 gnd vdd FILL
XOAI21X1_1519 INVX2_111/Y NOR2X1_226/B OAI21X1_1519/C gnd OAI21X1_1521/A vdd OAI21X1
XOAI21X1_1508 BUFX4_121/Y BUFX4_66/Y BUFX2_229/A gnd OAI21X1_1509/C vdd OAI21X1
XFILL_0_BUFX4_358 gnd vdd FILL
XFILL_1_OAI21X1_1706 gnd vdd FILL
XFILL_3_DFFPOSX1_440 gnd vdd FILL
XFILL_1_OAI21X1_1739 gnd vdd FILL
XFILL_1_OAI21X1_1728 gnd vdd FILL
XFILL_1_OAI21X1_1717 gnd vdd FILL
XFILL_3_DFFPOSX1_462 gnd vdd FILL
XOAI21X1_790 BUFX4_122/Y BUFX4_69/Y BUFX2_626/A gnd OAI21X1_792/C vdd OAI21X1
XFILL_3_DFFPOSX1_451 gnd vdd FILL
XFILL_3_DFFPOSX1_473 gnd vdd FILL
XFILL_0_BUFX4_369 gnd vdd FILL
XFILL_0_BUFX2_1007 gnd vdd FILL
XFILL_3_DFFPOSX1_484 gnd vdd FILL
XFILL_3_DFFPOSX1_495 gnd vdd FILL
XFILL_0_OAI21X1_508 gnd vdd FILL
XFILL_0_OAI21X1_519 gnd vdd FILL
XFILL_0_BUFX2_1018 gnd vdd FILL
XFILL_6_DFFPOSX1_900 gnd vdd FILL
XFILL_0_BUFX2_1029 gnd vdd FILL
XFILL_6_2 gnd vdd FILL
XFILL_17_16_0 gnd vdd FILL
XFILL_6_DFFPOSX1_988 gnd vdd FILL
XFILL_6_DFFPOSX1_999 gnd vdd FILL
XFILL_0_CLKBUF1_19 gnd vdd FILL
XFILL_30_18_0 gnd vdd FILL
XFILL_0_NAND2X1_525 gnd vdd FILL
XFILL_0_NAND2X1_514 gnd vdd FILL
XFILL_0_NAND2X1_503 gnd vdd FILL
XFILL_1_NAND2X1_729 gnd vdd FILL
XFILL_35_0_1 gnd vdd FILL
XFILL_2_XNOR2X1_91 gnd vdd FILL
XBUFX2_150 BUFX2_150/A gnd addr3_o[35] vdd BUFX2
XFILL_0_NAND2X1_558 gnd vdd FILL
XFILL_2_XNOR2X1_80 gnd vdd FILL
XFILL_0_OAI21X1_1329 gnd vdd FILL
XFILL_1_NAND2X1_718 gnd vdd FILL
XFILL_0_NAND2X1_536 gnd vdd FILL
XFILL_0_OAI21X1_1307 gnd vdd FILL
XFILL_0_OAI21X1_1318 gnd vdd FILL
XFILL_0_NAND2X1_547 gnd vdd FILL
XBUFX2_161 BUFX2_161/A gnd addr3_o[25] vdd BUFX2
XFILL_0_NAND2X1_569 gnd vdd FILL
XFILL_0_DFFPOSX1_919 gnd vdd FILL
XBUFX2_172 BUFX2_172/A gnd addr3_o[15] vdd BUFX2
XBUFX2_194 BUFX2_194/A gnd addr4_o[62] vdd BUFX2
XFILL_1_NAND2X1_2 gnd vdd FILL
XBUFX2_183 BUFX2_183/A gnd addr3_o[5] vdd BUFX2
XFILL_0_DFFPOSX1_908 gnd vdd FILL
XFILL_5_DFFPOSX1_512 gnd vdd FILL
XFILL_5_DFFPOSX1_501 gnd vdd FILL
XFILL_6_DFFPOSX1_78 gnd vdd FILL
XFILL_5_DFFPOSX1_545 gnd vdd FILL
XFILL_6_DFFPOSX1_89 gnd vdd FILL
XFILL_5_DFFPOSX1_534 gnd vdd FILL
XFILL_5_DFFPOSX1_523 gnd vdd FILL
XFILL_5_DFFPOSX1_578 gnd vdd FILL
XFILL_5_DFFPOSX1_567 gnd vdd FILL
XFILL_5_DFFPOSX1_556 gnd vdd FILL
XFILL_5_DFFPOSX1_589 gnd vdd FILL
XBUFX2_1020 BUFX2_1020/A gnd tid4_o[8] vdd BUFX2
XBUFX2_1031 BUFX2_1031/A gnd tid4_o[55] vdd BUFX2
XFILL_1_AOI21X1_7 gnd vdd FILL
XFILL_35_17_0 gnd vdd FILL
XCLKBUF1_32 BUFX4_87/Y gnd CLKBUF1_32/Y vdd CLKBUF1
XCLKBUF1_21 BUFX4_92/Y gnd CLKBUF1_21/Y vdd CLKBUF1
XCLKBUF1_10 BUFX4_90/Y gnd CLKBUF1_10/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_102 gnd vdd FILL
XFILL_4_DFFPOSX1_124 gnd vdd FILL
XCLKBUF1_65 BUFX4_84/Y gnd CLKBUF1_65/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_30 gnd vdd FILL
XCLKBUF1_43 BUFX4_86/Y gnd CLKBUF1_43/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_135 gnd vdd FILL
XCLKBUF1_54 BUFX4_90/Y gnd CLKBUF1_54/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_113 gnd vdd FILL
XFILL_1_DFFPOSX1_41 gnd vdd FILL
XFILL_4_DFFPOSX1_157 gnd vdd FILL
XFILL_4_DFFPOSX1_168 gnd vdd FILL
XCLKBUF1_98 BUFX4_85/Y gnd CLKBUF1_98/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_52 gnd vdd FILL
XFILL_1_DFFPOSX1_63 gnd vdd FILL
XCLKBUF1_87 BUFX4_83/Y gnd CLKBUF1_87/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_146 gnd vdd FILL
XFILL_1_DFFPOSX1_74 gnd vdd FILL
XCLKBUF1_76 BUFX4_89/Y gnd CLKBUF1_76/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_179 gnd vdd FILL
XFILL_1_DFFPOSX1_85 gnd vdd FILL
XFILL_1_DFFPOSX1_96 gnd vdd FILL
XFILL_26_0_1 gnd vdd FILL
XFILL_2_BUFX4_267 gnd vdd FILL
XFILL_1_0_1 gnd vdd FILL
XFILL_0_OAI21X1_1830 gnd vdd FILL
XFILL_0_BUFX2_829 gnd vdd FILL
XFILL_0_BUFX2_807 gnd vdd FILL
XFILL_0_BUFX2_818 gnd vdd FILL
XINVX1_106 bundle_i[34] gnd INVX1_106/Y vdd INVX1
XINVX1_139 bundle_i[65] gnd INVX1_139/Y vdd INVX1
XINVX1_117 bundle_i[87] gnd INVX1_117/Y vdd INVX1
XINVX1_128 bundle_i[76] gnd INVX1_128/Y vdd INVX1
XFILL_3_XNOR2X1_5 gnd vdd FILL
XFILL_9_1_1 gnd vdd FILL
XFILL_0_INVX2_27 gnd vdd FILL
XFILL_0_INVX2_16 gnd vdd FILL
XFILL_0_INVX2_38 gnd vdd FILL
XFILL_0_INVX2_49 gnd vdd FILL
XFILL_4_DFFPOSX1_691 gnd vdd FILL
XFILL_4_DFFPOSX1_680 gnd vdd FILL
XFILL_17_0_1 gnd vdd FILL
XFILL_0_CLKBUF1_6 gnd vdd FILL
XFILL_4_CLKBUF1_5 gnd vdd FILL
XFILL_0_BUFX4_100 gnd vdd FILL
XFILL_1_BUFX2_570 gnd vdd FILL
XFILL_0_BUFX4_111 gnd vdd FILL
XFILL_0_BUFX4_133 gnd vdd FILL
XFILL_0_BUFX4_122 gnd vdd FILL
XOAI21X1_1305 XNOR2X1_82/Y BUFX4_152/Y OAI21X1_1305/C gnd OAI21X1_1305/Y vdd OAI21X1
XOAI21X1_1338 NOR2X1_205/Y OAI21X1_1338/B OAI21X1_1338/C gnd OAI21X1_1338/Y vdd OAI21X1
XDFFPOSX1_906 BUFX2_157/A CLKBUF1_89/Y OAI21X1_1303/Y gnd vdd DFFPOSX1
XFILL_1_BUFX2_11 gnd vdd FILL
XFILL_0_BUFX4_166 gnd vdd FILL
XOAI21X1_1327 NAND2X1_616/Y BUFX4_160/Y OAI21X1_1327/C gnd OAI21X1_1327/Y vdd OAI21X1
XFILL_0_BUFX4_155 gnd vdd FILL
XFILL_1_OAI21X1_1514 gnd vdd FILL
XFILL_0_BUFX4_144 gnd vdd FILL
XOAI21X1_1316 BUFX4_6/A BUFX4_350/Y BUFX2_164/A gnd OAI21X1_1319/C vdd OAI21X1
XFILL_1_OAI21X1_1503 gnd vdd FILL
XFILL_3_DFFPOSX1_281 gnd vdd FILL
XDFFPOSX1_939 BUFX2_216/A CLKBUF1_43/Y OAI21X1_1391/Y gnd vdd DFFPOSX1
XFILL_1_BUFX2_44 gnd vdd FILL
XFILL_1_OAI21X1_1525 gnd vdd FILL
XFILL_1_BUFX2_55 gnd vdd FILL
XFILL_1_OAI21X1_1558 gnd vdd FILL
XDFFPOSX1_917 BUFX2_169/A CLKBUF1_77/Y OAI21X1_1332/Y gnd vdd DFFPOSX1
XFILL_0_BUFX4_177 gnd vdd FILL
XFILL_0_BUFX4_188 gnd vdd FILL
XFILL_1_OAI21X1_1536 gnd vdd FILL
XOAI21X1_1349 XNOR2X1_86/Y BUFX4_144/Y OAI21X1_1349/C gnd OAI21X1_1349/Y vdd OAI21X1
XFILL_1_OAI21X1_1547 gnd vdd FILL
XFILL_3_DFFPOSX1_270 gnd vdd FILL
XFILL_0_BUFX4_199 gnd vdd FILL
XDFFPOSX1_928 BUFX2_181/A CLKBUF1_37/Y OAI21X1_1364/Y gnd vdd DFFPOSX1
XFILL_1_BUFX2_88 gnd vdd FILL
XFILL_3_DFFPOSX1_292 gnd vdd FILL
XFILL_1_OAI21X1_1569 gnd vdd FILL
XFILL_1_OAI21X1_509 gnd vdd FILL
XFILL_0_OAI21X1_327 gnd vdd FILL
XFILL_0_OAI21X1_316 gnd vdd FILL
XFILL_0_OAI21X1_305 gnd vdd FILL
XFILL_1_BUFX2_99 gnd vdd FILL
XFILL_0_OAI21X1_349 gnd vdd FILL
XFILL_0_OAI21X1_338 gnd vdd FILL
XFILL_6_DFFPOSX1_741 gnd vdd FILL
XFILL_6_DFFPOSX1_752 gnd vdd FILL
XFILL_6_DFFPOSX1_763 gnd vdd FILL
XFILL_6_DFFPOSX1_774 gnd vdd FILL
XFILL_6_DFFPOSX1_785 gnd vdd FILL
XFILL_6_DFFPOSX1_796 gnd vdd FILL
XFILL_37_8_0 gnd vdd FILL
XFILL_0_NAND2X1_300 gnd vdd FILL
XFILL_1_NAND2X1_515 gnd vdd FILL
XFILL_0_OAI21X1_1104 gnd vdd FILL
XFILL_0_NAND2X1_333 gnd vdd FILL
XFILL_0_NAND2X1_322 gnd vdd FILL
XFILL_0_NAND2X1_344 gnd vdd FILL
XFILL_1_NAND2X1_504 gnd vdd FILL
XFILL_0_NAND2X1_311 gnd vdd FILL
XFILL_0_NAND2X1_377 gnd vdd FILL
XFILL_0_OAI21X1_1126 gnd vdd FILL
XFILL_0_NAND2X1_355 gnd vdd FILL
XFILL_0_OAI21X1_1115 gnd vdd FILL
XFILL_0_DFFPOSX1_716 gnd vdd FILL
XFILL_1_NAND2X1_526 gnd vdd FILL
XFILL_0_OAI21X1_1148 gnd vdd FILL
XFILL_0_NAND2X1_366 gnd vdd FILL
XFILL_1_NAND2X1_548 gnd vdd FILL
XFILL_0_DFFPOSX1_705 gnd vdd FILL
XFILL_0_OAI21X1_1137 gnd vdd FILL
XFILL_0_DFFPOSX1_749 gnd vdd FILL
XFILL_0_DFFPOSX1_727 gnd vdd FILL
XFILL_0_NAND2X1_399 gnd vdd FILL
XFILL_0_NAND2X1_388 gnd vdd FILL
XFILL_0_OAI21X1_1159 gnd vdd FILL
XFILL_0_DFFPOSX1_738 gnd vdd FILL
XFILL_5_DFFPOSX1_320 gnd vdd FILL
XFILL_5_DFFPOSX1_342 gnd vdd FILL
XFILL_5_DFFPOSX1_353 gnd vdd FILL
XFILL_5_DFFPOSX1_331 gnd vdd FILL
XFILL_20_7_0 gnd vdd FILL
XFILL_24_14_1 gnd vdd FILL
XFILL_5_DFFPOSX1_375 gnd vdd FILL
XFILL_5_DFFPOSX1_386 gnd vdd FILL
XFILL_5_DFFPOSX1_364 gnd vdd FILL
XFILL_5_DFFPOSX1_397 gnd vdd FILL
XFILL_1_NAND2X1_13 gnd vdd FILL
XFILL_1_NAND2X1_35 gnd vdd FILL
XINVX4_25 bundleStartMajId_i[6] gnd INVX4_25/Y vdd INVX4
XFILL_1_NAND2X1_57 gnd vdd FILL
XINVX4_14 bundleStartMajId_i[34] gnd INVX4_14/Y vdd INVX4
XINVX4_36 bundleAddress_i[42] gnd OR2X2_18/B vdd INVX4
XINVX4_47 INVX4_47/A gnd INVX4_47/Y vdd INVX4
XFILL_1_NAND2X1_79 gnd vdd FILL
XFILL_0_OAI21X1_850 gnd vdd FILL
XFILL_0_OAI21X1_883 gnd vdd FILL
XFILL_1_BUFX2_8 gnd vdd FILL
XFILL_0_OAI21X1_861 gnd vdd FILL
XFILL_0_OAI21X1_872 gnd vdd FILL
XFILL_0_OAI21X1_894 gnd vdd FILL
XFILL_2_DFFPOSX1_20 gnd vdd FILL
XBUFX2_908 BUFX2_908/A gnd tid3_o[52] vdd BUFX2
XBUFX2_919 BUFX2_919/A gnd tid3_o[42] vdd BUFX2
XFILL_2_DFFPOSX1_53 gnd vdd FILL
XFILL_28_8_0 gnd vdd FILL
XFILL_2_DFFPOSX1_64 gnd vdd FILL
XFILL_2_DFFPOSX1_31 gnd vdd FILL
XFILL_3_8_0 gnd vdd FILL
XFILL_2_DFFPOSX1_42 gnd vdd FILL
XFILL_2_DFFPOSX1_75 gnd vdd FILL
XFILL_2_DFFPOSX1_86 gnd vdd FILL
XFILL_2_DFFPOSX1_97 gnd vdd FILL
XFILL_0_OAI21X1_1660 gnd vdd FILL
XFILL_29_13_1 gnd vdd FILL
XFILL_0_OAI21X1_1693 gnd vdd FILL
XFILL_0_OAI21X1_1682 gnd vdd FILL
XFILL_0_OAI21X1_1671 gnd vdd FILL
XFILL_11_7_0 gnd vdd FILL
XFILL_0_BUFX4_2 gnd vdd FILL
XFILL_0_BUFX2_615 gnd vdd FILL
XFILL_0_BUFX2_604 gnd vdd FILL
XFILL_0_BUFX2_637 gnd vdd FILL
XFILL_0_BUFX2_648 gnd vdd FILL
XFILL_0_BUFX2_626 gnd vdd FILL
XFILL_4_DFFPOSX1_1032 gnd vdd FILL
XFILL_4_DFFPOSX1_1021 gnd vdd FILL
XFILL_0_BUFX2_659 gnd vdd FILL
XFILL_4_DFFPOSX1_1010 gnd vdd FILL
XBUFX4_212 BUFX4_21/Y gnd INVX8_1/A vdd BUFX4
XBUFX4_201 BUFX4_21/Y gnd BUFX4_201/Y vdd BUFX4
XFILL_2_OAI21X1_1710 gnd vdd FILL
XBUFX4_234 BUFX4_23/Y gnd BUFX4_234/Y vdd BUFX4
XBUFX4_223 BUFX4_22/Y gnd BUFX4_223/Y vdd BUFX4
XFILL_19_8_0 gnd vdd FILL
XBUFX4_245 INVX8_1/Y gnd BUFX4_245/Y vdd BUFX4
XFILL_0_INVX2_100 gnd vdd FILL
XFILL_4_14_1 gnd vdd FILL
XFILL_0_INVX2_133 gnd vdd FILL
XBUFX4_289 BUFX4_303/A gnd BUFX4_289/Y vdd BUFX4
XFILL_0_INVX2_111 gnd vdd FILL
XBUFX4_278 INVX8_7/Y gnd BUFX4_59/A vdd BUFX4
XBUFX4_256 INVX8_5/Y gnd BUFX4_2/A vdd BUFX4
XBUFX4_267 enable_i gnd BUFX4_267/Y vdd BUFX4
XFILL_0_INVX2_144 gnd vdd FILL
XFILL_0_INVX2_122 gnd vdd FILL
XFILL_0_INVX2_155 gnd vdd FILL
XFILL_0_INVX2_177 gnd vdd FILL
XFILL_0_INVX2_166 gnd vdd FILL
XFILL_0_INVX2_199 gnd vdd FILL
XFILL_0_INVX2_188 gnd vdd FILL
XFILL_0_INVX4_2 gnd vdd FILL
XFILL_18_3 gnd vdd FILL
XOAI21X1_1102 bundleAddress_i[61] BUFX4_216/Y NAND2X1_468/Y gnd OAI21X1_1102/Y vdd
+ OAI21X1
XOAI21X1_1113 NAND2X1_476/Y NOR2X1_216/A OAI21X1_1113/C gnd OAI21X1_1114/A vdd OAI21X1
XOAI21X1_1124 NAND2X1_488/Y NOR2X1_129/Y NAND2X1_486/Y gnd OAI21X1_1124/Y vdd OAI21X1
XOAI21X1_1146 OAI21X1_1146/A XNOR2X1_64/A NAND2X1_521/Y gnd OAI21X1_1146/Y vdd OAI21X1
XFILL_1_OAI21X1_1300 gnd vdd FILL
XDFFPOSX1_714 BUFX2_369/A CLKBUF1_26/Y OAI21X1_977/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1311 gnd vdd FILL
XFILL_1_OAI21X1_1322 gnd vdd FILL
XDFFPOSX1_703 BUFX2_341/A CLKBUF1_2/Y OAI21X1_955/Y gnd vdd DFFPOSX1
XOAI21X1_1135 NOR2X1_137/Y bundleAddress_i[43] BUFX4_239/Y gnd OAI21X1_1136/A vdd
+ OAI21X1
XDFFPOSX1_747 BUFX2_24/A CLKBUF1_74/Y OAI21X1_1039/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_102 gnd vdd FILL
XDFFPOSX1_725 BUFX2_362/A CLKBUF1_43/Y OAI21X1_999/Y gnd vdd DFFPOSX1
XDFFPOSX1_736 BUFX2_374/A CLKBUF1_61/Y OAI21X1_1021/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_934 gnd vdd FILL
XFILL_1_OAI21X1_1333 gnd vdd FILL
XFILL_1_DFFPOSX1_901 gnd vdd FILL
XFILL_1_OAI21X1_1344 gnd vdd FILL
XOAI21X1_1168 NOR2X1_160/Y bundleAddress_i[21] BUFX4_239/Y gnd OAI21X1_1169/B vdd
+ OAI21X1
XOAI21X1_1179 AOI21X1_41/Y NAND2X1_566/Y NAND2X1_562/Y gnd OAI21X1_1179/Y vdd OAI21X1
XOAI21X1_1157 AND2X2_24/A bundleAddress_i[29] BUFX4_239/Y gnd OAI21X1_1158/A vdd OAI21X1
XFILL_1_OAI21X1_1366 gnd vdd FILL
XFILL_1_DFFPOSX1_923 gnd vdd FILL
XFILL_1_DFFPOSX1_912 gnd vdd FILL
XFILL_1_OAI21X1_1355 gnd vdd FILL
XFILL_1_OAI21X1_306 gnd vdd FILL
XFILL_0_OAI21X1_124 gnd vdd FILL
XDFFPOSX1_758 BUFX2_7/A CLKBUF1_59/Y OAI21X1_1050/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_146 gnd vdd FILL
XFILL_1_OAI21X1_1399 gnd vdd FILL
XFILL_0_OAI21X1_113 gnd vdd FILL
XFILL_1_DFFPOSX1_967 gnd vdd FILL
XFILL_1_OAI21X1_1388 gnd vdd FILL
XFILL_1_DFFPOSX1_945 gnd vdd FILL
XFILL_0_OAI21X1_135 gnd vdd FILL
XDFFPOSX1_769 BUFX2_19/A CLKBUF1_60/Y OAI21X1_1061/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1377 gnd vdd FILL
XFILL_1_DFFPOSX1_956 gnd vdd FILL
XFILL_1_OAI21X1_317 gnd vdd FILL
XFILL_0_OAI21X1_179 gnd vdd FILL
XFILL_0_OAI21X1_168 gnd vdd FILL
XFILL_1_DFFPOSX1_978 gnd vdd FILL
XFILL_1_OAI21X1_328 gnd vdd FILL
XFILL_1_DFFPOSX1_989 gnd vdd FILL
XFILL_0_OAI21X1_157 gnd vdd FILL
XFILL_1_OAI21X1_339 gnd vdd FILL
XFILL_9_13_1 gnd vdd FILL
XFILL_0_BUFX4_34 gnd vdd FILL
XFILL_0_BUFX4_23 gnd vdd FILL
XFILL_0_BUFX4_45 gnd vdd FILL
XFILL_0_BUFX4_12 gnd vdd FILL
XFILL_0_NAND2X1_130 gnd vdd FILL
XFILL_0_BUFX4_67 gnd vdd FILL
XFILL_1_NAND2X1_301 gnd vdd FILL
XFILL_0_BUFX4_56 gnd vdd FILL
XFILL_1_NAND2X1_323 gnd vdd FILL
XFILL_0_NAND2X1_141 gnd vdd FILL
XFILL_0_BUFX4_78 gnd vdd FILL
XFILL_0_NAND2X1_152 gnd vdd FILL
XFILL_1_NAND2X1_312 gnd vdd FILL
XFILL_1_NAND2X1_334 gnd vdd FILL
XFILL_1_BUFX4_109 gnd vdd FILL
XFILL_1_NAND2X1_345 gnd vdd FILL
XFILL_0_BUFX4_89 gnd vdd FILL
XFILL_0_DFFPOSX1_513 gnd vdd FILL
XFILL_0_DFFPOSX1_502 gnd vdd FILL
XFILL_0_NAND2X1_174 gnd vdd FILL
XFILL_0_DFFPOSX1_524 gnd vdd FILL
XFILL_0_NAND2X1_163 gnd vdd FILL
XFILL_0_NAND2X1_185 gnd vdd FILL
XFILL_1_NAND2X1_367 gnd vdd FILL
XFILL_1_NAND2X1_378 gnd vdd FILL
XFILL_0_DFFPOSX1_546 gnd vdd FILL
XFILL_0_DFFPOSX1_535 gnd vdd FILL
XFILL_0_DFFPOSX1_557 gnd vdd FILL
XFILL_0_NAND2X1_196 gnd vdd FILL
XFILL_0_DFFPOSX1_568 gnd vdd FILL
XFILL_0_DFFPOSX1_579 gnd vdd FILL
XFILL_5_DFFPOSX1_150 gnd vdd FILL
XFILL_5_DFFPOSX1_161 gnd vdd FILL
XFILL_5_DFFPOSX1_194 gnd vdd FILL
XFILL_5_DFFPOSX1_183 gnd vdd FILL
XFILL_5_DFFPOSX1_172 gnd vdd FILL
XOAI21X1_1691 BUFX4_168/Y INVX2_139/Y OAI21X1_1691/C gnd DFFPOSX1_58/D vdd OAI21X1
XOAI21X1_1680 BUFX4_11/A BUFX4_318/Y BUFX2_722/A gnd OAI21X1_1681/C vdd OAI21X1
XFILL_0_OR2X2_15 gnd vdd FILL
XFILL_1_OAI21X1_873 gnd vdd FILL
XFILL_1_OAI21X1_862 gnd vdd FILL
XFILL_1_OAI21X1_840 gnd vdd FILL
XNAND3X1_12 bundleStartMajId_i[0] INVX4_28/A NOR3X1_4/Y gnd NAND3X1_13/B vdd NAND3X1
XFILL_0_OAI21X1_680 gnd vdd FILL
XNAND3X1_23 INVX1_33/A NOR2X1_90/Y INVX2_49/A gnd NOR2X1_91/B vdd NAND3X1
XFILL_0_OAI21X1_691 gnd vdd FILL
XFILL_1_OAI21X1_851 gnd vdd FILL
XFILL_1_OAI21X1_884 gnd vdd FILL
XNAND3X1_56 AND2X2_29/B NOR2X1_196/Y INVX1_205/A gnd NOR3X1_18/A vdd NAND3X1
XNAND3X1_45 bundleAddress_i[19] NOR2X1_162/Y NOR2X1_160/Y gnd XNOR2X1_73/A vdd NAND3X1
XNAND3X1_34 bundleStartMajId_i[8] INVX2_46/A NOR3X1_8/Y gnd NAND3X1_34/Y vdd NAND3X1
XFILL_1_OAI21X1_895 gnd vdd FILL
XFILL_2_OAI21X1_1006 gnd vdd FILL
XNAND3X1_67 INVX4_51/A AND2X2_23/B AND2X2_24/B gnd OR2X2_21/A vdd NAND3X1
XNOR2X1_12 OR2X2_5/A INVX1_10/A gnd NOR2X1_12/Y vdd NOR2X1
XFILL_3_DFFPOSX1_10 gnd vdd FILL
XFILL_3_DFFPOSX1_21 gnd vdd FILL
XFILL_3_DFFPOSX1_32 gnd vdd FILL
XFILL_3_DFFPOSX1_43 gnd vdd FILL
XBUFX2_716 BUFX2_716/A gnd pid3_o[20] vdd BUFX2
XBUFX2_727 BUFX2_727/A gnd pid3_o[10] vdd BUFX2
XNOR2X1_45 bundleStartMajId_i[13] NOR2X1_45/B gnd NOR2X1_45/Y vdd NOR2X1
XFILL_2_DFFPOSX1_607 gnd vdd FILL
XNOR2X1_34 NOR3X1_6/B NOR2X1_34/B gnd AND2X2_7/B vdd NOR2X1
XFILL_2_DFFPOSX1_629 gnd vdd FILL
XFILL_2_DFFPOSX1_618 gnd vdd FILL
XBUFX2_705 BUFX2_705/A gnd pid2_o[1] vdd BUFX2
XNOR2X1_23 NOR2X1_23/A NOR3X1_9/C gnd INVX1_16/A vdd NOR2X1
XFILL_3_DFFPOSX1_76 gnd vdd FILL
XNOR2X1_56 bundleStartMajId_i[2] NOR3X1_4/Y gnd NOR2X1_56/Y vdd NOR2X1
XFILL_3_DFFPOSX1_54 gnd vdd FILL
XBUFX2_749 BUFX2_749/A gnd pid4_o[19] vdd BUFX2
XNOR2X1_78 OR2X2_9/B OR2X2_9/A gnd OAI22X1_2/C vdd NOR2X1
XFILL_3_DFFPOSX1_65 gnd vdd FILL
XNOR2X1_67 OR2X2_5/A OR2X2_2/B gnd NOR2X1_67/Y vdd NOR2X1
XBUFX2_738 BUFX2_738/A gnd pid3_o[0] vdd BUFX2
XFILL_3_DFFPOSX1_87 gnd vdd FILL
XNOR2X1_89 NOR2X1_89/A NOR2X1_89/B gnd NOR2X1_89/Y vdd NOR2X1
XFILL_3_DFFPOSX1_98 gnd vdd FILL
XFILL_0_OAI21X1_1490 gnd vdd FILL
XFILL_0_BUFX2_412 gnd vdd FILL
XFILL_0_BUFX2_423 gnd vdd FILL
XINVX2_201 bundleTid_i[8] gnd INVX2_201/Y vdd INVX2
XFILL_0_BUFX2_401 gnd vdd FILL
XFILL_1_DFFPOSX1_208 gnd vdd FILL
XFILL_1_DFFPOSX1_219 gnd vdd FILL
XFILL_0_BUFX2_445 gnd vdd FILL
XFILL_0_BUFX2_434 gnd vdd FILL
XFILL_0_BUFX2_456 gnd vdd FILL
XFILL_0_BUFX2_489 gnd vdd FILL
XFILL_0_BUFX2_478 gnd vdd FILL
XFILL_0_BUFX2_467 gnd vdd FILL
XFILL_14_14_0 gnd vdd FILL
XFILL_0_NAND2X1_10 gnd vdd FILL
XFILL_0_NAND2X1_21 gnd vdd FILL
XFILL_0_NAND2X1_32 gnd vdd FILL
XNOR2X1_124 INVX1_183/A NOR2X1_124/B gnd INVX4_47/A vdd NOR2X1
XFILL_0_NAND2X1_65 gnd vdd FILL
XFILL_0_NAND2X1_43 gnd vdd FILL
XNOR2X1_113 NOR3X1_6/A AND2X2_21/A gnd NOR2X1_113/Y vdd NOR2X1
XFILL_0_NAND2X1_54 gnd vdd FILL
XNOR2X1_102 NOR2X1_4/A INVX2_52/Y gnd INVX1_34/A vdd NOR2X1
XFILL_34_6_0 gnd vdd FILL
XNOR2X1_146 bundleAddress_i[33] NOR2X1_146/B gnd NOR2X1_146/Y vdd NOR2X1
XFILL_0_NAND2X1_98 gnd vdd FILL
XNOR2X1_135 OR2X2_18/A INVX1_187/A gnd NOR2X1_138/B vdd NOR2X1
XFILL_0_NAND2X1_76 gnd vdd FILL
XFILL_0_NAND2X1_87 gnd vdd FILL
XNOR2X1_157 NOR3X1_16/B INVX1_193/A gnd NOR2X1_157/Y vdd NOR2X1
XNOR2X1_179 INVX2_62/Y INVX2_93/Y gnd XNOR2X1_75/A vdd NOR2X1
XFILL_23_1 gnd vdd FILL
XNOR2X1_168 INVX2_84/Y INVX2_85/Y gnd INVX2_103/A vdd NOR2X1
XOAI21X1_608 OAI21X1_608/A AOI21X1_13/Y OAI21X1_608/C gnd OAI21X1_608/Y vdd OAI21X1
XOAI21X1_619 INVX2_50/Y INVX1_33/Y NOR2X1_89/B gnd OAI21X1_620/A vdd OAI21X1
XFILL_1_OAI21X1_1130 gnd vdd FILL
XFILL_1_OAI21X1_1141 gnd vdd FILL
XDFFPOSX1_500 BUFX2_529/A CLKBUF1_46/Y OAI21X1_546/Y gnd vdd DFFPOSX1
XDFFPOSX1_522 BUFX2_553/A CLKBUF1_33/Y OAI21X1_602/Y gnd vdd DFFPOSX1
XDFFPOSX1_511 BUFX2_541/A CLKBUF1_63/Y OAI21X1_574/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_742 gnd vdd FILL
XDFFPOSX1_544 BUFX2_578/A CLKBUF1_29/Y OAI21X1_651/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1152 gnd vdd FILL
XFILL_1_OAI21X1_1174 gnd vdd FILL
XDFFPOSX1_555 BUFX2_646/A CLKBUF1_91/Y OAI21X1_681/Y gnd vdd DFFPOSX1
XDFFPOSX1_533 BUFX2_565/A CLKBUF1_87/Y OAI21X1_625/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_720 gnd vdd FILL
XFILL_1_DFFPOSX1_731 gnd vdd FILL
XFILL_1_OAI21X1_1163 gnd vdd FILL
XFILL_1_OAI21X1_103 gnd vdd FILL
XFILL_1_OAI21X1_125 gnd vdd FILL
XFILL_1_OAI21X1_114 gnd vdd FILL
XFILL_1_DFFPOSX1_753 gnd vdd FILL
XFILL_1_DFFPOSX1_775 gnd vdd FILL
XDFFPOSX1_599 BUFX2_632/A CLKBUF1_72/Y OAI21X1_809/Y gnd vdd DFFPOSX1
XNAND2X1_603 bundleAddress_i[38] bundleAddress_i[37] gnd OR2X2_19/B vdd NAND2X1
XDFFPOSX1_588 BUFX2_620/A CLKBUF1_1/Y OAI21X1_772/Y gnd vdd DFFPOSX1
XDFFPOSX1_566 BUFX2_595/A CLKBUF1_88/Y OAI21X1_711/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1196 gnd vdd FILL
XDFFPOSX1_577 BUFX2_607/A CLKBUF1_63/Y OAI21X1_743/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1185 gnd vdd FILL
XFILL_0_BUFX2_990 gnd vdd FILL
XFILL_1_DFFPOSX1_764 gnd vdd FILL
XFILL_1_OAI21X1_158 gnd vdd FILL
XFILL_1_OAI21X1_147 gnd vdd FILL
XNAND2X1_625 NAND2X1_625/A INVX2_108/Y gnd NAND2X1_625/Y vdd NAND2X1
XNAND2X1_636 INVX1_223/A NAND2X1_636/B gnd NAND2X1_636/Y vdd NAND2X1
XFILL_1_INVX2_109 gnd vdd FILL
XFILL_19_13_0 gnd vdd FILL
XFILL_1_DFFPOSX1_786 gnd vdd FILL
XNAND2X1_614 AND2X2_31/B NOR2X1_201/Y gnd NOR3X1_17/B vdd NAND2X1
XFILL_1_DFFPOSX1_797 gnd vdd FILL
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XFILL_1_OAI21X1_136 gnd vdd FILL
XFILL_2_OAI21X1_318 gnd vdd FILL
XNAND2X1_658 BUFX2_679/A BUFX4_349/Y gnd NAND2X1_658/Y vdd NAND2X1
XFILL_1_OAI21X1_169 gnd vdd FILL
XNAND2X1_647 NAND3X1_69/Y NAND2X1_647/B gnd NAND2X1_647/Y vdd NAND2X1
XNAND2X1_669 BUFX2_660/A BUFX4_321/Y gnd NAND2X1_669/Y vdd NAND2X1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XINVX1_26 NOR2X1_8/Y gnd INVX1_26/Y vdd INVX1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XINVX1_59 INVX1_59/A gnd INVX1_59/Y vdd INVX1
XFILL_6_DFFPOSX1_390 gnd vdd FILL
XFILL_32_15_0 gnd vdd FILL
XFILL_1_NAND2X1_131 gnd vdd FILL
XFILL_25_6_0 gnd vdd FILL
XFILL_0_XNOR2X1_100 gnd vdd FILL
XFILL_0_6_0 gnd vdd FILL
XFILL_0_DFFPOSX1_321 gnd vdd FILL
XFILL_0_DFFPOSX1_310 gnd vdd FILL
XFILL_0_DFFPOSX1_332 gnd vdd FILL
XFILL_1_NAND2X1_164 gnd vdd FILL
XFILL_1_NAND2X1_153 gnd vdd FILL
XFILL_0_DFFPOSX1_343 gnd vdd FILL
XFILL_1_NAND2X1_175 gnd vdd FILL
XFILL_0_DFFPOSX1_354 gnd vdd FILL
XFILL_0_DFFPOSX1_365 gnd vdd FILL
XFILL_0_DFFPOSX1_398 gnd vdd FILL
XFILL_0_DFFPOSX1_376 gnd vdd FILL
XFILL_0_DFFPOSX1_387 gnd vdd FILL
XFILL_3_DFFPOSX1_814 gnd vdd FILL
XFILL_3_DFFPOSX1_803 gnd vdd FILL
XFILL_3_DFFPOSX1_825 gnd vdd FILL
XFILL_3_DFFPOSX1_836 gnd vdd FILL
XFILL_3_DFFPOSX1_847 gnd vdd FILL
XFILL_3_DFFPOSX1_869 gnd vdd FILL
XFILL_3_DFFPOSX1_858 gnd vdd FILL
XFILL_37_14_0 gnd vdd FILL
XFILL_1_NOR2X1_220 gnd vdd FILL
XFILL_8_7_0 gnd vdd FILL
XFILL_1_OAI21X1_681 gnd vdd FILL
XFILL_1_OAI21X1_670 gnd vdd FILL
XFILL_1_OAI21X1_692 gnd vdd FILL
XFILL_2_OAI21X1_874 gnd vdd FILL
XFILL_1_INVX1_153 gnd vdd FILL
XFILL_1_INVX1_186 gnd vdd FILL
XFILL_2_DFFPOSX1_404 gnd vdd FILL
XBUFX2_502 BUFX2_502/A gnd majID2_o[58] vdd BUFX2
XFILL_4_DFFPOSX1_11 gnd vdd FILL
XFILL_2_DFFPOSX1_415 gnd vdd FILL
XFILL_4_DFFPOSX1_22 gnd vdd FILL
XFILL_4_DFFPOSX1_33 gnd vdd FILL
XBUFX2_524 BUFX2_524/A gnd majID3_o[52] vdd BUFX2
XBUFX2_535 MUX2X1_1/B gnd majID3_o[42] vdd BUFX2
XBUFX2_513 BUFX2_513/A gnd majID2_o[57] vdd BUFX2
XFILL_2_DFFPOSX1_426 gnd vdd FILL
XFILL_2_DFFPOSX1_437 gnd vdd FILL
XBUFX2_579 BUFX2_579/A gnd majID3_o[2] vdd BUFX2
XFILL_4_DFFPOSX1_44 gnd vdd FILL
XBUFX2_546 BUFX2_546/A gnd majID3_o[32] vdd BUFX2
XBUFX2_568 BUFX2_568/A gnd majID3_o[12] vdd BUFX2
XBUFX2_557 BUFX2_557/A gnd majID3_o[22] vdd BUFX2
XFILL_2_DFFPOSX1_459 gnd vdd FILL
XFILL_4_DFFPOSX1_55 gnd vdd FILL
XFILL_16_6_0 gnd vdd FILL
XFILL_4_DFFPOSX1_66 gnd vdd FILL
XFILL_2_DFFPOSX1_448 gnd vdd FILL
XFILL_4_DFFPOSX1_77 gnd vdd FILL
XFILL_4_DFFPOSX1_88 gnd vdd FILL
XFILL_4_DFFPOSX1_99 gnd vdd FILL
XFILL_5_DFFPOSX1_919 gnd vdd FILL
XFILL_5_DFFPOSX1_908 gnd vdd FILL
XFILL_0_BUFX2_220 gnd vdd FILL
XFILL_0_BUFX2_231 gnd vdd FILL
XFILL_0_BUFX2_264 gnd vdd FILL
XFILL_0_BUFX2_253 gnd vdd FILL
XFILL_0_BUFX2_242 gnd vdd FILL
XFILL_0_BUFX2_297 gnd vdd FILL
XFILL_0_BUFX2_286 gnd vdd FILL
XFILL_0_BUFX2_275 gnd vdd FILL
XFILL_4_DFFPOSX1_509 gnd vdd FILL
XFILL_2_OAI21X1_1392 gnd vdd FILL
XFILL_2_DFFPOSX1_960 gnd vdd FILL
XFILL_2_DFFPOSX1_982 gnd vdd FILL
XFILL_2_DFFPOSX1_993 gnd vdd FILL
XFILL_2_DFFPOSX1_971 gnd vdd FILL
XFILL_0_NAND3X1_5 gnd vdd FILL
XOAI21X1_405 INVX2_40/Y NOR2X1_4/A INVX4_2/Y gnd OAI21X1_406/C vdd OAI21X1
XOAI21X1_438 NOR3X1_1/C INVX1_12/Y INVX2_22/Y gnd OAI21X1_438/Y vdd OAI21X1
XOAI21X1_427 OAI21X1_427/A NOR2X1_12/Y OAI21X1_427/C gnd OAI21X1_427/Y vdd OAI21X1
XOAI21X1_416 XNOR2X1_2/Y BUFX4_225/Y OAI21X1_416/C gnd OAI21X1_416/Y vdd OAI21X1
XOAI21X1_449 INVX1_15/Y OAI21X1_449/B OAI21X1_449/C gnd OAI21X1_449/Y vdd OAI21X1
XFILL_21_12_1 gnd vdd FILL
XFILL_3_XNOR2X1_40 gnd vdd FILL
XDFFPOSX1_330 BUFX2_1001/A CLKBUF1_17/Y OAI21X1_277/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_73 gnd vdd FILL
XFILL_3_XNOR2X1_84 gnd vdd FILL
XDFFPOSX1_341 BUFX2_1013/A CLKBUF1_8/Y OAI21X1_299/Y gnd vdd DFFPOSX1
XDFFPOSX1_374 BUFX2_403/A CLKBUF1_19/Y OAI21X1_346/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_550 gnd vdd FILL
XFILL_3_XNOR2X1_95 gnd vdd FILL
XDFFPOSX1_352 BUFX2_1026/A CLKBUF1_83/Y OAI21X1_321/Y gnd vdd DFFPOSX1
XDFFPOSX1_363 BUFX2_454/A CLKBUF1_66/Y OAI21X1_335/Y gnd vdd DFFPOSX1
XNAND2X1_411 BUFX2_64/A BUFX4_382/Y gnd NAND2X1_411/Y vdd NAND2X1
XFILL_1_DFFPOSX1_583 gnd vdd FILL
XDFFPOSX1_396 BUFX2_428/A CLKBUF1_80/Y OAI21X1_368/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_572 gnd vdd FILL
XDFFPOSX1_385 BUFX2_415/A CLKBUF1_63/Y OAI21X1_357/Y gnd vdd DFFPOSX1
XNAND2X1_400 BUFX2_317/A BUFX4_228/Y gnd OAI21X1_906/C vdd NAND2X1
XFILL_1_DFFPOSX1_561 gnd vdd FILL
XNAND2X1_433 BUFX2_26/A BUFX4_341/Y gnd NAND2X1_433/Y vdd NAND2X1
XNAND2X1_444 BUFX2_38/A BUFX4_342/Y gnd NAND2X1_444/Y vdd NAND2X1
XFILL_1_DFFPOSX1_594 gnd vdd FILL
XNAND2X1_422 BUFX2_14/A BUFX4_354/Y gnd NAND2X1_422/Y vdd NAND2X1
XNAND2X1_466 BUFX2_65/A BUFX4_234/Y gnd NAND2X1_466/Y vdd NAND2X1
XNAND2X1_488 BUFX4_241/Y NAND2X1_488/B gnd NAND2X1_488/Y vdd NAND2X1
XNAND2X1_477 bundleAddress_i[57] bundleAddress_i[56] gnd NOR2X1_216/A vdd NAND2X1
XNAND2X1_455 BUFX2_50/A NAND2X1_7/B gnd NAND2X1_455/Y vdd NAND2X1
XNAND2X1_499 BUFX2_74/A OAI21X1_8/B gnd NAND2X1_499/Y vdd NAND2X1
XFILL_0_INVX1_209 gnd vdd FILL
XFILL_1_XNOR2X1_101 gnd vdd FILL
XFILL_0_DFFPOSX1_140 gnd vdd FILL
XFILL_0_DFFPOSX1_173 gnd vdd FILL
XFILL_0_DFFPOSX1_151 gnd vdd FILL
XFILL_0_DFFPOSX1_162 gnd vdd FILL
XFILL_0_DFFPOSX1_184 gnd vdd FILL
XFILL_1_BUFX2_900 gnd vdd FILL
XFILL_1_BUFX2_944 gnd vdd FILL
XFILL_1_BUFX2_933 gnd vdd FILL
XFILL_0_OAI21X1_19 gnd vdd FILL
XFILL_1_BUFX2_955 gnd vdd FILL
XFILL_26_11_1 gnd vdd FILL
XFILL_0_DFFPOSX1_195 gnd vdd FILL
XFILL_1_BUFX2_988 gnd vdd FILL
XOAI21X1_950 BUFX4_8/Y BUFX4_368/Y BUFX2_339/A gnd OAI21X1_951/C vdd OAI21X1
XFILL_1_BUFX2_977 gnd vdd FILL
XFILL_3_DFFPOSX1_600 gnd vdd FILL
XFILL_3_DFFPOSX1_611 gnd vdd FILL
XFILL_3_DFFPOSX1_622 gnd vdd FILL
XOAI21X1_961 BUFX4_153/Y INVX1_135/Y OAI21X1_961/C gnd OAI21X1_961/Y vdd OAI21X1
XFILL_1_BUFX2_999 gnd vdd FILL
XFILL_3_DFFPOSX1_655 gnd vdd FILL
XFILL_3_DFFPOSX1_633 gnd vdd FILL
XFILL_3_DFFPOSX1_644 gnd vdd FILL
XOAI21X1_983 BUFX4_294/Y INVX1_146/Y OAI21X1_983/C gnd OAI21X1_983/Y vdd OAI21X1
XOAI21X1_994 BUFX4_177/Y BUFX4_74/Y BUFX2_360/A gnd OAI21X1_995/C vdd OAI21X1
XOAI21X1_972 BUFX4_133/Y BUFX4_56/Y BUFX2_357/A gnd OAI21X1_973/C vdd OAI21X1
XFILL_3_DFFPOSX1_688 gnd vdd FILL
XFILL_3_DFFPOSX1_677 gnd vdd FILL
XFILL_3_DFFPOSX1_666 gnd vdd FILL
XFILL_3_DFFPOSX1_699 gnd vdd FILL
XINVX2_91 bundleAddress_i[2] gnd INVX2_91/Y vdd INVX2
XINVX2_80 bundleAddress_i[21] gnd INVX2_80/Y vdd INVX2
XBUFX2_310 BUFX2_310/A gnd instr2_o[7] vdd BUFX2
XFILL_2_DFFPOSX1_212 gnd vdd FILL
XFILL_2_DFFPOSX1_201 gnd vdd FILL
XFILL_0_NAND2X1_707 gnd vdd FILL
XFILL_0_NAND2X1_718 gnd vdd FILL
XFILL_2_DFFPOSX1_245 gnd vdd FILL
XFILL_0_NAND2X1_729 gnd vdd FILL
XFILL_5_DFFPOSX1_12 gnd vdd FILL
XFILL_2_DFFPOSX1_234 gnd vdd FILL
XBUFX2_321 BUFX2_321/A gnd instr2_o[25] vdd BUFX2
XBUFX2_354 BUFX2_354/A gnd instr3_o[24] vdd BUFX2
XBUFX2_332 BUFX2_332/A gnd instr3_o[16] vdd BUFX2
XFILL_1_12_1 gnd vdd FILL
XFILL_2_DFFPOSX1_223 gnd vdd FILL
XFILL_2_DFFPOSX1_256 gnd vdd FILL
XBUFX2_343 BUFX2_343/A gnd instr3_o[6] vdd BUFX2
XFILL_2_DFFPOSX1_278 gnd vdd FILL
XFILL_5_DFFPOSX1_45 gnd vdd FILL
XFILL_2_DFFPOSX1_289 gnd vdd FILL
XFILL_2_DFFPOSX1_267 gnd vdd FILL
XBUFX2_376 BUFX2_376/A gnd instr4_o[5] vdd BUFX2
XFILL_5_DFFPOSX1_23 gnd vdd FILL
XFILL_5_DFFPOSX1_34 gnd vdd FILL
XBUFX2_387 BUFX2_387/A gnd instr4_o[23] vdd BUFX2
XBUFX2_365 BUFX2_365/A gnd instr4_o[15] vdd BUFX2
XFILL_5_DFFPOSX1_78 gnd vdd FILL
XFILL_32_9_1 gnd vdd FILL
XFILL_5_DFFPOSX1_89 gnd vdd FILL
XFILL_5_DFFPOSX1_56 gnd vdd FILL
XFILL_1_NOR3X1_15 gnd vdd FILL
XOAI21X1_10 INVX2_148/Y BUFX4_233/Y OAI21X1_10/C gnd OAI21X1_10/Y vdd OAI21X1
XBUFX2_398 BUFX2_398/A gnd majID1_o[50] vdd BUFX2
XFILL_5_DFFPOSX1_67 gnd vdd FILL
XOAI21X1_32 INVX2_170/Y BUFX4_207/Y OAI21X1_32/C gnd OAI21X1_32/Y vdd OAI21X1
XFILL_31_4_0 gnd vdd FILL
XFILL_5_DFFPOSX1_716 gnd vdd FILL
XFILL_5_DFFPOSX1_727 gnd vdd FILL
XOAI21X1_43 INVX2_181/Y BUFX4_183/Y OAI21X1_43/C gnd OAI21X1_43/Y vdd OAI21X1
XOAI21X1_54 INVX2_192/Y BUFX4_222/Y OAI21X1_54/C gnd OAI21X1_54/Y vdd OAI21X1
XOAI21X1_21 INVX2_159/Y BUFX4_237/Y OAI21X1_21/C gnd OAI21X1_21/Y vdd OAI21X1
XFILL_5_DFFPOSX1_705 gnd vdd FILL
XFILL_5_DFFPOSX1_749 gnd vdd FILL
XOAI21X1_65 INVX2_1/Y BUFX4_223/Y OAI21X1_65/C gnd OAI21X1_65/Y vdd OAI21X1
XFILL_1_BUFX4_281 gnd vdd FILL
XFILL_1_BUFX4_270 gnd vdd FILL
XOAI21X1_87 BUFX4_162/Y INVX2_153/Y OAI21X1_87/C gnd OAI21X1_87/Y vdd OAI21X1
XOAI21X1_76 BUFX4_101/Y BUFX4_373/Y BUFX2_917/A gnd OAI21X1_77/C vdd OAI21X1
XFILL_5_DFFPOSX1_738 gnd vdd FILL
XFILL_1_BUFX4_292 gnd vdd FILL
XOAI21X1_98 BUFX4_7/A BUFX4_315/Y BUFX2_910/A gnd OAI21X1_99/C vdd OAI21X1
XFILL_4_DFFPOSX1_306 gnd vdd FILL
XFILL_0_DFFPOSX1_30 gnd vdd FILL
XFILL_0_DFFPOSX1_52 gnd vdd FILL
XFILL_4_DFFPOSX1_317 gnd vdd FILL
XFILL_0_DFFPOSX1_41 gnd vdd FILL
XFILL_4_DFFPOSX1_328 gnd vdd FILL
XFILL_4_DFFPOSX1_339 gnd vdd FILL
XFILL_0_DFFPOSX1_85 gnd vdd FILL
XFILL_0_DFFPOSX1_63 gnd vdd FILL
XFILL_6_11_1 gnd vdd FILL
XFILL_0_DFFPOSX1_74 gnd vdd FILL
XFILL_0_DFFPOSX1_96 gnd vdd FILL
XFILL_2_DFFPOSX1_1009 gnd vdd FILL
XFILL_2_DFFPOSX1_790 gnd vdd FILL
XFILL_23_9_1 gnd vdd FILL
XFILL_1_BUFX2_218 gnd vdd FILL
XFILL_22_4_0 gnd vdd FILL
XOAI21X1_213 INVX2_152/Y INVX8_2/A OAI21X1_213/C gnd OAI21X1_213/Y vdd OAI21X1
XFILL_1_BUFX2_229 gnd vdd FILL
XOAI21X1_202 BUFX4_169/Y BUFX4_78/Y BUFX2_970/A gnd OAI21X1_203/C vdd OAI21X1
XOAI21X1_224 BUFX4_165/Y BUFX4_34/Y BUFX2_973/A gnd OAI21X1_225/C vdd OAI21X1
XOAI21X1_235 INVX2_163/Y BUFX4_289/Y OAI21X1_235/C gnd OAI21X1_235/Y vdd OAI21X1
XOAI21X1_246 BUFX4_172/Y BUFX4_50/Y BUFX2_985/A gnd OAI21X1_247/C vdd OAI21X1
XOAI21X1_268 BUFX4_172/Y BUFX4_66/Y BUFX2_997/A gnd OAI21X1_269/C vdd OAI21X1
XOAI21X1_279 INVX2_185/Y BUFX4_297/Y OAI21X1_279/C gnd OAI21X1_279/Y vdd OAI21X1
XOAI21X1_257 INVX2_174/Y BUFX4_303/Y OAI21X1_257/C gnd OAI21X1_257/Y vdd OAI21X1
XAND2X2_13 NOR2X1_62/Y INVX4_30/A gnd AND2X2_13/Y vdd AND2X2
XAND2X2_24 AND2X2_24/A AND2X2_24/B gnd AND2X2_24/Y vdd AND2X2
XDFFPOSX1_171 BUFX2_902/A CLKBUF1_26/Y OAI21X1_15/Y gnd vdd DFFPOSX1
XDFFPOSX1_182 BUFX2_851/A CLKBUF1_30/Y OAI21X1_26/Y gnd vdd DFFPOSX1
XFILL_0_NOR3X1_3 gnd vdd FILL
XDFFPOSX1_160 NAND2X1_4/A CLKBUF1_52/Y OAI21X1_4/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_391 gnd vdd FILL
XFILL_1_DFFPOSX1_380 gnd vdd FILL
XDFFPOSX1_193 BUFX2_863/A CLKBUF1_76/Y OAI21X1_37/Y gnd vdd DFFPOSX1
XNAND2X1_241 bundleStartMajId_i[13] NOR2X1_45/B gnd XNOR2X1_21/A vdd NAND2X1
XNAND2X1_252 NOR2X1_53/Y NOR2X1_52/Y gnd XNOR2X1_23/A vdd NAND2X1
XNAND2X1_230 bundleStartMajId_i[20] bundleStartMajId_i[19] gnd NOR3X1_3/B vdd NAND2X1
XFILL_4_DFFPOSX1_840 gnd vdd FILL
XNAND2X1_263 BUFX2_516/A BUFX4_221/Y gnd OAI21X1_498/C vdd NAND2X1
XNAND2X1_296 INVX1_32/Y NOR2X1_84/Y gnd OAI21X1_610/A vdd NAND2X1
XNAND2X1_285 bundleStartMajId_i[34] bundleStartMajId_i[33] gnd NOR2X1_74/A vdd NAND2X1
XNAND2X1_274 OAI21X1_539/Y XNOR2X1_27/A gnd OAI21X1_541/A vdd NAND2X1
XFILL_5_5_0 gnd vdd FILL
XFILL_4_DFFPOSX1_851 gnd vdd FILL
XFILL_4_DFFPOSX1_873 gnd vdd FILL
XFILL_4_DFFPOSX1_862 gnd vdd FILL
XFILL_4_DFFPOSX1_884 gnd vdd FILL
XFILL_12_17_1 gnd vdd FILL
XFILL_4_DFFPOSX1_895 gnd vdd FILL
XFILL_0_OAI21X1_2 gnd vdd FILL
XFILL_14_9_1 gnd vdd FILL
XFILL_2_XNOR2X1_102 gnd vdd FILL
XFILL_13_4_0 gnd vdd FILL
XFILL_1_BUFX2_730 gnd vdd FILL
XFILL_1_BUFX2_752 gnd vdd FILL
XFILL_0_BUFX4_304 gnd vdd FILL
XFILL_1_NOR2X1_70 gnd vdd FILL
XFILL_0_BUFX4_315 gnd vdd FILL
XFILL_1_BUFX2_741 gnd vdd FILL
XFILL_1_BUFX2_796 gnd vdd FILL
XFILL_1_BUFX2_785 gnd vdd FILL
XFILL_1_NOR2X1_92 gnd vdd FILL
XFILL_0_BUFX4_348 gnd vdd FILL
XOAI21X1_1509 OAI21X1_1509/A BUFX4_297/Y OAI21X1_1509/C gnd OAI21X1_1509/Y vdd OAI21X1
XFILL_3_DFFPOSX1_430 gnd vdd FILL
XFILL_1_OAI21X1_1707 gnd vdd FILL
XFILL_0_BUFX4_326 gnd vdd FILL
XFILL_0_BUFX4_337 gnd vdd FILL
XFILL_0_BUFX4_359 gnd vdd FILL
XFILL_1_OAI21X1_1729 gnd vdd FILL
XFILL_3_DFFPOSX1_463 gnd vdd FILL
XOAI21X1_780 NOR3X1_2/B NOR2X1_114/B OAI21X1_780/C gnd OAI21X1_782/A vdd OAI21X1
XFILL_1_OAI21X1_1718 gnd vdd FILL
XOAI21X1_791 INVX4_31/Y OAI21X1_793/B BUFX4_285/Y gnd OAI21X1_792/B vdd OAI21X1
XFILL_3_DFFPOSX1_452 gnd vdd FILL
XFILL_3_DFFPOSX1_441 gnd vdd FILL
XFILL_3_DFFPOSX1_474 gnd vdd FILL
XFILL_3_DFFPOSX1_485 gnd vdd FILL
XFILL_0_OAI21X1_509 gnd vdd FILL
XFILL_3_DFFPOSX1_496 gnd vdd FILL
XFILL_0_BUFX2_1008 gnd vdd FILL
XFILL_0_BUFX2_1019 gnd vdd FILL
XFILL_6_DFFPOSX1_945 gnd vdd FILL
XFILL_6_DFFPOSX1_934 gnd vdd FILL
XFILL_6_DFFPOSX1_923 gnd vdd FILL
XFILL_6_DFFPOSX1_967 gnd vdd FILL
XFILL_17_16_1 gnd vdd FILL
XFILL_6_DFFPOSX1_978 gnd vdd FILL
XFILL_6_DFFPOSX1_956 gnd vdd FILL
XFILL_6_3 gnd vdd FILL
XFILL_2_OAI21X1_490 gnd vdd FILL
XFILL_0_NAND2X1_515 gnd vdd FILL
XFILL_30_18_1 gnd vdd FILL
XFILL_0_NAND2X1_526 gnd vdd FILL
XFILL_11_12_0 gnd vdd FILL
XFILL_0_NAND2X1_504 gnd vdd FILL
XFILL_2_XNOR2X1_92 gnd vdd FILL
XFILL_0_NAND2X1_559 gnd vdd FILL
XFILL_2_XNOR2X1_81 gnd vdd FILL
XBUFX2_151 BUFX2_151/A gnd addr3_o[34] vdd BUFX2
XBUFX2_162 BUFX2_162/A gnd addr3_o[24] vdd BUFX2
XFILL_0_NAND2X1_537 gnd vdd FILL
XFILL_0_NAND2X1_548 gnd vdd FILL
XBUFX2_140 BUFX2_140/A gnd addr3_o[44] vdd BUFX2
XFILL_2_XNOR2X1_70 gnd vdd FILL
XFILL_0_OAI21X1_1319 gnd vdd FILL
XFILL_0_OAI21X1_1308 gnd vdd FILL
XFILL_6_DFFPOSX1_13 gnd vdd FILL
XBUFX2_195 BUFX2_195/A gnd addr4_o[53] vdd BUFX2
XFILL_6_DFFPOSX1_24 gnd vdd FILL
XBUFX2_173 BUFX2_173/A gnd addr3_o[14] vdd BUFX2
XBUFX2_184 BUFX2_184/A gnd addr3_o[4] vdd BUFX2
XFILL_0_DFFPOSX1_909 gnd vdd FILL
XFILL_1_NAND2X1_3 gnd vdd FILL
XFILL_6_DFFPOSX1_35 gnd vdd FILL
XFILL_6_DFFPOSX1_68 gnd vdd FILL
XFILL_6_DFFPOSX1_57 gnd vdd FILL
XFILL_6_DFFPOSX1_46 gnd vdd FILL
XFILL_5_DFFPOSX1_502 gnd vdd FILL
XFILL_5_DFFPOSX1_535 gnd vdd FILL
XFILL_5_DFFPOSX1_513 gnd vdd FILL
XFILL_5_DFFPOSX1_524 gnd vdd FILL
XFILL_5_DFFPOSX1_546 gnd vdd FILL
XFILL_5_DFFPOSX1_568 gnd vdd FILL
XFILL_5_DFFPOSX1_579 gnd vdd FILL
XFILL_5_DFFPOSX1_557 gnd vdd FILL
XBUFX2_1021 BUFX2_1021/A gnd tid4_o[7] vdd BUFX2
XBUFX2_1010 BUFX2_1010/A gnd tid4_o[17] vdd BUFX2
XBUFX2_1032 BUFX2_1032/A gnd tid4_o[54] vdd BUFX2
XFILL_1_AOI21X1_8 gnd vdd FILL
XFILL_35_17_1 gnd vdd FILL
XCLKBUF1_11 BUFX4_84/Y gnd CLKBUF1_11/Y vdd CLKBUF1
XCLKBUF1_22 BUFX4_83/Y gnd CLKBUF1_22/Y vdd CLKBUF1
XCLKBUF1_33 BUFX4_91/Y gnd CLKBUF1_33/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_114 gnd vdd FILL
XFILL_4_DFFPOSX1_125 gnd vdd FILL
XFILL_1_DFFPOSX1_20 gnd vdd FILL
XFILL_4_DFFPOSX1_136 gnd vdd FILL
XCLKBUF1_55 BUFX4_86/Y gnd CLKBUF1_55/Y vdd CLKBUF1
XFILL_16_11_0 gnd vdd FILL
XCLKBUF1_44 BUFX4_84/Y gnd CLKBUF1_44/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_103 gnd vdd FILL
XFILL_1_DFFPOSX1_31 gnd vdd FILL
XFILL_1_DFFPOSX1_42 gnd vdd FILL
XCLKBUF1_66 BUFX4_90/Y gnd CLKBUF1_66/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_75 gnd vdd FILL
XCLKBUF1_99 BUFX4_87/Y gnd CLKBUF1_99/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_147 gnd vdd FILL
XFILL_1_DFFPOSX1_53 gnd vdd FILL
XFILL_1_DFFPOSX1_64 gnd vdd FILL
XCLKBUF1_88 BUFX4_91/Y gnd CLKBUF1_88/Y vdd CLKBUF1
XCLKBUF1_77 BUFX4_88/Y gnd CLKBUF1_77/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_158 gnd vdd FILL
XFILL_4_DFFPOSX1_169 gnd vdd FILL
XFILL_2_BUFX4_235 gnd vdd FILL
XFILL_2_BUFX4_202 gnd vdd FILL
XFILL_1_DFFPOSX1_86 gnd vdd FILL
XFILL_1_DFFPOSX1_97 gnd vdd FILL
XFILL_0_OAI21X1_1820 gnd vdd FILL
XFILL_0_BUFX2_808 gnd vdd FILL
XFILL_0_BUFX2_819 gnd vdd FILL
XINVX1_107 bundle_i[33] gnd INVX1_107/Y vdd INVX1
XINVX1_129 bundle_i[75] gnd INVX1_129/Y vdd INVX1
XINVX1_118 bundle_i[86] gnd INVX1_118/Y vdd INVX1
XFILL_3_XNOR2X1_6 gnd vdd FILL
XFILL_6_DFFPOSX1_208 gnd vdd FILL
XFILL_6_DFFPOSX1_219 gnd vdd FILL
XFILL_34_12_0 gnd vdd FILL
XFILL_0_INVX2_28 gnd vdd FILL
XFILL_0_INVX2_17 gnd vdd FILL
XFILL_0_INVX2_39 gnd vdd FILL
XFILL_4_DFFPOSX1_670 gnd vdd FILL
XFILL_4_DFFPOSX1_692 gnd vdd FILL
XFILL_4_DFFPOSX1_681 gnd vdd FILL
XFILL_0_CLKBUF1_7 gnd vdd FILL
XFILL_4_CLKBUF1_6 gnd vdd FILL
XFILL_3_XNOR2X1_103 gnd vdd FILL
XFILL_0_BUFX4_123 gnd vdd FILL
XFILL_0_BUFX4_101 gnd vdd FILL
XFILL_0_BUFX4_112 gnd vdd FILL
XFILL_1_BUFX2_582 gnd vdd FILL
XFILL_0_BUFX4_156 gnd vdd FILL
XFILL_1_OAI21X1_1515 gnd vdd FILL
XFILL_0_BUFX4_145 gnd vdd FILL
XOAI21X1_1328 BUFX4_6/A BUFX4_344/Y BUFX2_168/A gnd OAI21X1_1330/C vdd OAI21X1
XFILL_0_BUFX4_134 gnd vdd FILL
XFILL_0_BUFX4_167 gnd vdd FILL
XOAI21X1_1306 INVX2_106/Y INVX2_76/Y INVX2_77/Y gnd OAI21X1_1307/C vdd OAI21X1
XFILL_1_OAI21X1_1504 gnd vdd FILL
XFILL_1_BUFX2_593 gnd vdd FILL
XOAI21X1_1317 NOR3X1_16/C INVX8_3/Y INVX2_79/Y gnd OAI21X1_1318/C vdd OAI21X1
XFILL_3_DFFPOSX1_282 gnd vdd FILL
XFILL_3_DFFPOSX1_271 gnd vdd FILL
XFILL_0_BUFX4_178 gnd vdd FILL
XFILL_1_BUFX2_23 gnd vdd FILL
XOAI21X1_1339 BUFX4_99/Y BUFX4_342/Y BUFX2_172/A gnd OAI21X1_1341/C vdd OAI21X1
XFILL_1_OAI21X1_1526 gnd vdd FILL
XFILL_1_BUFX2_45 gnd vdd FILL
XDFFPOSX1_918 BUFX2_170/A CLKBUF1_68/Y OAI21X1_1335/Y gnd vdd DFFPOSX1
XDFFPOSX1_929 BUFX2_182/A CLKBUF1_36/Y OAI21X1_1367/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1537 gnd vdd FILL
XFILL_1_BUFX2_34 gnd vdd FILL
XFILL_0_BUFX4_189 gnd vdd FILL
XFILL_3_DFFPOSX1_260 gnd vdd FILL
XFILL_1_OAI21X1_1548 gnd vdd FILL
XDFFPOSX1_907 BUFX2_158/A CLKBUF1_53/Y OAI21X1_1305/Y gnd vdd DFFPOSX1
XFILL_1_BUFX2_67 gnd vdd FILL
XFILL_0_OAI21X1_306 gnd vdd FILL
XFILL_1_OAI21X1_1559 gnd vdd FILL
XFILL_0_OAI21X1_328 gnd vdd FILL
XFILL_0_OAI21X1_317 gnd vdd FILL
XFILL_1_BUFX2_78 gnd vdd FILL
XFILL_3_DFFPOSX1_293 gnd vdd FILL
XFILL_1_BUFX2_89 gnd vdd FILL
XFILL_6_DFFPOSX1_720 gnd vdd FILL
XFILL_0_OAI21X1_339 gnd vdd FILL
XFILL_6_DFFPOSX1_731 gnd vdd FILL
XFILL_5_DFFPOSX1_1 gnd vdd FILL
XFILL_37_8_1 gnd vdd FILL
XFILL_0_NAND2X1_301 gnd vdd FILL
XFILL_36_3_0 gnd vdd FILL
XFILL_0_OAI21X1_1105 gnd vdd FILL
XFILL_0_NAND2X1_334 gnd vdd FILL
XFILL_0_NAND2X1_323 gnd vdd FILL
XFILL_0_NAND2X1_312 gnd vdd FILL
XFILL_0_NAND2X1_367 gnd vdd FILL
XFILL_0_NAND2X1_356 gnd vdd FILL
XFILL_0_OAI21X1_1116 gnd vdd FILL
XFILL_0_OAI21X1_1127 gnd vdd FILL
XFILL_1_NAND2X1_516 gnd vdd FILL
XFILL_1_NAND2X1_527 gnd vdd FILL
XFILL_0_NAND2X1_345 gnd vdd FILL
XFILL_1_NOR2X1_3 gnd vdd FILL
XFILL_1_NAND2X1_538 gnd vdd FILL
XFILL_0_DFFPOSX1_706 gnd vdd FILL
XFILL_0_OAI21X1_1138 gnd vdd FILL
XFILL_0_NAND2X1_378 gnd vdd FILL
XFILL_0_OAI21X1_1149 gnd vdd FILL
XFILL_0_DFFPOSX1_728 gnd vdd FILL
XFILL_0_NAND2X1_389 gnd vdd FILL
XFILL_0_DFFPOSX1_717 gnd vdd FILL
XFILL_0_DFFPOSX1_739 gnd vdd FILL
XFILL_5_DFFPOSX1_310 gnd vdd FILL
XFILL_5_DFFPOSX1_321 gnd vdd FILL
XFILL_20_7_1 gnd vdd FILL
XFILL_5_DFFPOSX1_343 gnd vdd FILL
XFILL_5_DFFPOSX1_354 gnd vdd FILL
XFILL_5_DFFPOSX1_332 gnd vdd FILL
XFILL_5_DFFPOSX1_365 gnd vdd FILL
XFILL_5_DFFPOSX1_376 gnd vdd FILL
XFILL_0_MUX2X1_1 gnd vdd FILL
XFILL_5_DFFPOSX1_387 gnd vdd FILL
XFILL_1_NAND2X1_14 gnd vdd FILL
XFILL_5_DFFPOSX1_398 gnd vdd FILL
XFILL_1_NAND2X1_25 gnd vdd FILL
XINVX4_26 bundleStartMajId_i[5] gnd INVX4_26/Y vdd INVX4
XFILL_1_NAND2X1_47 gnd vdd FILL
XFILL_1_NAND2X1_36 gnd vdd FILL
XINVX4_15 bundleStartMajId_i[30] gnd INVX4_15/Y vdd INVX4
XFILL_1_NAND2X1_69 gnd vdd FILL
XINVX4_37 bundleAddress_i[38] gnd INVX4_37/Y vdd INVX4
XINVX4_48 INVX4_48/A gnd INVX4_48/Y vdd INVX4
XFILL_0_OAI21X1_840 gnd vdd FILL
XFILL_0_OAI21X1_873 gnd vdd FILL
XFILL_0_OAI21X1_884 gnd vdd FILL
XFILL_0_OAI21X1_862 gnd vdd FILL
XFILL_0_OAI21X1_851 gnd vdd FILL
XFILL_0_OAI21X1_895 gnd vdd FILL
XFILL_2_DFFPOSX1_21 gnd vdd FILL
XFILL_2_DFFPOSX1_10 gnd vdd FILL
XBUFX2_909 BUFX2_909/A gnd tid3_o[51] vdd BUFX2
XFILL_2_DFFPOSX1_32 gnd vdd FILL
XFILL_2_DFFPOSX1_43 gnd vdd FILL
XFILL_28_8_1 gnd vdd FILL
XFILL_2_DFFPOSX1_54 gnd vdd FILL
XFILL_3_8_1 gnd vdd FILL
XFILL_2_DFFPOSX1_76 gnd vdd FILL
XFILL_27_3_0 gnd vdd FILL
XFILL_2_DFFPOSX1_87 gnd vdd FILL
XFILL_2_DFFPOSX1_65 gnd vdd FILL
XFILL_2_3_0 gnd vdd FILL
XFILL_2_DFFPOSX1_98 gnd vdd FILL
XFILL_0_OAI21X1_1661 gnd vdd FILL
XFILL_0_OAI21X1_1650 gnd vdd FILL
XFILL_0_OAI21X1_1694 gnd vdd FILL
XFILL_0_OAI21X1_1683 gnd vdd FILL
XFILL_0_OAI21X1_1672 gnd vdd FILL
XFILL_11_7_1 gnd vdd FILL
XFILL_0_BUFX4_3 gnd vdd FILL
XFILL_10_2_0 gnd vdd FILL
XFILL_0_BUFX2_605 gnd vdd FILL
XFILL_0_BUFX2_616 gnd vdd FILL
XFILL_0_BUFX2_638 gnd vdd FILL
XFILL_4_DFFPOSX1_1000 gnd vdd FILL
XFILL_0_BUFX2_627 gnd vdd FILL
XFILL_20_18_0 gnd vdd FILL
XFILL_4_DFFPOSX1_1011 gnd vdd FILL
XFILL_0_BUFX2_649 gnd vdd FILL
XFILL_4_DFFPOSX1_1022 gnd vdd FILL
XBUFX4_202 BUFX4_26/Y gnd BUFX4_202/Y vdd BUFX4
XBUFX4_235 BUFX4_25/Y gnd BUFX4_235/Y vdd BUFX4
XBUFX4_246 INVX8_5/Y gnd BUFX4_3/A vdd BUFX4
XBUFX4_224 BUFX4_22/Y gnd BUFX4_224/Y vdd BUFX4
XBUFX4_213 BUFX4_25/Y gnd BUFX4_213/Y vdd BUFX4
XFILL_19_8_1 gnd vdd FILL
XFILL_0_INVX2_101 gnd vdd FILL
XFILL_0_INVX2_134 gnd vdd FILL
XFILL_2_OAI21X1_1755 gnd vdd FILL
XBUFX4_279 INVX8_7/Y gnd BUFX4_67/A vdd BUFX4
XBUFX4_257 INVX8_5/Y gnd BUFX4_11/A vdd BUFX4
XFILL_18_3_0 gnd vdd FILL
XFILL_0_INVX2_112 gnd vdd FILL
XBUFX4_268 enable_i gnd BUFX4_268/Y vdd BUFX4
XFILL_0_INVX2_123 gnd vdd FILL
XFILL_0_INVX2_145 gnd vdd FILL
XFILL_0_INVX2_167 gnd vdd FILL
XFILL_0_INVX2_156 gnd vdd FILL
XFILL_0_INVX2_189 gnd vdd FILL
XFILL_0_INVX2_178 gnd vdd FILL
XFILL_0_INVX4_3 gnd vdd FILL
XFILL_18_4 gnd vdd FILL
XFILL_25_17_0 gnd vdd FILL
XFILL_1_BUFX2_390 gnd vdd FILL
XOAI21X1_1103 INVX1_182/Y BUFX4_238/Y NAND2X1_469/Y gnd OAI21X1_1103/Y vdd OAI21X1
XDFFPOSX1_704 BUFX2_342/A CLKBUF1_96/Y OAI21X1_957/Y gnd vdd DFFPOSX1
XOAI21X1_1114 OAI21X1_1114/A BUFX4_216/Y NAND2X1_478/Y gnd OAI21X1_1114/Y vdd OAI21X1
XOAI21X1_1125 INVX2_95/Y INVX2_96/A INVX2_65/Y gnd NAND2X1_490/A vdd OAI21X1
XOAI21X1_1147 XNOR2X1_64/Y BUFX4_229/Y NAND2X1_522/Y gnd OAI21X1_1147/Y vdd OAI21X1
XFILL_1_OAI21X1_1301 gnd vdd FILL
XFILL_1_OAI21X1_1323 gnd vdd FILL
XFILL_1_OAI21X1_1312 gnd vdd FILL
XOAI21X1_1136 OAI21X1_1136/A NOR2X1_138/B NAND2X1_506/Y gnd OAI21X1_1136/Y vdd OAI21X1
XDFFPOSX1_715 BUFX2_380/A CLKBUF1_102/Y OAI21X1_979/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_103 gnd vdd FILL
XDFFPOSX1_737 BUFX2_375/A CLKBUF1_64/Y OAI21X1_1023/Y gnd vdd DFFPOSX1
XDFFPOSX1_748 BUFX2_35/A CLKBUF1_31/Y OAI21X1_1040/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_902 gnd vdd FILL
XFILL_1_OAI21X1_1334 gnd vdd FILL
XFILL_1_OAI21X1_1345 gnd vdd FILL
XOAI21X1_1169 INVX1_194/Y OAI21X1_1169/B NAND2X1_550/Y gnd OAI21X1_1169/Y vdd OAI21X1
XFILL_1_DFFPOSX1_924 gnd vdd FILL
XOAI21X1_1158 OAI21X1_1158/A XNOR2X1_67/A NAND2X1_534/Y gnd OAI21X1_1158/Y vdd OAI21X1
XFILL_1_OAI21X1_1356 gnd vdd FILL
XDFFPOSX1_726 BUFX2_363/A CLKBUF1_81/Y OAI21X1_1001/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_913 gnd vdd FILL
XFILL_1_OAI21X1_307 gnd vdd FILL
XFILL_0_OAI21X1_125 gnd vdd FILL
XDFFPOSX1_759 BUFX2_8/A CLKBUF1_59/Y OAI21X1_1051/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_114 gnd vdd FILL
XFILL_1_DFFPOSX1_946 gnd vdd FILL
XFILL_1_OAI21X1_1389 gnd vdd FILL
XFILL_1_DFFPOSX1_935 gnd vdd FILL
XFILL_1_OAI21X1_1378 gnd vdd FILL
XFILL_1_OAI21X1_1367 gnd vdd FILL
XFILL_1_DFFPOSX1_957 gnd vdd FILL
XFILL_0_OAI21X1_136 gnd vdd FILL
XFILL_0_OAI21X1_158 gnd vdd FILL
XFILL_0_OAI21X1_169 gnd vdd FILL
XFILL_0_OAI21X1_147 gnd vdd FILL
XFILL_1_DFFPOSX1_968 gnd vdd FILL
XFILL_1_OAI21X1_329 gnd vdd FILL
XFILL_1_DFFPOSX1_979 gnd vdd FILL
XFILL_1_OAI21X1_318 gnd vdd FILL
XFILL_6_DFFPOSX1_572 gnd vdd FILL
XFILL_6_DFFPOSX1_583 gnd vdd FILL
XFILL_6_DFFPOSX1_594 gnd vdd FILL
XFILL_0_BUFX4_35 gnd vdd FILL
XFILL_0_BUFX4_24 gnd vdd FILL
XFILL_0_BUFX4_13 gnd vdd FILL
XFILL_0_NAND2X1_131 gnd vdd FILL
XFILL_0_BUFX4_57 gnd vdd FILL
XFILL_0_BUFX4_46 gnd vdd FILL
XFILL_1_NAND2X1_302 gnd vdd FILL
XFILL_0_NAND2X1_142 gnd vdd FILL
XFILL_0_NAND2X1_120 gnd vdd FILL
XFILL_0_18_0 gnd vdd FILL
XFILL_0_BUFX4_68 gnd vdd FILL
XFILL_1_NAND2X1_346 gnd vdd FILL
XFILL_1_NAND2X1_335 gnd vdd FILL
XFILL_0_DFFPOSX1_503 gnd vdd FILL
XFILL_0_DFFPOSX1_514 gnd vdd FILL
XFILL_0_BUFX4_79 gnd vdd FILL
XFILL_1_NAND2X1_324 gnd vdd FILL
XFILL_0_NAND2X1_175 gnd vdd FILL
XFILL_0_NAND2X1_186 gnd vdd FILL
XFILL_0_NAND2X1_164 gnd vdd FILL
XFILL_0_NAND2X1_153 gnd vdd FILL
XFILL_0_DFFPOSX1_547 gnd vdd FILL
XFILL_0_DFFPOSX1_525 gnd vdd FILL
XFILL_0_DFFPOSX1_536 gnd vdd FILL
XFILL_1_NAND2X1_379 gnd vdd FILL
XFILL_0_DFFPOSX1_558 gnd vdd FILL
XFILL_0_NAND2X1_197 gnd vdd FILL
XFILL_0_DFFPOSX1_569 gnd vdd FILL
XFILL_5_DFFPOSX1_151 gnd vdd FILL
XFILL_5_DFFPOSX1_162 gnd vdd FILL
XFILL_5_DFFPOSX1_140 gnd vdd FILL
XFILL_5_DFFPOSX1_195 gnd vdd FILL
XFILL_5_DFFPOSX1_173 gnd vdd FILL
XFILL_5_DFFPOSX1_184 gnd vdd FILL
XOAI21X1_1692 BUFX4_11/A BUFX4_332/Y BUFX2_729/A gnd OAI21X1_1693/C vdd OAI21X1
XOAI21X1_1681 BUFX4_178/Y INVX2_134/Y OAI21X1_1681/C gnd DFFPOSX1_53/D vdd OAI21X1
XOAI21X1_1670 BUFX4_98/Y BUFX4_376/Y BUFX2_717/A gnd OAI21X1_1671/C vdd OAI21X1
XFILL_0_OR2X2_16 gnd vdd FILL
XFILL_1_OAI21X1_830 gnd vdd FILL
XFILL_1_OAI21X1_852 gnd vdd FILL
XNAND3X1_13 BUFX4_240/Y NAND3X1_13/B NAND3X1_13/C gnd NAND3X1_13/Y vdd NAND3X1
XFILL_0_OAI21X1_681 gnd vdd FILL
XFILL_1_OAI21X1_841 gnd vdd FILL
XFILL_0_OAI21X1_692 gnd vdd FILL
XFILL_0_OAI21X1_670 gnd vdd FILL
XFILL_1_OAI21X1_863 gnd vdd FILL
XFILL_1_OAI21X1_896 gnd vdd FILL
XNAND3X1_46 bundleAddress_i[17] INVX2_111/A NOR2X1_160/Y gnd INVX2_102/A vdd NAND3X1
XNAND3X1_35 bundleStartMajId_i[7] INVX2_47/Y NOR3X1_9/Y gnd XNOR2X1_55/A vdd NAND3X1
XNAND3X1_57 INVX2_107/Y AND2X2_26/Y INVX1_210/Y gnd NOR2X1_203/B vdd NAND3X1
XNAND3X1_24 NOR2X1_76/Y NOR2X1_91/Y AND2X2_13/Y gnd NOR2X1_97/B vdd NAND3X1
XFILL_1_OAI21X1_874 gnd vdd FILL
XFILL_1_OAI21X1_885 gnd vdd FILL
XNAND3X1_68 BUFX4_286/Y OR2X2_21/Y NAND3X1_68/C gnd NAND3X1_68/Y vdd NAND3X1
XFILL_5_17_0 gnd vdd FILL
XFILL_3_DFFPOSX1_11 gnd vdd FILL
XBUFX2_728 BUFX2_728/A gnd pid3_o[9] vdd BUFX2
XFILL_3_DFFPOSX1_44 gnd vdd FILL
XNOR2X1_46 INVX4_23/Y INVX2_33/Y gnd INVX2_51/A vdd NOR2X1
XFILL_3_DFFPOSX1_22 gnd vdd FILL
XBUFX2_717 BUFX2_717/A gnd pid3_o[19] vdd BUFX2
XNOR2X1_35 INVX4_19/Y NOR3X1_2/C gnd NOR2X1_35/Y vdd NOR2X1
XFILL_3_DFFPOSX1_33 gnd vdd FILL
XFILL_2_DFFPOSX1_608 gnd vdd FILL
XFILL_2_DFFPOSX1_619 gnd vdd FILL
XBUFX2_706 BUFX2_706/A gnd pid2_o[0] vdd BUFX2
XNOR2X1_24 OR2X2_8/A INVX1_15/A gnd NOR2X1_24/Y vdd NOR2X1
XNOR2X1_13 OR2X2_2/Y INVX1_10/A gnd XNOR2X1_7/A vdd NOR2X1
XFILL_3_DFFPOSX1_77 gnd vdd FILL
XNOR2X1_57 INVX4_27/Y INVX1_5/Y gnd INVX4_28/A vdd NOR2X1
XFILL_3_DFFPOSX1_55 gnd vdd FILL
XBUFX2_739 BUFX2_739/A gnd pid3_o[27] vdd BUFX2
XNOR2X1_79 INVX2_26/Y NOR3X1_5/C gnd NOR2X1_79/Y vdd NOR2X1
XNOR2X1_68 NOR2X1_69/A OR2X2_6/A gnd NOR2X1_68/Y vdd NOR2X1
XFILL_3_DFFPOSX1_66 gnd vdd FILL
XFILL_3_DFFPOSX1_88 gnd vdd FILL
XFILL_3_DFFPOSX1_99 gnd vdd FILL
XFILL_0_OAI21X1_1480 gnd vdd FILL
XFILL_0_OAI21X1_1491 gnd vdd FILL
XINVX2_202 bundleTid_i[7] gnd INVX2_202/Y vdd INVX2
XFILL_0_BUFX2_402 gnd vdd FILL
XFILL_0_BUFX2_413 gnd vdd FILL
XFILL_1_DFFPOSX1_209 gnd vdd FILL
XFILL_0_BUFX2_446 gnd vdd FILL
XFILL_0_BUFX2_435 gnd vdd FILL
XFILL_0_BUFX2_457 gnd vdd FILL
XFILL_0_BUFX2_424 gnd vdd FILL
XFILL_0_BUFX2_468 gnd vdd FILL
XFILL_0_BUFX2_479 gnd vdd FILL
XFILL_14_14_1 gnd vdd FILL
XFILL_0_NAND2X1_22 gnd vdd FILL
XFILL_0_NAND2X1_11 gnd vdd FILL
XFILL_0_NAND2X1_55 gnd vdd FILL
XFILL_0_NAND2X1_33 gnd vdd FILL
XFILL_0_NAND2X1_44 gnd vdd FILL
XFILL_2_OAI21X1_1574 gnd vdd FILL
XNOR2X1_114 INVX4_19/Y NOR2X1_114/B gnd INVX4_31/A vdd NOR2X1
XNOR2X1_103 INVX4_2/Y INVX1_34/Y gnd NOR2X1_103/Y vdd NOR2X1
XFILL_34_6_1 gnd vdd FILL
XNOR2X1_125 NOR2X1_180/A INVX4_47/Y gnd INVX2_93/A vdd NOR2X1
XNOR2X1_147 bundleAddress_i[32] NOR2X1_148/B gnd NOR2X1_147/Y vdd NOR2X1
XNOR2X1_136 INVX2_69/Y INVX4_35/Y gnd INVX2_97/A vdd NOR2X1
XFILL_2_OAI21X1_1585 gnd vdd FILL
XFILL_0_NAND2X1_66 gnd vdd FILL
XFILL_0_NAND2X1_77 gnd vdd FILL
XFILL_0_NAND2X1_88 gnd vdd FILL
XNOR2X1_158 INVX2_78/Y INVX8_3/Y gnd NOR2X1_158/Y vdd NOR2X1
XFILL_33_1_0 gnd vdd FILL
XNOR2X1_169 INVX2_86/Y INVX1_196/A gnd INVX4_48/A vdd NOR2X1
XFILL_0_NAND2X1_99 gnd vdd FILL
XOAI21X1_609 BUFX4_2/A BUFX4_362/Y BUFX2_559/A gnd OAI21X1_611/C vdd OAI21X1
XFILL_16_1 gnd vdd FILL
XFILL_1_OAI21X1_1131 gnd vdd FILL
XFILL_1_OAI21X1_1120 gnd vdd FILL
XDFFPOSX1_512 INVX1_28/A CLKBUF1_88/Y OAI21X1_576/Y gnd vdd DFFPOSX1
XDFFPOSX1_501 BUFX2_530/A CLKBUF1_80/Y OAI21X1_548/Y gnd vdd DFFPOSX1
XDFFPOSX1_523 INVX1_29/A CLKBUF1_44/Y OAI21X1_604/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_710 gnd vdd FILL
XDFFPOSX1_545 BUFX2_579/A CLKBUF1_70/Y OAI21X1_654/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_721 gnd vdd FILL
XFILL_1_OAI21X1_1153 gnd vdd FILL
XDFFPOSX1_534 BUFX2_567/A CLKBUF1_100/Y OAI21X1_628/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_732 gnd vdd FILL
XFILL_1_OAI21X1_1164 gnd vdd FILL
XDFFPOSX1_556 BUFX2_647/A CLKBUF1_13/Y OAI21X1_683/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1142 gnd vdd FILL
XFILL_1_OAI21X1_126 gnd vdd FILL
XFILL_0_BUFX2_980 gnd vdd FILL
XFILL_1_OAI21X1_115 gnd vdd FILL
XFILL_1_DFFPOSX1_754 gnd vdd FILL
XFILL_1_DFFPOSX1_776 gnd vdd FILL
XFILL_0_BUFX2_991 gnd vdd FILL
XFILL_1_OAI21X1_1175 gnd vdd FILL
XFILL_1_OAI21X1_104 gnd vdd FILL
XDFFPOSX1_578 BUFX2_609/A CLKBUF1_1/Y OAI21X1_745/Y gnd vdd DFFPOSX1
XDFFPOSX1_567 BUFX2_596/A CLKBUF1_1/Y OAI21X1_715/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_743 gnd vdd FILL
XFILL_1_OAI21X1_1197 gnd vdd FILL
XDFFPOSX1_589 BUFX2_621/A CLKBUF1_80/Y OAI21X1_774/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1186 gnd vdd FILL
XFILL_1_DFFPOSX1_765 gnd vdd FILL
XFILL_1_OAI21X1_159 gnd vdd FILL
XFILL_1_OAI21X1_148 gnd vdd FILL
XNAND2X1_626 INVX2_105/A INVX1_221/A gnd XNOR2X1_93/A vdd NAND2X1
XFILL_1_DFFPOSX1_787 gnd vdd FILL
XNAND2X1_604 bundleAddress_i[36] bundleAddress_i[35] gnd INVX1_207/A vdd NAND2X1
XFILL_19_13_1 gnd vdd FILL
XNAND2X1_615 bundleAddress_i[20] NOR3X1_17/Y gnd NAND2X1_616/A vdd NAND2X1
XFILL_1_DFFPOSX1_798 gnd vdd FILL
XFILL_1_OAI21X1_137 gnd vdd FILL
XNAND2X1_659 BUFX2_680/A BUFX4_380/Y gnd NAND2X1_659/Y vdd NAND2X1
XNAND2X1_648 BUFX2_389/A BUFX4_328/Y gnd NAND2X1_648/Y vdd NAND2X1
XINVX1_27 OR2X2_6/A gnd INVX1_27/Y vdd INVX1
XNAND2X1_637 bundleAddress_i[29] INVX1_208/Y gnd NAND2X1_637/Y vdd NAND2X1
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XINVX1_49 INVX1_49/A gnd INVX1_49/Y vdd INVX1
XFILL_6_DFFPOSX1_380 gnd vdd FILL
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XFILL_32_15_1 gnd vdd FILL
XNAND2X1_90 BUFX2_403/A BUFX4_351/Y gnd NAND2X1_90/Y vdd NAND2X1
XFILL_1_NAND2X1_110 gnd vdd FILL
XFILL_25_6_1 gnd vdd FILL
XFILL_1_NAND2X1_121 gnd vdd FILL
XFILL_0_6_1 gnd vdd FILL
XFILL_0_XNOR2X1_101 gnd vdd FILL
XFILL_0_DFFPOSX1_322 gnd vdd FILL
XFILL_0_DFFPOSX1_333 gnd vdd FILL
XFILL_0_DFFPOSX1_311 gnd vdd FILL
XFILL_24_1_0 gnd vdd FILL
XFILL_0_DFFPOSX1_300 gnd vdd FILL
XFILL_1_NAND2X1_143 gnd vdd FILL
XFILL_1_NAND2X1_165 gnd vdd FILL
XFILL_1_NAND2X1_187 gnd vdd FILL
XFILL_0_DFFPOSX1_366 gnd vdd FILL
XFILL_0_DFFPOSX1_355 gnd vdd FILL
XFILL_1_NAND2X1_198 gnd vdd FILL
XFILL_0_DFFPOSX1_344 gnd vdd FILL
XFILL_0_DFFPOSX1_399 gnd vdd FILL
XFILL_0_DFFPOSX1_388 gnd vdd FILL
XFILL_0_DFFPOSX1_377 gnd vdd FILL
XFILL_3_DFFPOSX1_804 gnd vdd FILL
XFILL_3_DFFPOSX1_815 gnd vdd FILL
XFILL_3_DFFPOSX1_837 gnd vdd FILL
XFILL_3_DFFPOSX1_848 gnd vdd FILL
XFILL_3_DFFPOSX1_826 gnd vdd FILL
XFILL_3_DFFPOSX1_859 gnd vdd FILL
XFILL_37_14_1 gnd vdd FILL
XFILL_1_NOR2X1_232 gnd vdd FILL
XFILL_1_NOR2X1_221 gnd vdd FILL
XFILL_8_7_1 gnd vdd FILL
XFILL_1_OAI21X1_671 gnd vdd FILL
XFILL_7_2_0 gnd vdd FILL
XFILL_1_OAI21X1_660 gnd vdd FILL
XFILL_1_OAI21X1_693 gnd vdd FILL
XFILL_1_OAI21X1_682 gnd vdd FILL
XFILL_31_10_0 gnd vdd FILL
XBUFX2_503 BUFX2_503/A gnd majID2_o[13] vdd BUFX2
XFILL_4_DFFPOSX1_12 gnd vdd FILL
XFILL_2_DFFPOSX1_416 gnd vdd FILL
XFILL_2_DFFPOSX1_405 gnd vdd FILL
XBUFX2_514 BUFX2_514/A gnd majID2_o[3] vdd BUFX2
XFILL_2_DFFPOSX1_427 gnd vdd FILL
XFILL_4_DFFPOSX1_23 gnd vdd FILL
XBUFX2_536 BUFX2_536/A gnd majID3_o[41] vdd BUFX2
XBUFX2_525 BUFX2_525/A gnd majID3_o[51] vdd BUFX2
XFILL_2_DFFPOSX1_438 gnd vdd FILL
XBUFX2_558 BUFX2_558/A gnd majID3_o[21] vdd BUFX2
XFILL_4_DFFPOSX1_45 gnd vdd FILL
XFILL_4_DFFPOSX1_56 gnd vdd FILL
XBUFX2_569 BUFX2_569/A gnd majID3_o[11] vdd BUFX2
XBUFX2_547 NOR2X1_73/A gnd majID3_o[31] vdd BUFX2
XFILL_16_6_1 gnd vdd FILL
XFILL_4_DFFPOSX1_34 gnd vdd FILL
XFILL_2_DFFPOSX1_449 gnd vdd FILL
XFILL_4_DFFPOSX1_78 gnd vdd FILL
XFILL_4_DFFPOSX1_89 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XFILL_4_DFFPOSX1_67 gnd vdd FILL
XFILL_5_DFFPOSX1_909 gnd vdd FILL
XDFFPOSX1_1030 BUFX2_668/A CLKBUF1_99/Y OAI21X1_1607/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_232 gnd vdd FILL
XFILL_0_BUFX2_210 gnd vdd FILL
XFILL_0_BUFX2_221 gnd vdd FILL
XFILL_0_BUFX2_254 gnd vdd FILL
XFILL_0_BUFX2_265 gnd vdd FILL
XFILL_0_BUFX2_243 gnd vdd FILL
XFILL_0_BUFX2_298 gnd vdd FILL
XFILL_0_BUFX2_276 gnd vdd FILL
XFILL_0_BUFX2_287 gnd vdd FILL
XFILL_2_DFFPOSX1_950 gnd vdd FILL
XFILL_2_DFFPOSX1_961 gnd vdd FILL
XFILL_2_DFFPOSX1_983 gnd vdd FILL
XFILL_2_DFFPOSX1_994 gnd vdd FILL
XFILL_2_DFFPOSX1_972 gnd vdd FILL
XFILL_0_NAND3X1_6 gnd vdd FILL
XOAI21X1_428 INVX1_10/A OR2X2_5/A OR2X2_5/B gnd OAI21X1_428/Y vdd OAI21X1
XOAI21X1_439 OAI21X1_439/A BUFX4_214/Y OAI21X1_439/C gnd OAI21X1_439/Y vdd OAI21X1
XOAI21X1_406 INVX1_8/A NOR2X1_60/A OAI21X1_406/C gnd OAI21X1_407/A vdd OAI21X1
XOAI21X1_417 XNOR2X1_2/A INVX4_4/Y INVX4_5/Y gnd OAI21X1_418/C vdd OAI21X1
XFILL_3_XNOR2X1_41 gnd vdd FILL
XFILL_3_XNOR2X1_74 gnd vdd FILL
XDFFPOSX1_331 BUFX2_1002/A CLKBUF1_26/Y OAI21X1_279/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_63 gnd vdd FILL
XFILL_3_XNOR2X1_52 gnd vdd FILL
XDFFPOSX1_320 BUFX2_990/A CLKBUF1_71/Y OAI21X1_257/Y gnd vdd DFFPOSX1
XDFFPOSX1_342 BUFX2_1015/A CLKBUF1_25/Y OAI21X1_301/Y gnd vdd DFFPOSX1
XDFFPOSX1_353 BUFX2_1027/A CLKBUF1_22/Y OAI21X1_323/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_551 gnd vdd FILL
XFILL_3_XNOR2X1_85 gnd vdd FILL
XFILL_3_XNOR2X1_96 gnd vdd FILL
XFILL_1_DFFPOSX1_540 gnd vdd FILL
XDFFPOSX1_364 BUFX2_455/A CLKBUF1_6/Y OAI21X1_336/Y gnd vdd DFFPOSX1
XNAND2X1_401 BUFX2_318/A BUFX4_184/Y gnd OAI21X1_907/C vdd NAND2X1
XDFFPOSX1_375 BUFX2_404/A CLKBUF1_1/Y OAI21X1_347/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_584 gnd vdd FILL
XDFFPOSX1_397 BUFX2_429/A CLKBUF1_84/Y OAI21X1_369/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_573 gnd vdd FILL
XDFFPOSX1_386 BUFX2_417/A CLKBUF1_63/Y OAI21X1_358/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_562 gnd vdd FILL
XNAND2X1_412 BUFX2_3/A BUFX4_328/Y gnd NAND2X1_412/Y vdd NAND2X1
XNAND2X1_434 BUFX2_27/A BUFX4_381/Y gnd NAND2X1_434/Y vdd NAND2X1
XFILL_1_DFFPOSX1_595 gnd vdd FILL
XNAND2X1_445 BUFX2_39/A BUFX4_344/Y gnd NAND2X1_445/Y vdd NAND2X1
XFILL_2_OAI21X1_116 gnd vdd FILL
XNAND2X1_423 BUFX2_15/A BUFX4_354/Y gnd NAND2X1_423/Y vdd NAND2X1
XNAND2X1_478 BUFX2_126/A BUFX4_216/Y gnd NAND2X1_478/Y vdd NAND2X1
XFILL_2_OAI21X1_149 gnd vdd FILL
XNAND2X1_467 BUFX2_66/A BUFX4_230/Y gnd NAND2X1_467/Y vdd NAND2X1
XNAND2X1_456 BUFX2_51/A BUFX4_374/Y gnd NAND2X1_456/Y vdd NAND2X1
XNAND2X1_489 bundleAddress_i[50] NOR2X1_129/Y gnd NAND2X1_492/B vdd NAND2X1
XFILL_0_DFFPOSX1_130 gnd vdd FILL
XFILL_1_XNOR2X1_102 gnd vdd FILL
XFILL_0_DFFPOSX1_141 gnd vdd FILL
XFILL_1_BUFX2_912 gnd vdd FILL
XFILL_0_DFFPOSX1_163 gnd vdd FILL
XFILL_0_DFFPOSX1_152 gnd vdd FILL
XFILL_0_DFFPOSX1_174 gnd vdd FILL
XFILL_1_BUFX2_923 gnd vdd FILL
XFILL_0_DFFPOSX1_185 gnd vdd FILL
XFILL_1_BUFX2_934 gnd vdd FILL
XFILL_0_DFFPOSX1_196 gnd vdd FILL
XFILL_1_BUFX2_978 gnd vdd FILL
XOAI21X1_951 BUFX4_136/Y INVX1_130/Y OAI21X1_951/C gnd OAI21X1_951/Y vdd OAI21X1
XOAI21X1_940 BUFX4_105/Y NAND2X1_7/B BUFX2_333/A gnd OAI21X1_941/C vdd OAI21X1
XFILL_3_DFFPOSX1_601 gnd vdd FILL
XFILL_3_DFFPOSX1_612 gnd vdd FILL
XFILL_1_BUFX2_967 gnd vdd FILL
XOAI21X1_984 BUFX4_137/Y BUFX4_34/Y BUFX2_385/A gnd OAI21X1_985/C vdd OAI21X1
XFILL_3_DFFPOSX1_645 gnd vdd FILL
XFILL_3_DFFPOSX1_634 gnd vdd FILL
XFILL_3_DFFPOSX1_656 gnd vdd FILL
XOAI21X1_962 BUFX4_7/A BUFX4_315/Y BUFX2_345/A gnd OAI21X1_963/C vdd OAI21X1
XFILL_3_DFFPOSX1_623 gnd vdd FILL
XOAI21X1_973 BUFX4_295/Y INVX1_141/Y OAI21X1_973/C gnd OAI21X1_973/Y vdd OAI21X1
XFILL_3_DFFPOSX1_678 gnd vdd FILL
XFILL_3_DFFPOSX1_667 gnd vdd FILL
XFILL_3_DFFPOSX1_689 gnd vdd FILL
XOAI21X1_995 BUFX4_300/Y INVX1_152/Y OAI21X1_995/C gnd OAI21X1_995/Y vdd OAI21X1
XFILL_2_OAI21X1_650 gnd vdd FILL
XFILL_1_OAI21X1_490 gnd vdd FILL
XINVX2_81 bundleAddress_i[18] gnd INVX2_81/Y vdd INVX2
XINVX2_70 bundleAddress_i[41] gnd INVX2_70/Y vdd INVX2
XINVX2_92 bundleAddress_i[1] gnd INVX2_92/Y vdd INVX2
XFILL_0_NAND2X1_708 gnd vdd FILL
XFILL_2_DFFPOSX1_202 gnd vdd FILL
XFILL_2_DFFPOSX1_213 gnd vdd FILL
XBUFX2_300 BUFX2_300/A gnd instr2_o[16] vdd BUFX2
XBUFX2_311 BUFX2_311/A gnd instr2_o[6] vdd BUFX2
XBUFX2_322 BUFX2_322/A gnd instr2_o[24] vdd BUFX2
XFILL_0_NAND2X1_719 gnd vdd FILL
XFILL_2_DFFPOSX1_246 gnd vdd FILL
XFILL_2_DFFPOSX1_235 gnd vdd FILL
XBUFX2_333 BUFX2_333/A gnd instr3_o[15] vdd BUFX2
XBUFX2_344 BUFX2_344/A gnd instr3_o[5] vdd BUFX2
XFILL_2_DFFPOSX1_224 gnd vdd FILL
XFILL_5_DFFPOSX1_13 gnd vdd FILL
XBUFX2_355 BUFX2_355/A gnd instr3_o[23] vdd BUFX2
XFILL_5_DFFPOSX1_46 gnd vdd FILL
XBUFX2_366 BUFX2_366/A gnd instr4_o[14] vdd BUFX2
XFILL_5_DFFPOSX1_24 gnd vdd FILL
XFILL_2_DFFPOSX1_279 gnd vdd FILL
XFILL_2_DFFPOSX1_268 gnd vdd FILL
XBUFX2_377 BUFX2_377/A gnd instr4_o[4] vdd BUFX2
XFILL_2_DFFPOSX1_257 gnd vdd FILL
XFILL_5_DFFPOSX1_35 gnd vdd FILL
XFILL_5_DFFPOSX1_68 gnd vdd FILL
XBUFX2_388 BUFX2_388/A gnd instr4_o[22] vdd BUFX2
XFILL_5_DFFPOSX1_57 gnd vdd FILL
XFILL_5_DFFPOSX1_79 gnd vdd FILL
XFILL_1_NOR3X1_16 gnd vdd FILL
XBUFX2_399 BUFX2_399/A gnd majID1_o[49] vdd BUFX2
XOAI21X1_11 INVX2_149/Y BUFX4_222/Y OAI21X1_11/C gnd OAI21X1_11/Y vdd OAI21X1
XOAI21X1_22 INVX2_160/Y BUFX4_218/Y OAI21X1_22/C gnd OAI21X1_22/Y vdd OAI21X1
XOAI21X1_33 INVX2_171/Y BUFX4_229/Y OAI21X1_33/C gnd OAI21X1_33/Y vdd OAI21X1
XOAI21X1_44 INVX2_182/Y BUFX4_229/Y OAI21X1_44/C gnd OAI21X1_44/Y vdd OAI21X1
XFILL_31_4_1 gnd vdd FILL
XFILL_5_DFFPOSX1_728 gnd vdd FILL
XFILL_5_DFFPOSX1_706 gnd vdd FILL
XFILL_5_DFFPOSX1_717 gnd vdd FILL
XOAI21X1_55 INVX2_193/Y BUFX4_207/Y OAI21X1_55/C gnd OAI21X1_55/Y vdd OAI21X1
XFILL_1_BUFX4_282 gnd vdd FILL
XFILL_1_BUFX4_260 gnd vdd FILL
XFILL_1_BUFX4_271 gnd vdd FILL
XOAI21X1_66 INVX2_2/Y BUFX4_190/Y OAI21X1_66/C gnd OAI21X1_66/Y vdd OAI21X1
XOAI21X1_77 BUFX4_131/Y INVX2_148/Y OAI21X1_77/C gnd OAI21X1_77/Y vdd OAI21X1
XFILL_5_DFFPOSX1_739 gnd vdd FILL
XFILL_1_BUFX4_293 gnd vdd FILL
XOAI21X1_99 BUFX4_153/Y INVX2_159/Y OAI21X1_99/C gnd OAI21X1_99/Y vdd OAI21X1
XOAI21X1_88 BUFX4_7/A BUFX4_315/Y BUFX2_967/A gnd OAI21X1_89/C vdd OAI21X1
XFILL_22_15_0 gnd vdd FILL
XFILL_0_DFFPOSX1_20 gnd vdd FILL
XFILL_4_DFFPOSX1_318 gnd vdd FILL
XFILL_4_DFFPOSX1_307 gnd vdd FILL
XFILL_0_DFFPOSX1_53 gnd vdd FILL
XFILL_0_DFFPOSX1_31 gnd vdd FILL
XFILL_0_DFFPOSX1_42 gnd vdd FILL
XFILL_0_DFFPOSX1_75 gnd vdd FILL
XFILL_4_DFFPOSX1_329 gnd vdd FILL
XFILL_0_DFFPOSX1_64 gnd vdd FILL
XFILL_0_DFFPOSX1_86 gnd vdd FILL
XFILL_38_0_0 gnd vdd FILL
XFILL_0_DFFPOSX1_97 gnd vdd FILL
XFILL_2_DFFPOSX1_791 gnd vdd FILL
XFILL_2_DFFPOSX1_780 gnd vdd FILL
XFILL_22_4_1 gnd vdd FILL
XFILL_1_BUFX2_208 gnd vdd FILL
XFILL_6_DFFPOSX1_5 gnd vdd FILL
XFILL_1_BUFX2_219 gnd vdd FILL
XFILL_27_14_0 gnd vdd FILL
XOAI21X1_203 OAI21X1_9/A BUFX4_294/Y OAI21X1_203/C gnd OAI21X1_203/Y vdd OAI21X1
XOAI21X1_225 INVX2_158/Y BUFX4_293/Y OAI21X1_225/C gnd OAI21X1_225/Y vdd OAI21X1
XOAI21X1_247 INVX2_169/Y BUFX4_301/Y OAI21X1_247/C gnd OAI21X1_247/Y vdd OAI21X1
XOAI21X1_214 BUFX4_162/Y BUFX4_51/Y BUFX2_1030/A gnd OAI21X1_215/C vdd OAI21X1
XOAI21X1_236 BUFX4_129/Y BUFX4_67/Y BUFX2_979/A gnd OAI21X1_237/C vdd OAI21X1
XOAI21X1_269 INVX2_180/Y BUFX4_301/Y OAI21X1_269/C gnd OAI21X1_269/Y vdd OAI21X1
XOAI21X1_258 OR2X2_20/B BUFX4_59/A BUFX2_991/A gnd OAI21X1_259/C vdd OAI21X1
XAND2X2_25 NOR3X1_15/Y bundleAddress_i[0] gnd AND2X2_25/Y vdd AND2X2
XAND2X2_14 NOR2X1_19/Y NOR2X1_74/Y gnd AND2X2_14/Y vdd AND2X2
XDFFPOSX1_150 BUFX2_823/A CLKBUF1_102/Y OAI21X1_1824/Y gnd vdd DFFPOSX1
XDFFPOSX1_161 NAND2X1_5/A CLKBUF1_60/Y OAI21X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_172 BUFX2_903/A CLKBUF1_10/Y OAI21X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_194 BUFX2_865/A CLKBUF1_102/Y OAI21X1_38/Y gnd vdd DFFPOSX1
XDFFPOSX1_183 BUFX2_852/A CLKBUF1_98/Y OAI21X1_27/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_392 gnd vdd FILL
XFILL_1_DFFPOSX1_381 gnd vdd FILL
XFILL_0_NOR3X1_4 gnd vdd FILL
XNAND2X1_220 BUFX2_493/A BUFX4_204/Y gnd OAI21X1_461/C vdd NAND2X1
XFILL_1_DFFPOSX1_370 gnd vdd FILL
XNAND2X1_242 bundleStartMajId_i[15] INVX2_51/A gnd INVX2_45/A vdd NAND2X1
XNAND2X1_253 INVX2_47/Y INVX1_19/Y gnd OAI21X1_493/A vdd NAND2X1
XNAND2X1_231 NOR3X1_3/Y AND2X2_7/Y gnd NOR3X1_9/B vdd NAND2X1
XNAND2X1_264 BUFX2_517/A BUFX4_235/Y gnd NAND2X1_265/A vdd NAND2X1
XNAND2X1_286 OR2X2_7/A OAI21X1_582/Y gnd OAI21X1_584/A vdd NAND2X1
XNAND2X1_275 INVX4_30/A NOR2X1_62/Y gnd OR2X2_10/B vdd NAND2X1
XFILL_5_5_1 gnd vdd FILL
XFILL_4_DFFPOSX1_830 gnd vdd FILL
XFILL_4_DFFPOSX1_874 gnd vdd FILL
XFILL_4_DFFPOSX1_841 gnd vdd FILL
XFILL_29_0_0 gnd vdd FILL
XFILL_4_DFFPOSX1_852 gnd vdd FILL
XNAND2X1_297 NOR2X1_96/B OAI21X1_610/A gnd OAI21X1_608/A vdd NAND2X1
XFILL_4_0_0 gnd vdd FILL
XFILL_4_DFFPOSX1_863 gnd vdd FILL
XFILL_4_DFFPOSX1_885 gnd vdd FILL
XFILL_4_DFFPOSX1_896 gnd vdd FILL
XFILL_2_15_0 gnd vdd FILL
XFILL_0_OAI21X1_3 gnd vdd FILL
XFILL_13_4_1 gnd vdd FILL
XFILL_2_XNOR2X1_103 gnd vdd FILL
XFILL_1_BUFX2_720 gnd vdd FILL
XFILL_0_BUFX2_90 gnd vdd FILL
XFILL_1_BUFX2_731 gnd vdd FILL
XFILL_1_BUFX2_764 gnd vdd FILL
XFILL_0_BUFX4_316 gnd vdd FILL
XFILL_0_BUFX4_305 gnd vdd FILL
XFILL_1_NOR2X1_82 gnd vdd FILL
XFILL_1_NOR2X1_60 gnd vdd FILL
XFILL_1_BUFX2_775 gnd vdd FILL
XFILL_1_BUFX2_786 gnd vdd FILL
XFILL_0_BUFX4_349 gnd vdd FILL
XFILL_0_BUFX4_327 gnd vdd FILL
XFILL_3_DFFPOSX1_431 gnd vdd FILL
XFILL_3_DFFPOSX1_420 gnd vdd FILL
XFILL_0_BUFX4_338 gnd vdd FILL
XOAI21X1_781 BUFX4_161/Y BUFX4_82/Y BUFX2_623/A gnd OAI21X1_782/C vdd OAI21X1
XOAI21X1_770 OR2X2_15/A NOR2X1_42/A INVX4_19/Y gnd OAI21X1_770/Y vdd OAI21X1
XFILL_1_OAI21X1_1719 gnd vdd FILL
XOAI21X1_792 AND2X2_22/Y OAI21X1_792/B OAI21X1_792/C gnd OAI21X1_792/Y vdd OAI21X1
XFILL_3_DFFPOSX1_442 gnd vdd FILL
XFILL_3_DFFPOSX1_453 gnd vdd FILL
XFILL_3_DFFPOSX1_464 gnd vdd FILL
XFILL_1_OAI21X1_1708 gnd vdd FILL
XFILL_3_DFFPOSX1_486 gnd vdd FILL
XFILL_3_DFFPOSX1_497 gnd vdd FILL
XFILL_3_DFFPOSX1_475 gnd vdd FILL
XFILL_0_BUFX2_1009 gnd vdd FILL
XFILL_6_DFFPOSX1_902 gnd vdd FILL
XFILL_6_DFFPOSX1_913 gnd vdd FILL
XFILL_7_14_0 gnd vdd FILL
XFILL_0_NAND2X1_516 gnd vdd FILL
XFILL_0_NAND2X1_505 gnd vdd FILL
XBUFX2_141 BUFX2_141/A gnd addr3_o[61] vdd BUFX2
XBUFX2_152 BUFX2_152/A gnd addr3_o[60] vdd BUFX2
XFILL_0_NAND2X1_527 gnd vdd FILL
XBUFX2_130 BUFX2_130/A gnd addr3_o[62] vdd BUFX2
XFILL_0_NAND2X1_549 gnd vdd FILL
XFILL_0_NAND2X1_538 gnd vdd FILL
XFILL_11_12_1 gnd vdd FILL
XFILL_2_XNOR2X1_82 gnd vdd FILL
XFILL_1_NAND2X1_709 gnd vdd FILL
XFILL_2_XNOR2X1_71 gnd vdd FILL
XFILL_0_OAI21X1_1309 gnd vdd FILL
XFILL_2_XNOR2X1_60 gnd vdd FILL
XBUFX2_196 BUFX2_196/A gnd addr4_o[52] vdd BUFX2
XBUFX2_163 BUFX2_163/A gnd addr3_o[59] vdd BUFX2
XBUFX2_185 BUFX2_185/A gnd addr3_o[57] vdd BUFX2
XBUFX2_174 BUFX2_174/A gnd addr3_o[58] vdd BUFX2
XFILL_2_XNOR2X1_93 gnd vdd FILL
XFILL_1_NAND2X1_4 gnd vdd FILL
XFILL_5_DFFPOSX1_503 gnd vdd FILL
XFILL_5_DFFPOSX1_525 gnd vdd FILL
XFILL_5_DFFPOSX1_536 gnd vdd FILL
XFILL_5_DFFPOSX1_514 gnd vdd FILL
XFILL_5_DFFPOSX1_547 gnd vdd FILL
XFILL_5_DFFPOSX1_569 gnd vdd FILL
XFILL_5_DFFPOSX1_558 gnd vdd FILL
XBUFX2_1011 BUFX2_1011/A gnd tid4_o[16] vdd BUFX2
XBUFX2_1000 BUFX2_1000/A gnd tid4_o[26] vdd BUFX2
XBUFX2_1022 BUFX2_1022/A gnd tid4_o[6] vdd BUFX2
XCLKBUF1_12 BUFX4_85/Y gnd CLKBUF1_12/Y vdd CLKBUF1
XCLKBUF1_23 BUFX4_91/Y gnd CLKBUF1_23/Y vdd CLKBUF1
XFILL_1_AOI21X1_9 gnd vdd FILL
XFILL_1_DFFPOSX1_21 gnd vdd FILL
XFILL_4_DFFPOSX1_104 gnd vdd FILL
XFILL_1_DFFPOSX1_32 gnd vdd FILL
XFILL_4_DFFPOSX1_126 gnd vdd FILL
XFILL_4_DFFPOSX1_115 gnd vdd FILL
XCLKBUF1_45 BUFX4_83/Y gnd CLKBUF1_45/Y vdd CLKBUF1
XFILL_16_11_1 gnd vdd FILL
XCLKBUF1_34 BUFX4_88/Y gnd CLKBUF1_34/Y vdd CLKBUF1
XCLKBUF1_56 BUFX4_90/Y gnd CLKBUF1_56/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_10 gnd vdd FILL
XFILL_1_DFFPOSX1_43 gnd vdd FILL
XFILL_4_DFFPOSX1_137 gnd vdd FILL
XFILL_4_DFFPOSX1_148 gnd vdd FILL
XCLKBUF1_67 BUFX4_87/Y gnd CLKBUF1_67/Y vdd CLKBUF1
XCLKBUF1_89 BUFX4_92/Y gnd CLKBUF1_89/Y vdd CLKBUF1
XCLKBUF1_78 BUFX4_83/Y gnd CLKBUF1_78/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_54 gnd vdd FILL
XFILL_1_DFFPOSX1_65 gnd vdd FILL
XFILL_4_DFFPOSX1_159 gnd vdd FILL
XFILL_1_DFFPOSX1_76 gnd vdd FILL
XFILL_1_DFFPOSX1_87 gnd vdd FILL
XFILL_1_DFFPOSX1_98 gnd vdd FILL
XFILL_0_OAI21X1_1810 gnd vdd FILL
XFILL_0_OAI21X1_1821 gnd vdd FILL
XFILL_0_BUFX2_809 gnd vdd FILL
XINVX1_119 bundle_i[85] gnd INVX1_119/Y vdd INVX1
XINVX1_108 bundle_i[32] gnd INVX1_108/Y vdd INVX1
XFILL_3_XNOR2X1_7 gnd vdd FILL
XFILL_2_AOI21X1_60 gnd vdd FILL
XFILL_34_12_1 gnd vdd FILL
XFILL_0_INVX2_18 gnd vdd FILL
XFILL_0_INVX2_29 gnd vdd FILL
XFILL_4_DFFPOSX1_660 gnd vdd FILL
XFILL_4_DFFPOSX1_671 gnd vdd FILL
XFILL_4_DFFPOSX1_682 gnd vdd FILL
XFILL_4_DFFPOSX1_693 gnd vdd FILL
XFILL_0_CLKBUF1_8 gnd vdd FILL
XFILL_4_CLKBUF1_7 gnd vdd FILL
XFILL_3_XNOR2X1_104 gnd vdd FILL
XFILL_1_BUFX2_572 gnd vdd FILL
XFILL_0_BUFX4_113 gnd vdd FILL
XFILL_0_BUFX4_102 gnd vdd FILL
XFILL_1_BUFX2_561 gnd vdd FILL
XFILL_0_BUFX4_124 gnd vdd FILL
XFILL_0_BUFX4_146 gnd vdd FILL
XOAI21X1_1329 NOR2X1_203/B NOR2X1_204/A BUFX4_310/Y gnd OAI21X1_1330/A vdd OAI21X1
XFILL_0_BUFX4_157 gnd vdd FILL
XFILL_0_BUFX4_135 gnd vdd FILL
XOAI21X1_1307 INVX1_208/A INVX2_106/Y OAI21X1_1307/C gnd OAI21X1_1309/A vdd OAI21X1
XFILL_1_OAI21X1_1505 gnd vdd FILL
XFILL_1_BUFX2_583 gnd vdd FILL
XOAI21X1_1318 NOR3X1_16/B NOR3X1_16/C OAI21X1_1318/C gnd OAI21X1_1319/A vdd OAI21X1
XFILL_1_BUFX2_24 gnd vdd FILL
XFILL_1_BUFX2_13 gnd vdd FILL
XFILL_3_DFFPOSX1_261 gnd vdd FILL
XFILL_3_DFFPOSX1_272 gnd vdd FILL
XFILL_0_BUFX4_168 gnd vdd FILL
XDFFPOSX1_919 BUFX2_171/A CLKBUF1_21/Y OAI21X1_1338/Y gnd vdd DFFPOSX1
XFILL_0_BUFX4_179 gnd vdd FILL
XFILL_1_OAI21X1_1527 gnd vdd FILL
XFILL_1_OAI21X1_1516 gnd vdd FILL
XFILL_3_DFFPOSX1_250 gnd vdd FILL
XFILL_1_OAI21X1_1538 gnd vdd FILL
XFILL_1_OAI21X1_1549 gnd vdd FILL
XDFFPOSX1_908 BUFX2_159/A CLKBUF1_62/Y OAI21X1_1309/Y gnd vdd DFFPOSX1
XFILL_1_BUFX2_68 gnd vdd FILL
XFILL_0_OAI21X1_307 gnd vdd FILL
XFILL_1_BUFX2_57 gnd vdd FILL
XFILL_3_DFFPOSX1_283 gnd vdd FILL
XFILL_3_DFFPOSX1_294 gnd vdd FILL
XFILL_0_OAI21X1_318 gnd vdd FILL
XFILL_0_OAI21X1_329 gnd vdd FILL
XFILL_6_DFFPOSX1_754 gnd vdd FILL
XFILL_4_1 gnd vdd FILL
XFILL_6_DFFPOSX1_776 gnd vdd FILL
XFILL_6_DFFPOSX1_787 gnd vdd FILL
XFILL_5_DFFPOSX1_2 gnd vdd FILL
XFILL_6_DFFPOSX1_765 gnd vdd FILL
XFILL_6_DFFPOSX1_798 gnd vdd FILL
XFILL_36_3_1 gnd vdd FILL
XFILL_0_NAND2X1_335 gnd vdd FILL
XFILL_0_NAND2X1_302 gnd vdd FILL
XFILL_0_NAND2X1_324 gnd vdd FILL
XFILL_0_NAND2X1_313 gnd vdd FILL
XFILL_0_OAI21X1_1106 gnd vdd FILL
XFILL_0_NAND2X1_346 gnd vdd FILL
XFILL_0_OAI21X1_1128 gnd vdd FILL
XFILL_0_OAI21X1_1117 gnd vdd FILL
XFILL_1_NAND2X1_528 gnd vdd FILL
XFILL_1_NAND2X1_539 gnd vdd FILL
XFILL_0_DFFPOSX1_707 gnd vdd FILL
XFILL_0_NAND2X1_357 gnd vdd FILL
XFILL_0_NAND2X1_368 gnd vdd FILL
XFILL_0_OAI21X1_1139 gnd vdd FILL
XFILL_0_DFFPOSX1_718 gnd vdd FILL
XFILL_0_DFFPOSX1_729 gnd vdd FILL
XFILL_0_NAND2X1_379 gnd vdd FILL
XFILL_1_DFFPOSX1_1030 gnd vdd FILL
XFILL_5_DFFPOSX1_311 gnd vdd FILL
XFILL_5_DFFPOSX1_300 gnd vdd FILL
XFILL_5_DFFPOSX1_322 gnd vdd FILL
XFILL_5_DFFPOSX1_333 gnd vdd FILL
XFILL_5_DFFPOSX1_344 gnd vdd FILL
XFILL_0_MUX2X1_2 gnd vdd FILL
XFILL_5_DFFPOSX1_377 gnd vdd FILL
XFILL_5_DFFPOSX1_366 gnd vdd FILL
XFILL_5_DFFPOSX1_355 gnd vdd FILL
XFILL_5_DFFPOSX1_399 gnd vdd FILL
XFILL_5_DFFPOSX1_388 gnd vdd FILL
XOAI21X1_1830 BUFX4_361/Y INVX2_202/Y NAND2X1_771/Y gnd OAI21X1_1830/Y vdd OAI21X1
XINVX4_27 bundleStartMajId_i[2] gnd INVX4_27/Y vdd INVX4
XFILL_1_NAND2X1_26 gnd vdd FILL
XFILL_1_NAND2X1_48 gnd vdd FILL
XINVX4_16 bundleStartMajId_i[28] gnd OR2X2_8/B vdd INVX4
XINVX4_38 bundleAddress_i[34] gnd INVX4_38/Y vdd INVX4
XINVX4_49 INVX4_49/A gnd INVX4_49/Y vdd INVX4
XFILL_0_OAI21X1_830 gnd vdd FILL
XFILL_0_OAI21X1_841 gnd vdd FILL
XFILL_0_OAI21X1_852 gnd vdd FILL
XFILL_0_OAI21X1_874 gnd vdd FILL
XFILL_0_OAI21X1_863 gnd vdd FILL
XFILL_0_OAI21X1_896 gnd vdd FILL
XFILL_0_OAI21X1_885 gnd vdd FILL
XFILL_2_DFFPOSX1_11 gnd vdd FILL
XFILL_2_DFFPOSX1_44 gnd vdd FILL
XFILL_2_DFFPOSX1_22 gnd vdd FILL
XFILL_2_DFFPOSX1_55 gnd vdd FILL
XFILL_2_DFFPOSX1_33 gnd vdd FILL
XFILL_2_DFFPOSX1_77 gnd vdd FILL
XFILL_27_3_1 gnd vdd FILL
XFILL_2_DFFPOSX1_88 gnd vdd FILL
XFILL_2_3_1 gnd vdd FILL
XFILL_2_DFFPOSX1_66 gnd vdd FILL
XFILL_2_DFFPOSX1_99 gnd vdd FILL
XFILL_0_OAI21X1_1651 gnd vdd FILL
XFILL_0_OAI21X1_1640 gnd vdd FILL
XFILL_0_OAI21X1_1662 gnd vdd FILL
XFILL_0_OAI21X1_1695 gnd vdd FILL
XFILL_0_OAI21X1_1684 gnd vdd FILL
XFILL_0_OAI21X1_1673 gnd vdd FILL
XFILL_0_BUFX4_4 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XFILL_0_BUFX2_606 gnd vdd FILL
XFILL_0_BUFX2_639 gnd vdd FILL
XFILL_0_BUFX2_628 gnd vdd FILL
XFILL_20_18_1 gnd vdd FILL
XFILL_0_BUFX2_617 gnd vdd FILL
XFILL_4_DFFPOSX1_1012 gnd vdd FILL
XFILL_1_XNOR2X1_90 gnd vdd FILL
XFILL_4_DFFPOSX1_1001 gnd vdd FILL
XFILL_4_DFFPOSX1_1023 gnd vdd FILL
XBUFX4_203 BUFX4_23/Y gnd BUFX4_203/Y vdd BUFX4
XBUFX4_225 BUFX4_20/Y gnd BUFX4_225/Y vdd BUFX4
XBUFX4_236 BUFX4_22/Y gnd BUFX4_236/Y vdd BUFX4
XBUFX4_214 BUFX4_22/Y gnd BUFX4_214/Y vdd BUFX4
XFILL_2_OAI21X1_1723 gnd vdd FILL
XFILL_0_INVX2_124 gnd vdd FILL
XBUFX4_247 INVX8_5/Y gnd BUFX4_247/Y vdd BUFX4
XBUFX4_269 INVX8_7/Y gnd BUFX4_75/A vdd BUFX4
XFILL_0_INVX2_135 gnd vdd FILL
XFILL_0_INVX2_102 gnd vdd FILL
XFILL_18_3_1 gnd vdd FILL
XBUFX4_258 INVX8_5/Y gnd BUFX4_1/A vdd BUFX4
XFILL_4_DFFPOSX1_490 gnd vdd FILL
XFILL_0_INVX2_113 gnd vdd FILL
XFILL_0_INVX2_157 gnd vdd FILL
XFILL_2_OAI21X1_1778 gnd vdd FILL
XFILL_0_INVX2_146 gnd vdd FILL
XFILL_0_INVX2_168 gnd vdd FILL
XFILL_0_INVX2_179 gnd vdd FILL
XFILL_0_INVX4_4 gnd vdd FILL
XFILL_25_17_1 gnd vdd FILL
XFILL_1_BUFX2_380 gnd vdd FILL
XOAI21X1_1104 INVX4_32/Y INVX2_56/Y INVX2_57/Y gnd OAI21X1_1105/C vdd OAI21X1
XOAI21X1_1126 NAND2X1_490/Y BUFX4_235/Y NAND2X1_491/Y gnd OAI21X1_1126/Y vdd OAI21X1
XOAI21X1_1115 NAND2X1_476/Y NOR2X1_216/A INVX2_61/Y gnd NAND2X1_481/B vdd OAI21X1
XFILL_1_OAI21X1_1302 gnd vdd FILL
XFILL_1_OAI21X1_1313 gnd vdd FILL
XDFFPOSX1_705 BUFX2_343/A CLKBUF1_37/Y OAI21X1_959/Y gnd vdd DFFPOSX1
XOAI21X1_1137 NAND2X1_507/Y OR2X2_18/B BUFX4_239/Y gnd OAI21X1_1138/A vdd OAI21X1
XFILL_1_DFFPOSX1_903 gnd vdd FILL
XDFFPOSX1_716 BUFX2_383/A CLKBUF1_21/Y OAI21X1_981/Y gnd vdd DFFPOSX1
XDFFPOSX1_727 BUFX2_364/A CLKBUF1_38/Y OAI21X1_1003/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1335 gnd vdd FILL
XOAI21X1_1148 XNOR2X1_65/Y BUFX4_209/Y NAND2X1_524/Y gnd OAI21X1_1148/Y vdd OAI21X1
XFILL_1_DFFPOSX1_914 gnd vdd FILL
XFILL_1_OAI21X1_1346 gnd vdd FILL
XFILL_1_DFFPOSX1_925 gnd vdd FILL
XFILL_1_OAI21X1_1324 gnd vdd FILL
XFILL_1_OAI21X1_1357 gnd vdd FILL
XOAI21X1_1159 XNOR2X1_67/Y BUFX4_226/Y NAND2X1_535/Y gnd OAI21X1_1159/Y vdd OAI21X1
XDFFPOSX1_738 BUFX2_376/A CLKBUF1_37/Y OAI21X1_1025/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_126 gnd vdd FILL
XFILL_1_DFFPOSX1_936 gnd vdd FILL
XFILL_0_OAI21X1_115 gnd vdd FILL
XFILL_1_OAI21X1_308 gnd vdd FILL
XDFFPOSX1_749 BUFX2_46/A CLKBUF1_31/Y OAI21X1_1041/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_947 gnd vdd FILL
XFILL_0_OAI21X1_104 gnd vdd FILL
XFILL_1_OAI21X1_1379 gnd vdd FILL
XFILL_1_OAI21X1_1368 gnd vdd FILL
XFILL_1_DFFPOSX1_958 gnd vdd FILL
XFILL_0_OAI21X1_137 gnd vdd FILL
XFILL_0_OAI21X1_159 gnd vdd FILL
XFILL_0_OAI21X1_148 gnd vdd FILL
XFILL_1_DFFPOSX1_969 gnd vdd FILL
XFILL_1_OAI21X1_319 gnd vdd FILL
XFILL_6_DFFPOSX1_551 gnd vdd FILL
XFILL_6_DFFPOSX1_540 gnd vdd FILL
XFILL_6_DFFPOSX1_562 gnd vdd FILL
XFILL_0_BUFX4_36 gnd vdd FILL
XFILL_0_BUFX4_14 gnd vdd FILL
XFILL_0_BUFX4_25 gnd vdd FILL
XFILL_0_NAND2X1_132 gnd vdd FILL
XFILL_0_NAND2X1_110 gnd vdd FILL
XFILL_0_NAND2X1_121 gnd vdd FILL
XFILL_0_BUFX4_47 gnd vdd FILL
XFILL_0_BUFX4_69 gnd vdd FILL
XFILL_0_BUFX4_58 gnd vdd FILL
XFILL_1_NAND2X1_314 gnd vdd FILL
XFILL_0_NAND2X1_143 gnd vdd FILL
XFILL_0_DFFPOSX1_515 gnd vdd FILL
XFILL_0_NAND2X1_176 gnd vdd FILL
XFILL_1_NAND2X1_336 gnd vdd FILL
XFILL_0_DFFPOSX1_504 gnd vdd FILL
XFILL_1_NAND2X1_325 gnd vdd FILL
XFILL_0_18_1 gnd vdd FILL
XFILL_0_NAND2X1_154 gnd vdd FILL
XFILL_1_NAND2X1_347 gnd vdd FILL
XFILL_0_NAND2X1_165 gnd vdd FILL
XFILL_1_NAND2X1_358 gnd vdd FILL
XFILL_0_INVX1_190 gnd vdd FILL
XFILL_0_DFFPOSX1_537 gnd vdd FILL
XFILL_0_DFFPOSX1_526 gnd vdd FILL
XFILL_0_DFFPOSX1_548 gnd vdd FILL
XFILL_0_NAND2X1_187 gnd vdd FILL
XFILL_0_NAND2X1_198 gnd vdd FILL
XFILL_0_DFFPOSX1_559 gnd vdd FILL
XFILL_5_DFFPOSX1_130 gnd vdd FILL
XFILL_5_DFFPOSX1_152 gnd vdd FILL
XFILL_5_DFFPOSX1_141 gnd vdd FILL
XFILL_5_DFFPOSX1_185 gnd vdd FILL
XFILL_24_12_0 gnd vdd FILL
XFILL_5_DFFPOSX1_163 gnd vdd FILL
XFILL_5_DFFPOSX1_196 gnd vdd FILL
XFILL_5_DFFPOSX1_174 gnd vdd FILL
XOAI21X1_1660 BUFX4_248/Y BUFX4_361/Y BUFX2_742/A gnd OAI21X1_1661/C vdd OAI21X1
XOAI21X1_1693 BUFX4_123/Y INVX2_140/Y OAI21X1_1693/C gnd DFFPOSX1_59/D vdd OAI21X1
XOAI21X1_1682 BUFX4_2/A BUFX4_366/Y BUFX2_723/A gnd OAI21X1_1683/C vdd OAI21X1
XOAI21X1_1671 BUFX4_176/Y INVX2_129/Y OAI21X1_1671/C gnd DFFPOSX1_48/D vdd OAI21X1
XFILL_1_OAI21X1_820 gnd vdd FILL
XFILL_0_OR2X2_17 gnd vdd FILL
XFILL_1_OAI21X1_864 gnd vdd FILL
XFILL_1_OAI21X1_831 gnd vdd FILL
XFILL_1_OAI21X1_842 gnd vdd FILL
XFILL_0_OAI21X1_671 gnd vdd FILL
XFILL_1_OAI21X1_853 gnd vdd FILL
XFILL_0_OAI21X1_682 gnd vdd FILL
XFILL_0_OAI21X1_660 gnd vdd FILL
XNAND3X1_14 bundleStartMajId_i[52] INVX1_9/Y INVX4_30/A gnd OAI22X1_1/B vdd NAND3X1
XNAND3X1_36 INVX2_47/Y INVX1_44/A NOR3X1_9/Y gnd NOR3X1_11/C vdd NAND3X1
XNAND3X1_25 bundleStartMajId_i[8] bundleStartMajId_i[7] INVX2_46/A gnd OR2X2_13/A
+ vdd NAND3X1
XNAND3X1_47 bundleAddress_i[13] bundleAddress_i[12] AND2X2_24/Y gnd NOR3X1_13/C vdd
+ NAND3X1
XFILL_0_OAI21X1_693 gnd vdd FILL
XFILL_1_OAI21X1_897 gnd vdd FILL
XFILL_1_OAI21X1_886 gnd vdd FILL
XFILL_1_OAI21X1_875 gnd vdd FILL
XNAND3X1_69 bundleAddress_i[1] INVX4_49/A NOR2X1_231/Y gnd NAND3X1_69/Y vdd NAND3X1
XNAND3X1_58 INVX1_195/Y INVX1_211/A NOR3X1_17/Y gnd INVX1_213/A vdd NAND3X1
XFILL_5_17_1 gnd vdd FILL
XFILL_3_DFFPOSX1_12 gnd vdd FILL
XFILL_2_DFFPOSX1_609 gnd vdd FILL
XNOR2X1_36 NOR2X1_36/A NOR3X1_2/C gnd NOR2X1_37/B vdd NOR2X1
XBUFX2_707 BUFX2_707/A gnd pid2_o[27] vdd BUFX2
XNOR2X1_25 OR2X2_15/B INVX4_15/Y gnd INVX2_43/A vdd NOR2X1
XBUFX2_718 BUFX2_718/A gnd pid3_o[18] vdd BUFX2
XFILL_3_DFFPOSX1_23 gnd vdd FILL
XFILL_3_DFFPOSX1_34 gnd vdd FILL
XNOR2X1_14 OR2X2_3/Y NOR2X1_23/A gnd AND2X2_3/A vdd NOR2X1
XBUFX2_729 BUFX2_729/A gnd pid3_o[8] vdd BUFX2
XFILL_3_DFFPOSX1_45 gnd vdd FILL
XFILL_3_DFFPOSX1_56 gnd vdd FILL
XNOR2X1_47 NOR3X1_8/B NOR3X1_4/C gnd NOR2X1_47/Y vdd NOR2X1
XNOR2X1_69 NOR2X1_69/A NOR2X1_69/B gnd NOR2X1_69/Y vdd NOR2X1
XNOR2X1_58 NOR2X1_4/A INVX1_25/A gnd INVX4_29/A vdd NOR2X1
XFILL_3_DFFPOSX1_67 gnd vdd FILL
XFILL_3_DFFPOSX1_78 gnd vdd FILL
XFILL_3_DFFPOSX1_89 gnd vdd FILL
XFILL_29_11_0 gnd vdd FILL
XFILL_0_OAI21X1_1470 gnd vdd FILL
XFILL_0_OAI21X1_1481 gnd vdd FILL
XFILL_0_OAI21X1_1492 gnd vdd FILL
XFILL_0_BUFX2_1 gnd vdd FILL
XFILL_0_BUFX2_403 gnd vdd FILL
XFILL_0_BUFX2_414 gnd vdd FILL
XFILL_0_BUFX2_447 gnd vdd FILL
XFILL_0_BUFX2_425 gnd vdd FILL
XFILL_0_BUFX2_436 gnd vdd FILL
XFILL_0_BUFX2_469 gnd vdd FILL
XFILL_0_BUFX2_458 gnd vdd FILL
XFILL_0_NAND2X1_12 gnd vdd FILL
XFILL_4_12_0 gnd vdd FILL
XFILL_0_NAND2X1_23 gnd vdd FILL
XFILL_0_NAND2X1_34 gnd vdd FILL
XFILL_0_NAND2X1_56 gnd vdd FILL
XFILL_0_NAND2X1_45 gnd vdd FILL
XNOR2X1_115 INVX4_22/Y NOR3X1_8/C gnd INVX2_53/A vdd NOR2X1
XNOR2X1_104 NOR2X1_104/A INVX1_35/A gnd AND2X2_19/A vdd NOR2X1
XNOR2X1_126 INVX4_32/Y INVX2_93/Y gnd NOR2X1_126/Y vdd NOR2X1
XNOR2X1_148 INVX4_39/Y NOR2X1_148/B gnd NOR2X1_149/B vdd NOR2X1
XNOR2X1_137 INVX2_97/Y INVX1_188/Y gnd NOR2X1_137/Y vdd NOR2X1
XFILL_0_NAND2X1_67 gnd vdd FILL
XFILL_0_NAND2X1_89 gnd vdd FILL
XFILL_0_NAND2X1_78 gnd vdd FILL
XFILL_0_INVX2_1 gnd vdd FILL
XFILL_33_1_1 gnd vdd FILL
XNOR2X1_159 INVX2_78/Y INVX4_42/Y gnd NOR2X1_159/Y vdd NOR2X1
XFILL_16_2 gnd vdd FILL
XFILL_1_DFFPOSX1_700 gnd vdd FILL
XFILL_1_OAI21X1_1110 gnd vdd FILL
XFILL_1_OAI21X1_1121 gnd vdd FILL
XDFFPOSX1_513 BUFX2_543/A CLKBUF1_63/Y OAI21X1_578/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1132 gnd vdd FILL
XDFFPOSX1_502 BUFX2_531/A CLKBUF1_63/Y OAI21X1_552/Y gnd vdd DFFPOSX1
XDFFPOSX1_546 BUFX2_580/A CLKBUF1_70/Y OAI21X1_657/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_711 gnd vdd FILL
XFILL_1_OAI21X1_1143 gnd vdd FILL
XFILL_1_DFFPOSX1_722 gnd vdd FILL
XFILL_1_OAI21X1_1154 gnd vdd FILL
XDFFPOSX1_535 BUFX2_568/A CLKBUF1_91/Y OAI21X1_630/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_733 gnd vdd FILL
XDFFPOSX1_524 NOR2X1_81/A CLKBUF1_44/Y AOI21X1_12/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_970 gnd vdd FILL
XFILL_1_OAI21X1_1165 gnd vdd FILL
XFILL_1_DFFPOSX1_755 gnd vdd FILL
XFILL_1_DFFPOSX1_744 gnd vdd FILL
XFILL_1_OAI21X1_1176 gnd vdd FILL
XFILL_1_OAI21X1_105 gnd vdd FILL
XFILL_1_OAI21X1_116 gnd vdd FILL
XDFFPOSX1_568 BUFX2_598/A CLKBUF1_88/Y OAI21X1_718/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1198 gnd vdd FILL
XDFFPOSX1_579 INVX1_39/A CLKBUF1_60/Y OAI21X1_747/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1187 gnd vdd FILL
XFILL_0_BUFX2_992 gnd vdd FILL
XFILL_0_BUFX2_981 gnd vdd FILL
XFILL_1_DFFPOSX1_766 gnd vdd FILL
XDFFPOSX1_557 BUFX2_648/A CLKBUF1_46/Y OAI21X1_685/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_138 gnd vdd FILL
XFILL_1_OAI21X1_127 gnd vdd FILL
XFILL_1_OAI21X1_149 gnd vdd FILL
XFILL_1_DFFPOSX1_788 gnd vdd FILL
XFILL_1_DFFPOSX1_777 gnd vdd FILL
XNAND2X1_605 INVX1_206/Y NOR2X1_190/Y gnd NOR2X1_194/B vdd NAND2X1
XNAND2X1_627 bundleAddress_i[45] INVX4_51/A gnd NOR2X1_222/B vdd NAND2X1
XNAND2X1_616 NAND2X1_616/A NAND2X1_616/B gnd NAND2X1_616/Y vdd NAND2X1
XFILL_1_DFFPOSX1_799 gnd vdd FILL
XNAND2X1_649 BUFX2_390/A BUFX4_213/Y gnd NAND2X1_649/Y vdd NAND2X1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XINVX1_17 NOR3X1_2/C gnd INVX1_17/Y vdd INVX1
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XFILL_9_11_0 gnd vdd FILL
XNAND2X1_638 NAND2X1_638/A NAND3X1_65/Y gnd NAND2X1_638/Y vdd NAND2X1
XNAND2X1_91 BUFX2_404/A BUFX4_351/Y gnd NAND2X1_91/Y vdd NAND2X1
XNAND2X1_80 BUFX2_455/A BUFX4_387/Y gnd NAND2X1_80/Y vdd NAND2X1
XFILL_0_XNOR2X1_102 gnd vdd FILL
XFILL_10_18_0 gnd vdd FILL
XFILL_0_DFFPOSX1_323 gnd vdd FILL
XFILL_0_DFFPOSX1_301 gnd vdd FILL
XFILL_0_DFFPOSX1_312 gnd vdd FILL
XFILL_24_1_1 gnd vdd FILL
XFILL_1_NAND2X1_133 gnd vdd FILL
XFILL_0_DFFPOSX1_345 gnd vdd FILL
XFILL_0_DFFPOSX1_356 gnd vdd FILL
XFILL_1_NAND2X1_199 gnd vdd FILL
XFILL_1_NAND2X1_166 gnd vdd FILL
XFILL_0_DFFPOSX1_334 gnd vdd FILL
XFILL_1_NAND2X1_177 gnd vdd FILL
XFILL_0_DFFPOSX1_378 gnd vdd FILL
XFILL_0_DFFPOSX1_367 gnd vdd FILL
XFILL_0_DFFPOSX1_389 gnd vdd FILL
XFILL_3_DFFPOSX1_805 gnd vdd FILL
XFILL_3_DFFPOSX1_816 gnd vdd FILL
XFILL_3_DFFPOSX1_838 gnd vdd FILL
XFILL_3_DFFPOSX1_827 gnd vdd FILL
XFILL_3_DFFPOSX1_849 gnd vdd FILL
XOAI21X1_1490 NAND2X1_637/Y INVX1_223/A OAI21X1_1490/C gnd OAI21X1_1492/A vdd OAI21X1
XFILL_2_OAI21X1_810 gnd vdd FILL
XFILL_1_NOR2X1_211 gnd vdd FILL
XFILL_1_NOR2X1_222 gnd vdd FILL
XFILL_1_NOR2X1_200 gnd vdd FILL
XFILL_1_OAI21X1_650 gnd vdd FILL
XFILL_0_OAI21X1_490 gnd vdd FILL
XFILL_1_NOR2X1_233 gnd vdd FILL
XFILL_3_NOR3X1_1 gnd vdd FILL
XFILL_7_2_1 gnd vdd FILL
XFILL_1_OAI21X1_672 gnd vdd FILL
XFILL_1_OAI21X1_661 gnd vdd FILL
XFILL_15_17_0 gnd vdd FILL
XFILL_1_OAI21X1_694 gnd vdd FILL
XFILL_1_OAI21X1_683 gnd vdd FILL
XFILL_1_INVX1_166 gnd vdd FILL
XFILL_1_INVX1_177 gnd vdd FILL
XFILL_2_OAI21X1_887 gnd vdd FILL
XFILL_4_DFFPOSX1_13 gnd vdd FILL
XFILL_31_10_1 gnd vdd FILL
XBUFX2_504 BUFX2_504/A gnd majID2_o[12] vdd BUFX2
XFILL_4_DFFPOSX1_24 gnd vdd FILL
XBUFX2_515 BUFX2_515/A gnd majID2_o[2] vdd BUFX2
XFILL_2_DFFPOSX1_406 gnd vdd FILL
XBUFX2_526 BUFX2_526/A gnd majID3_o[50] vdd BUFX2
XFILL_2_DFFPOSX1_428 gnd vdd FILL
XFILL_2_DFFPOSX1_417 gnd vdd FILL
XFILL_4_DFFPOSX1_57 gnd vdd FILL
XFILL_4_DFFPOSX1_46 gnd vdd FILL
XFILL_2_DFFPOSX1_439 gnd vdd FILL
XBUFX2_559 BUFX2_559/A gnd majID3_o[20] vdd BUFX2
XBUFX2_537 BUFX2_537/A gnd majID3_o[40] vdd BUFX2
XBUFX2_548 BUFX2_548/A gnd majID3_o[30] vdd BUFX2
XFILL_4_DFFPOSX1_35 gnd vdd FILL
XFILL_4_DFFPOSX1_68 gnd vdd FILL
XFILL_4_DFFPOSX1_79 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XDFFPOSX1_1020 BUFX2_657/A CLKBUF1_11/Y OAI21X1_1597/Y gnd vdd DFFPOSX1
XFILL_0_DFFPOSX1_890 gnd vdd FILL
XDFFPOSX1_1031 BUFX2_669/A CLKBUF1_16/Y OAI21X1_1608/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_211 gnd vdd FILL
XFILL_0_BUFX2_200 gnd vdd FILL
XFILL_0_BUFX2_222 gnd vdd FILL
XFILL_0_BUFX2_255 gnd vdd FILL
XFILL_0_BUFX2_233 gnd vdd FILL
XFILL_0_BUFX2_244 gnd vdd FILL
XFILL_0_BUFX2_299 gnd vdd FILL
XFILL_0_BUFX2_277 gnd vdd FILL
XFILL_0_BUFX2_288 gnd vdd FILL
XFILL_2_AND2X2_26 gnd vdd FILL
XFILL_0_BUFX2_266 gnd vdd FILL
XFILL_33_18_0 gnd vdd FILL
XFILL_35_9_0 gnd vdd FILL
XFILL_2_DFFPOSX1_951 gnd vdd FILL
XFILL_2_DFFPOSX1_940 gnd vdd FILL
XFILL_2_DFFPOSX1_962 gnd vdd FILL
XFILL_2_DFFPOSX1_984 gnd vdd FILL
XFILL_2_DFFPOSX1_973 gnd vdd FILL
XFILL_2_DFFPOSX1_995 gnd vdd FILL
XFILL_0_NAND3X1_7 gnd vdd FILL
XOAI21X1_429 OAI21X1_429/A BUFX4_224/Y OAI21X1_429/C gnd OAI21X1_429/Y vdd OAI21X1
XOAI21X1_407 OAI21X1_407/A BUFX4_199/Y OAI21X1_407/C gnd OAI21X1_407/Y vdd OAI21X1
XOAI21X1_418 NOR2X1_6/B OR2X2_1/Y OAI21X1_418/C gnd OAI21X1_419/A vdd OAI21X1
XFILL_3_XNOR2X1_31 gnd vdd FILL
XFILL_3_XNOR2X1_20 gnd vdd FILL
XFILL_3_XNOR2X1_64 gnd vdd FILL
XFILL_3_XNOR2X1_75 gnd vdd FILL
XDFFPOSX1_321 BUFX2_991/A CLKBUF1_49/Y OAI21X1_259/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_53 gnd vdd FILL
XDFFPOSX1_310 BUFX2_979/A CLKBUF1_77/Y OAI21X1_237/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_541 gnd vdd FILL
XFILL_3_XNOR2X1_97 gnd vdd FILL
XFILL_1_DFFPOSX1_530 gnd vdd FILL
XDFFPOSX1_343 BUFX2_1016/A CLKBUF1_69/Y OAI21X1_303/Y gnd vdd DFFPOSX1
XDFFPOSX1_354 BUFX2_1028/A CLKBUF1_4/Y OAI21X1_325/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_86 gnd vdd FILL
XDFFPOSX1_332 BUFX2_1004/A CLKBUF1_83/Y OAI21X1_281/Y gnd vdd DFFPOSX1
XDFFPOSX1_365 BUFX2_456/A CLKBUF1_6/Y OAI21X1_337/Y gnd vdd DFFPOSX1
XFILL_38_17_0 gnd vdd FILL
XNAND2X1_402 BUFX2_1/A BUFX4_322/Y gnd NAND2X1_402/Y vdd NAND2X1
XFILL_1_DFFPOSX1_563 gnd vdd FILL
XDFFPOSX1_398 BUFX2_430/A CLKBUF1_84/Y OAI21X1_370/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_574 gnd vdd FILL
XFILL_1_DFFPOSX1_552 gnd vdd FILL
XDFFPOSX1_376 BUFX2_406/A CLKBUF1_33/Y OAI21X1_348/Y gnd vdd DFFPOSX1
XDFFPOSX1_387 BUFX2_418/A CLKBUF1_15/Y OAI21X1_359/Y gnd vdd DFFPOSX1
XNAND2X1_413 BUFX2_4/A BUFX4_386/Y gnd NAND2X1_413/Y vdd NAND2X1
XFILL_1_DFFPOSX1_585 gnd vdd FILL
XNAND2X1_435 BUFX2_28/A BUFX4_381/Y gnd NAND2X1_435/Y vdd NAND2X1
XFILL_1_DFFPOSX1_596 gnd vdd FILL
XNAND2X1_424 BUFX2_16/A OAI21X1_4/A gnd NAND2X1_424/Y vdd NAND2X1
XNAND2X1_468 BUFX2_77/A BUFX4_197/Y gnd NAND2X1_468/Y vdd NAND2X1
XNAND2X1_446 BUFX2_40/A BUFX4_381/Y gnd NAND2X1_446/Y vdd NAND2X1
XNAND2X1_457 BUFX2_52/A BUFX4_357/Y gnd NAND2X1_457/Y vdd NAND2X1
XNAND2X1_479 BUFX2_127/A BUFX4_198/Y gnd NAND2X1_479/Y vdd NAND2X1
XFILL_26_9_0 gnd vdd FILL
XFILL_1_9_0 gnd vdd FILL
XFILL_0_DFFPOSX1_131 gnd vdd FILL
XFILL_0_DFFPOSX1_120 gnd vdd FILL
XFILL_1_XNOR2X1_103 gnd vdd FILL
XFILL_0_DFFPOSX1_153 gnd vdd FILL
XFILL_0_DFFPOSX1_175 gnd vdd FILL
XFILL_0_DFFPOSX1_164 gnd vdd FILL
XFILL_1_BUFX2_913 gnd vdd FILL
XFILL_1_BUFX2_902 gnd vdd FILL
XFILL_0_DFFPOSX1_142 gnd vdd FILL
XFILL_0_DFFPOSX1_197 gnd vdd FILL
XFILL_0_DFFPOSX1_186 gnd vdd FILL
XFILL_1_BUFX2_946 gnd vdd FILL
XFILL_1_BUFX2_957 gnd vdd FILL
XOAI21X1_930 BUFX4_11/A BUFX4_332/Y BUFX2_328/A gnd OAI21X1_931/C vdd OAI21X1
XFILL_1_BUFX2_968 gnd vdd FILL
XFILL_3_DFFPOSX1_613 gnd vdd FILL
XOAI21X1_952 BUFX4_1/Y BUFX4_330/Y BUFX2_340/A gnd OAI21X1_953/C vdd OAI21X1
XFILL_3_DFFPOSX1_602 gnd vdd FILL
XOAI21X1_941 BUFX4_144/Y INVX1_125/Y OAI21X1_941/C gnd OAI21X1_941/Y vdd OAI21X1
XOAI21X1_985 BUFX4_293/Y INVX1_147/Y OAI21X1_985/C gnd OAI21X1_985/Y vdd OAI21X1
XOAI21X1_974 BUFX4_137/Y BUFX4_53/Y BUFX2_358/A gnd OAI21X1_975/C vdd OAI21X1
XFILL_3_DFFPOSX1_624 gnd vdd FILL
XOAI21X1_963 BUFX4_153/Y INVX1_136/Y OAI21X1_963/C gnd OAI21X1_963/Y vdd OAI21X1
XFILL_3_DFFPOSX1_635 gnd vdd FILL
XFILL_3_DFFPOSX1_646 gnd vdd FILL
XFILL_3_DFFPOSX1_679 gnd vdd FILL
XFILL_3_DFFPOSX1_668 gnd vdd FILL
XFILL_3_DFFPOSX1_657 gnd vdd FILL
XOAI21X1_996 BUFX4_139/Y BUFX4_68/Y BUFX2_361/A gnd OAI21X1_997/C vdd OAI21X1
XINVX2_60 bundleAddress_i[56] gnd INVX2_60/Y vdd INVX2
XINVX2_82 bundleAddress_i[16] gnd INVX2_82/Y vdd INVX2
XINVX2_71 bundleAddress_i[37] gnd INVX2_71/Y vdd INVX2
XFILL_2_OAI21X1_640 gnd vdd FILL
XFILL_1_OAI21X1_480 gnd vdd FILL
XINVX2_93 INVX2_93/A gnd INVX2_93/Y vdd INVX2
XFILL_1_OAI21X1_491 gnd vdd FILL
XFILL_2_OAI21X1_662 gnd vdd FILL
XFILL_2_OAI21X1_695 gnd vdd FILL
XBUFX2_301 BUFX2_301/A gnd instr2_o[15] vdd BUFX2
XFILL_2_DFFPOSX1_203 gnd vdd FILL
XFILL_0_AOI21X1_1 gnd vdd FILL
XFILL_0_NAND2X1_709 gnd vdd FILL
XBUFX2_323 BUFX2_323/A gnd instr2_o[23] vdd BUFX2
XFILL_2_DFFPOSX1_214 gnd vdd FILL
XFILL_2_DFFPOSX1_225 gnd vdd FILL
XFILL_17_9_0 gnd vdd FILL
XBUFX2_345 BUFX2_345/A gnd instr3_o[4] vdd BUFX2
XBUFX2_334 BUFX2_334/A gnd instr3_o[14] vdd BUFX2
XBUFX2_312 BUFX2_312/A gnd instr2_o[5] vdd BUFX2
XFILL_2_DFFPOSX1_236 gnd vdd FILL
XBUFX2_378 BUFX2_378/A gnd instr4_o[3] vdd BUFX2
XFILL_2_DFFPOSX1_258 gnd vdd FILL
XFILL_5_DFFPOSX1_36 gnd vdd FILL
XFILL_5_DFFPOSX1_25 gnd vdd FILL
XFILL_5_DFFPOSX1_14 gnd vdd FILL
XFILL_2_DFFPOSX1_247 gnd vdd FILL
XBUFX2_356 BUFX2_356/A gnd instr3_o[22] vdd BUFX2
XBUFX2_367 BUFX2_367/A gnd instr4_o[13] vdd BUFX2
XFILL_2_DFFPOSX1_269 gnd vdd FILL
XFILL_5_DFFPOSX1_69 gnd vdd FILL
XFILL_5_DFFPOSX1_58 gnd vdd FILL
XBUFX2_389 BUFX2_389/A gnd is64b1_o vdd BUFX2
XFILL_5_DFFPOSX1_47 gnd vdd FILL
XFILL_1_NOR3X1_17 gnd vdd FILL
XOAI21X1_34 INVX2_172/Y BUFX4_191/Y OAI21X1_34/C gnd OAI21X1_34/Y vdd OAI21X1
XOAI21X1_23 INVX2_161/Y BUFX4_216/Y OAI21X1_23/C gnd OAI21X1_23/Y vdd OAI21X1
XOAI21X1_12 INVX2_150/Y BUFX4_197/Y OAI21X1_12/C gnd OAI21X1_12/Y vdd OAI21X1
XFILL_5_DFFPOSX1_718 gnd vdd FILL
XOAI21X1_45 INVX2_183/Y BUFX4_200/Y OAI21X1_45/C gnd OAI21X1_45/Y vdd OAI21X1
XFILL_5_DFFPOSX1_707 gnd vdd FILL
XOAI21X1_56 INVX2_194/Y BUFX4_191/Y OAI21X1_56/C gnd OAI21X1_56/Y vdd OAI21X1
XFILL_1_BUFX4_250 gnd vdd FILL
XFILL_1_BUFX4_272 gnd vdd FILL
XFILL_5_DFFPOSX1_729 gnd vdd FILL
XOAI21X1_78 BUFX4_98/Y BUFX4_321/Y BUFX2_928/A gnd OAI21X1_79/C vdd OAI21X1
XFILL_1_BUFX4_261 gnd vdd FILL
XOAI21X1_67 INVX2_3/Y OAI21X1_9/B OAI21X1_67/C gnd OAI21X1_67/Y vdd OAI21X1
XFILL_1_BUFX4_283 gnd vdd FILL
XFILL_1_BUFX4_294 gnd vdd FILL
XOAI21X1_89 BUFX4_153/Y INVX2_154/Y OAI21X1_89/C gnd OAI21X1_89/Y vdd OAI21X1
XFILL_22_15_1 gnd vdd FILL
XFILL_0_DFFPOSX1_10 gnd vdd FILL
XFILL_0_DFFPOSX1_21 gnd vdd FILL
XFILL_0_DFFPOSX1_32 gnd vdd FILL
XFILL_0_DFFPOSX1_43 gnd vdd FILL
XFILL_4_DFFPOSX1_308 gnd vdd FILL
XFILL_0_DFFPOSX1_76 gnd vdd FILL
XFILL_4_DFFPOSX1_319 gnd vdd FILL
XFILL_0_DFFPOSX1_54 gnd vdd FILL
XFILL_0_DFFPOSX1_65 gnd vdd FILL
XFILL_38_0_1 gnd vdd FILL
XFILL_0_DFFPOSX1_87 gnd vdd FILL
XFILL_0_DFFPOSX1_98 gnd vdd FILL
XBUFX2_890 BUFX2_890/A gnd tid2_o[10] vdd BUFX2
XFILL_2_DFFPOSX1_792 gnd vdd FILL
XFILL_2_DFFPOSX1_770 gnd vdd FILL
XFILL_2_DFFPOSX1_781 gnd vdd FILL
XFILL_0_NOR2X1_230 gnd vdd FILL
XFILL_27_14_1 gnd vdd FILL
XOAI21X1_204 BUFX4_177/Y BUFX4_74/Y BUFX2_981/A gnd OAI21X1_205/C vdd OAI21X1
XOAI21X1_215 INVX2_153/Y BUFX4_297/Y OAI21X1_215/C gnd OAI21X1_215/Y vdd OAI21X1
XOAI21X1_237 INVX2_164/Y BUFX4_294/Y OAI21X1_237/C gnd OAI21X1_237/Y vdd OAI21X1
XOAI21X1_226 BUFX4_163/Y BUFX4_30/Y BUFX2_974/A gnd OAI21X1_227/C vdd OAI21X1
XOAI21X1_248 BUFX4_164/Y BUFX4_44/Y BUFX2_986/A gnd OAI21X1_249/C vdd OAI21X1
XOAI21X1_259 INVX2_175/Y BUFX4_294/Y OAI21X1_259/C gnd OAI21X1_259/Y vdd OAI21X1
XFILL_21_10_0 gnd vdd FILL
XAND2X2_26 AND2X2_26/A INVX1_201/Y gnd AND2X2_26/Y vdd AND2X2
XAND2X2_15 NOR2X1_84/Y INVX1_32/Y gnd NOR2X1_85/B vdd AND2X2
XDFFPOSX1_173 BUFX2_904/A CLKBUF1_1/Y OAI21X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_151 BUFX2_824/A CLKBUF1_26/Y OAI21X1_1825/Y gnd vdd DFFPOSX1
XDFFPOSX1_162 NAND2X1_6/A CLKBUF1_4/Y OAI21X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_140 BUFX2_812/A CLKBUF1_2/Y OAI21X1_1814/Y gnd vdd DFFPOSX1
XDFFPOSX1_195 BUFX2_866/A CLKBUF1_78/Y OAI21X1_39/Y gnd vdd DFFPOSX1
XNAND2X1_210 BUFX2_487/A BUFX4_224/Y gnd OAI21X1_454/C vdd NAND2X1
XFILL_1_DFFPOSX1_382 gnd vdd FILL
XFILL_0_NOR3X1_5 gnd vdd FILL
XFILL_1_DFFPOSX1_393 gnd vdd FILL
XFILL_1_DFFPOSX1_360 gnd vdd FILL
XDFFPOSX1_184 BUFX2_854/A CLKBUF1_18/Y OAI21X1_28/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_371 gnd vdd FILL
XNAND2X1_243 bundleStartMajId_i[12] INVX2_45/Y gnd NOR3X1_8/B vdd NAND2X1
XNAND2X1_232 AND2X2_7/A AND2X2_7/B gnd NOR2X1_42/A vdd NAND2X1
XNAND2X1_221 bundleStartMajId_i[23] bundleStartMajId_i[22] gnd NOR2X1_36/A vdd NAND2X1
XNAND2X1_265 NAND2X1_265/A NAND3X1_13/Y gnd NAND2X1_265/Y vdd NAND2X1
XFILL_4_DFFPOSX1_820 gnd vdd FILL
XNAND2X1_254 XNOR2X1_23/A OAI21X1_488/Y gnd OAI21X1_489/A vdd NAND2X1
XNAND2X1_287 bundleStartMajId_i[32] bundleStartMajId_i[31] gnd NOR2X1_74/B vdd NAND2X1
XNAND2X1_276 OR2X2_10/B OAI21X1_545/Y gnd OAI21X1_546/A vdd NAND2X1
XFILL_4_DFFPOSX1_831 gnd vdd FILL
XFILL_29_0_1 gnd vdd FILL
XFILL_4_DFFPOSX1_853 gnd vdd FILL
XNAND2X1_298 INVX1_18/Y INVX2_50/A gnd OR2X2_11/A vdd NAND2X1
XFILL_4_DFFPOSX1_842 gnd vdd FILL
XFILL_4_DFFPOSX1_864 gnd vdd FILL
XFILL_4_0_1 gnd vdd FILL
XFILL_4_DFFPOSX1_875 gnd vdd FILL
XFILL_4_DFFPOSX1_886 gnd vdd FILL
XFILL_4_DFFPOSX1_897 gnd vdd FILL
XFILL_2_15_1 gnd vdd FILL
XFILL_0_OAI21X1_4 gnd vdd FILL
XFILL_2_XNOR2X1_104 gnd vdd FILL
XFILL_1_BUFX2_710 gnd vdd FILL
XFILL_1_BUFX2_721 gnd vdd FILL
XFILL_0_BUFX2_80 gnd vdd FILL
XFILL_0_BUFX2_91 gnd vdd FILL
XFILL_1_BUFX2_754 gnd vdd FILL
XFILL_0_BUFX4_306 gnd vdd FILL
XFILL_1_BUFX2_743 gnd vdd FILL
XFILL_1_BUFX2_765 gnd vdd FILL
XFILL_0_BUFX4_328 gnd vdd FILL
XFILL_0_BUFX4_339 gnd vdd FILL
XFILL_0_BUFX4_317 gnd vdd FILL
XOAI21X1_760 INVX1_41/A OR2X2_8/B INVX4_17/Y gnd OAI21X1_761/C vdd OAI21X1
XFILL_1_NOR2X1_83 gnd vdd FILL
XFILL_3_DFFPOSX1_421 gnd vdd FILL
XFILL_3_DFFPOSX1_410 gnd vdd FILL
XFILL_1_BUFX2_798 gnd vdd FILL
XOAI21X1_782 OAI21X1_782/A BUFX4_289/Y OAI21X1_782/C gnd OAI21X1_782/Y vdd OAI21X1
XOAI21X1_771 BUFX4_175/Y BUFX4_31/Y BUFX2_620/A gnd OAI21X1_772/C vdd OAI21X1
XOAI21X1_793 INVX4_31/Y OAI21X1_793/B INVX2_32/Y gnd OAI21X1_794/C vdd OAI21X1
XFILL_3_DFFPOSX1_443 gnd vdd FILL
XFILL_3_DFFPOSX1_432 gnd vdd FILL
XFILL_3_DFFPOSX1_454 gnd vdd FILL
XFILL_1_OAI21X1_1709 gnd vdd FILL
XFILL_3_DFFPOSX1_476 gnd vdd FILL
XFILL_3_DFFPOSX1_498 gnd vdd FILL
XFILL_3_DFFPOSX1_487 gnd vdd FILL
XFILL_3_DFFPOSX1_465 gnd vdd FILL
XFILL_6_DFFPOSX1_936 gnd vdd FILL
XFILL_6_DFFPOSX1_947 gnd vdd FILL
XFILL_6_DFFPOSX1_969 gnd vdd FILL
XFILL_6_DFFPOSX1_958 gnd vdd FILL
XFILL_7_14_1 gnd vdd FILL
XFILL_2_OAI21X1_470 gnd vdd FILL
XFILL_0_NAND2X1_517 gnd vdd FILL
XBUFX2_120 BUFX2_120/A gnd addr2_o[4] vdd BUFX2
XFILL_2_XNOR2X1_50 gnd vdd FILL
XFILL_0_NAND2X1_506 gnd vdd FILL
XBUFX2_131 BUFX2_131/A gnd addr3_o[53] vdd BUFX2
XBUFX2_153 BUFX2_153/A gnd addr3_o[33] vdd BUFX2
XFILL_0_NAND2X1_528 gnd vdd FILL
XFILL_2_XNOR2X1_72 gnd vdd FILL
XFILL_2_XNOR2X1_83 gnd vdd FILL
XFILL_0_NAND2X1_539 gnd vdd FILL
XFILL_1_10_0 gnd vdd FILL
XFILL_2_XNOR2X1_61 gnd vdd FILL
XBUFX2_142 BUFX2_142/A gnd addr3_o[43] vdd BUFX2
XFILL_6_DFFPOSX1_26 gnd vdd FILL
XBUFX2_186 BUFX2_186/A gnd addr3_o[3] vdd BUFX2
XBUFX2_175 BUFX2_175/A gnd addr3_o[13] vdd BUFX2
XFILL_1_NAND2X1_5 gnd vdd FILL
XFILL_2_XNOR2X1_94 gnd vdd FILL
XBUFX2_164 BUFX2_164/A gnd addr3_o[23] vdd BUFX2
XBUFX2_197 BUFX2_197/A gnd addr4_o[51] vdd BUFX2
XFILL_6_DFFPOSX1_59 gnd vdd FILL
XFILL_6_DFFPOSX1_37 gnd vdd FILL
XFILL_32_7_0 gnd vdd FILL
XFILL_6_DFFPOSX1_48 gnd vdd FILL
XFILL_5_DFFPOSX1_515 gnd vdd FILL
XFILL_5_DFFPOSX1_526 gnd vdd FILL
XFILL_5_DFFPOSX1_504 gnd vdd FILL
XFILL_5_DFFPOSX1_537 gnd vdd FILL
XFILL_5_DFFPOSX1_548 gnd vdd FILL
XFILL_5_DFFPOSX1_559 gnd vdd FILL
XBUFX2_1001 BUFX2_1001/A gnd tid4_o[25] vdd BUFX2
XBUFX2_1012 BUFX2_1012/A gnd tid4_o[15] vdd BUFX2
XBUFX2_1023 BUFX2_1023/A gnd tid4_o[5] vdd BUFX2
XCLKBUF1_24 BUFX4_84/Y gnd CLKBUF1_24/Y vdd CLKBUF1
XCLKBUF1_13 BUFX4_90/Y gnd CLKBUF1_13/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_127 gnd vdd FILL
XFILL_1_DFFPOSX1_11 gnd vdd FILL
XCLKBUF1_57 BUFX4_92/Y gnd CLKBUF1_57/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_116 gnd vdd FILL
XCLKBUF1_35 BUFX4_86/Y gnd CLKBUF1_35/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_22 gnd vdd FILL
XFILL_4_DFFPOSX1_105 gnd vdd FILL
XCLKBUF1_46 BUFX4_90/Y gnd CLKBUF1_46/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_138 gnd vdd FILL
XFILL_1_DFFPOSX1_44 gnd vdd FILL
XFILL_4_DFFPOSX1_149 gnd vdd FILL
XCLKBUF1_68 BUFX4_92/Y gnd CLKBUF1_68/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_55 gnd vdd FILL
XCLKBUF1_79 BUFX4_84/Y gnd CLKBUF1_79/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_33 gnd vdd FILL
XFILL_1_DFFPOSX1_66 gnd vdd FILL
XFILL_1_DFFPOSX1_77 gnd vdd FILL
XFILL_1_DFFPOSX1_88 gnd vdd FILL
XFILL_2_BUFX4_215 gnd vdd FILL
XFILL_1_DFFPOSX1_99 gnd vdd FILL
XFILL_0_OAI21X1_1800 gnd vdd FILL
XFILL_2_BUFX4_248 gnd vdd FILL
XFILL_0_OAI21X1_1811 gnd vdd FILL
XFILL_0_OAI21X1_1822 gnd vdd FILL
XFILL_23_7_0 gnd vdd FILL
XINVX1_109 bundle_i[95] gnd INVX1_109/Y vdd INVX1
XFILL_3_XNOR2X1_8 gnd vdd FILL
XFILL_1_DFFPOSX1_190 gnd vdd FILL
XFILL_0_INVX2_19 gnd vdd FILL
XFILL_6_8_0 gnd vdd FILL
XFILL_4_DFFPOSX1_672 gnd vdd FILL
XFILL_4_DFFPOSX1_650 gnd vdd FILL
XFILL_4_DFFPOSX1_661 gnd vdd FILL
XFILL_4_DFFPOSX1_683 gnd vdd FILL
XFILL_4_DFFPOSX1_694 gnd vdd FILL
XFILL_12_15_0 gnd vdd FILL
XFILL_0_CLKBUF1_9 gnd vdd FILL
XFILL_14_7_0 gnd vdd FILL
XFILL_4_CLKBUF1_8 gnd vdd FILL
XFILL_0_BUFX4_103 gnd vdd FILL
XFILL_0_BUFX4_114 gnd vdd FILL
XFILL_1_BUFX2_551 gnd vdd FILL
XFILL_1_BUFX2_562 gnd vdd FILL
XFILL_0_BUFX4_136 gnd vdd FILL
XFILL_1_BUFX2_595 gnd vdd FILL
XFILL_0_BUFX4_125 gnd vdd FILL
XFILL_0_BUFX4_147 gnd vdd FILL
XFILL_1_OAI21X1_1506 gnd vdd FILL
XFILL_0_BUFX4_158 gnd vdd FILL
XOAI21X1_1319 OAI21X1_1319/A BUFX4_152/Y OAI21X1_1319/C gnd OAI21X1_1319/Y vdd OAI21X1
XOAI21X1_1308 BUFX4_4/Y BUFX4_370/Y BUFX2_159/A gnd OAI21X1_1309/C vdd OAI21X1
XFILL_3_DFFPOSX1_273 gnd vdd FILL
XFILL_3_DFFPOSX1_262 gnd vdd FILL
XFILL_3_DFFPOSX1_240 gnd vdd FILL
XFILL_3_DFFPOSX1_251 gnd vdd FILL
XFILL_1_OAI21X1_1528 gnd vdd FILL
XFILL_1_OAI21X1_1517 gnd vdd FILL
XDFFPOSX1_909 BUFX2_160/A CLKBUF1_77/Y OAI21X1_1311/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1539 gnd vdd FILL
XFILL_0_BUFX4_169 gnd vdd FILL
XFILL_1_BUFX2_36 gnd vdd FILL
XOAI21X1_590 OAI21X1_590/A BUFX4_131/Y OAI21X1_590/C gnd OAI21X1_590/Y vdd OAI21X1
XFILL_3_DFFPOSX1_284 gnd vdd FILL
XFILL_0_OAI21X1_308 gnd vdd FILL
XFILL_3_DFFPOSX1_295 gnd vdd FILL
XFILL_1_BUFX2_58 gnd vdd FILL
XFILL_1_BUFX2_47 gnd vdd FILL
XFILL_0_OAI21X1_319 gnd vdd FILL
XFILL_6_DFFPOSX1_700 gnd vdd FILL
XFILL_6_DFFPOSX1_711 gnd vdd FILL
XFILL_6_DFFPOSX1_744 gnd vdd FILL
XFILL_6_DFFPOSX1_722 gnd vdd FILL
XFILL_6_DFFPOSX1_733 gnd vdd FILL
XFILL_17_14_0 gnd vdd FILL
XFILL_4_2 gnd vdd FILL
XFILL_5_DFFPOSX1_3 gnd vdd FILL
XFILL_30_16_0 gnd vdd FILL
XFILL_0_NAND2X1_303 gnd vdd FILL
XFILL_0_NAND2X1_325 gnd vdd FILL
XFILL_0_NAND2X1_314 gnd vdd FILL
XFILL_39_1 gnd vdd FILL
XFILL_0_NAND2X1_358 gnd vdd FILL
XFILL_0_OAI21X1_1107 gnd vdd FILL
XFILL_0_OAI21X1_1118 gnd vdd FILL
XFILL_0_OAI21X1_1129 gnd vdd FILL
XFILL_0_NAND2X1_336 gnd vdd FILL
XFILL_1_NAND2X1_518 gnd vdd FILL
XFILL_0_NAND2X1_347 gnd vdd FILL
XFILL_1_NOR2X1_5 gnd vdd FILL
XFILL_1_NAND2X1_507 gnd vdd FILL
XFILL_0_DFFPOSX1_719 gnd vdd FILL
XFILL_0_DFFPOSX1_708 gnd vdd FILL
XFILL_0_NAND2X1_369 gnd vdd FILL
XFILL_1_DFFPOSX1_1020 gnd vdd FILL
XFILL_1_DFFPOSX1_1031 gnd vdd FILL
XFILL_5_DFFPOSX1_301 gnd vdd FILL
XFILL_5_DFFPOSX1_345 gnd vdd FILL
XFILL_5_DFFPOSX1_323 gnd vdd FILL
XFILL_5_DFFPOSX1_312 gnd vdd FILL
XFILL_5_DFFPOSX1_334 gnd vdd FILL
XFILL_5_DFFPOSX1_356 gnd vdd FILL
XFILL_5_DFFPOSX1_378 gnd vdd FILL
XFILL_5_DFFPOSX1_367 gnd vdd FILL
XFILL_5_DFFPOSX1_389 gnd vdd FILL
XFILL_1_NAND2X1_38 gnd vdd FILL
XFILL_1_NAND2X1_27 gnd vdd FILL
XINVX4_17 bundleStartMajId_i[27] gnd INVX4_17/Y vdd INVX4
XOAI21X1_1820 OAI21X1_6/A INVX2_192/Y NAND2X1_761/Y gnd OAI21X1_1820/Y vdd OAI21X1
XINVX4_28 INVX4_28/A gnd INVX4_28/Y vdd INVX4
XINVX4_39 bundleAddress_i[32] gnd INVX4_39/Y vdd INVX4
XFILL_1_NAND2X1_49 gnd vdd FILL
XFILL_0_OAI21X1_831 gnd vdd FILL
XFILL_0_OAI21X1_820 gnd vdd FILL
XFILL_0_OAI21X1_864 gnd vdd FILL
XFILL_0_OAI21X1_842 gnd vdd FILL
XFILL_0_OAI21X1_875 gnd vdd FILL
XFILL_0_OAI21X1_853 gnd vdd FILL
XFILL_35_15_0 gnd vdd FILL
XFILL_0_OAI21X1_897 gnd vdd FILL
XFILL_0_OAI21X1_886 gnd vdd FILL
XFILL_2_DFFPOSX1_12 gnd vdd FILL
XFILL_2_DFFPOSX1_45 gnd vdd FILL
XFILL_2_DFFPOSX1_23 gnd vdd FILL
XFILL_2_DFFPOSX1_34 gnd vdd FILL
XFILL_2_DFFPOSX1_78 gnd vdd FILL
XFILL_2_DFFPOSX1_89 gnd vdd FILL
XFILL_2_DFFPOSX1_56 gnd vdd FILL
XFILL_2_DFFPOSX1_67 gnd vdd FILL
XFILL_0_OAI21X1_1630 gnd vdd FILL
XFILL_0_OAI21X1_1652 gnd vdd FILL
XFILL_0_OAI21X1_1641 gnd vdd FILL
XFILL_0_OAI21X1_1674 gnd vdd FILL
XFILL_0_OAI21X1_1663 gnd vdd FILL
XFILL_0_OAI21X1_1685 gnd vdd FILL
XFILL_0_OAI21X1_1696 gnd vdd FILL
XFILL_0_BUFX4_5 gnd vdd FILL
XFILL_5_DFFPOSX1_890 gnd vdd FILL
XFILL_0_BUFX2_618 gnd vdd FILL
XFILL_0_BUFX2_629 gnd vdd FILL
XFILL_0_BUFX2_607 gnd vdd FILL
XFILL_4_DFFPOSX1_1013 gnd vdd FILL
XFILL_4_DFFPOSX1_1024 gnd vdd FILL
XFILL_1_XNOR2X1_91 gnd vdd FILL
XFILL_1_XNOR2X1_80 gnd vdd FILL
XFILL_4_DFFPOSX1_1002 gnd vdd FILL
XBUFX4_204 BUFX4_25/Y gnd BUFX4_204/Y vdd BUFX4
XBUFX4_215 BUFX4_20/Y gnd BUFX4_215/Y vdd BUFX4
XBUFX4_237 BUFX4_20/Y gnd BUFX4_237/Y vdd BUFX4
XBUFX4_226 BUFX4_21/Y gnd BUFX4_226/Y vdd BUFX4
XFILL_0_INVX2_125 gnd vdd FILL
XBUFX4_248 INVX8_5/Y gnd BUFX4_248/Y vdd BUFX4
XFILL_4_DFFPOSX1_480 gnd vdd FILL
XBUFX4_259 INVX8_5/Y gnd BUFX4_6/A vdd BUFX4
XFILL_0_INVX2_103 gnd vdd FILL
XFILL_4_DFFPOSX1_491 gnd vdd FILL
XFILL_0_INVX2_114 gnd vdd FILL
XFILL_0_INVX2_158 gnd vdd FILL
XFILL_2_OAI21X1_1768 gnd vdd FILL
XFILL_0_INVX2_136 gnd vdd FILL
XFILL_0_INVX2_147 gnd vdd FILL
XFILL_0_INVX2_169 gnd vdd FILL
XFILL_0_INVX4_5 gnd vdd FILL
XFILL_1_BUFX2_370 gnd vdd FILL
XOAI21X1_1116 NOR2X1_126/Y NAND2X1_481/Y NAND2X1_479/Y gnd OAI21X1_1116/Y vdd OAI21X1
XOAI21X1_1105 INVX4_32/Y INVX1_183/A OAI21X1_1105/C gnd OAI21X1_1106/A vdd OAI21X1
XOAI21X1_1127 INVX2_95/Y NOR2X1_185/A NAND2X1_492/Y gnd OAI21X1_1128/A vdd OAI21X1
XFILL_1_OAI21X1_1303 gnd vdd FILL
XFILL_1_BUFX2_392 gnd vdd FILL
XFILL_1_OAI21X1_1314 gnd vdd FILL
XOAI21X1_1138 OAI21X1_1138/A NOR2X1_138/Y NAND2X1_508/Y gnd OAI21X1_1138/Y vdd OAI21X1
XOAI21X1_1149 XNOR2X1_66/Y BUFX4_202/Y NAND2X1_525/Y gnd OAI21X1_1149/Y vdd OAI21X1
XFILL_1_OAI21X1_1336 gnd vdd FILL
XFILL_1_DFFPOSX1_904 gnd vdd FILL
XFILL_1_DFFPOSX1_915 gnd vdd FILL
XFILL_1_OAI21X1_1325 gnd vdd FILL
XFILL_1_OAI21X1_1347 gnd vdd FILL
XDFFPOSX1_728 BUFX2_365/A CLKBUF1_38/Y OAI21X1_1005/Y gnd vdd DFFPOSX1
XDFFPOSX1_706 BUFX2_344/A CLKBUF1_54/Y OAI21X1_961/Y gnd vdd DFFPOSX1
XDFFPOSX1_717 BUFX2_384/A CLKBUF1_62/Y OAI21X1_983/Y gnd vdd DFFPOSX1
XDFFPOSX1_739 BUFX2_377/A CLKBUF1_56/Y OAI21X1_1027/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_127 gnd vdd FILL
XFILL_1_DFFPOSX1_948 gnd vdd FILL
XFILL_0_OAI21X1_105 gnd vdd FILL
XFILL_1_DFFPOSX1_937 gnd vdd FILL
XFILL_0_OAI21X1_116 gnd vdd FILL
XFILL_1_OAI21X1_1369 gnd vdd FILL
XFILL_1_OAI21X1_1358 gnd vdd FILL
XFILL_1_DFFPOSX1_926 gnd vdd FILL
XFILL_0_OAI21X1_138 gnd vdd FILL
XFILL_0_OAI21X1_149 gnd vdd FILL
XFILL_1_OAI21X1_309 gnd vdd FILL
XFILL_1_DFFPOSX1_959 gnd vdd FILL
XFILL_6_DFFPOSX1_585 gnd vdd FILL
XFILL_6_DFFPOSX1_596 gnd vdd FILL
XFILL_37_6_0 gnd vdd FILL
XFILL_0_BUFX4_26 gnd vdd FILL
XFILL_0_BUFX4_15 gnd vdd FILL
XFILL_0_NAND2X1_100 gnd vdd FILL
XFILL_1_NAND2X1_304 gnd vdd FILL
XFILL_0_NAND2X1_122 gnd vdd FILL
XFILL_0_BUFX4_48 gnd vdd FILL
XFILL_0_NAND2X1_111 gnd vdd FILL
XFILL_0_BUFX4_59 gnd vdd FILL
XFILL_0_BUFX4_37 gnd vdd FILL
XFILL_0_NAND2X1_133 gnd vdd FILL
XFILL_1_NAND2X1_348 gnd vdd FILL
XFILL_0_NAND2X1_144 gnd vdd FILL
XFILL_0_DFFPOSX1_505 gnd vdd FILL
XFILL_0_NAND2X1_155 gnd vdd FILL
XFILL_0_NAND2X1_166 gnd vdd FILL
XFILL_0_NAND2X1_177 gnd vdd FILL
XFILL_0_INVX1_191 gnd vdd FILL
XFILL_0_DFFPOSX1_516 gnd vdd FILL
XFILL_0_DFFPOSX1_527 gnd vdd FILL
XFILL_0_DFFPOSX1_538 gnd vdd FILL
XFILL_0_NAND2X1_199 gnd vdd FILL
XFILL_0_INVX1_180 gnd vdd FILL
XFILL_1_NAND2X1_359 gnd vdd FILL
XFILL_0_DFFPOSX1_549 gnd vdd FILL
XFILL_0_NAND2X1_188 gnd vdd FILL
XFILL_5_DFFPOSX1_120 gnd vdd FILL
XFILL_5_DFFPOSX1_153 gnd vdd FILL
XFILL_5_DFFPOSX1_131 gnd vdd FILL
XFILL_20_5_0 gnd vdd FILL
XFILL_5_DFFPOSX1_142 gnd vdd FILL
XFILL_5_DFFPOSX1_175 gnd vdd FILL
XFILL_5_DFFPOSX1_164 gnd vdd FILL
XFILL_5_DFFPOSX1_186 gnd vdd FILL
XFILL_24_12_1 gnd vdd FILL
XFILL_5_DFFPOSX1_197 gnd vdd FILL
XOAI21X1_1650 BUFX4_11/A BUFX4_332/Y BUFX2_725/A gnd OAI21X1_1651/C vdd OAI21X1
XOAI21X1_1661 BUFX4_168/Y INVX2_124/Y OAI21X1_1661/C gnd DFFPOSX1_43/D vdd OAI21X1
XOAI21X1_1683 BUFX4_125/Y INVX2_135/Y OAI21X1_1683/C gnd DFFPOSX1_54/D vdd OAI21X1
XOAI21X1_1672 BUFX4_95/Y BUFX4_324/Y BUFX2_718/A gnd OAI21X1_1673/C vdd OAI21X1
XOAI21X1_1694 BUFX4_110/Y BUFX4_359/Y BUFX2_730/A gnd OAI21X1_1695/C vdd OAI21X1
XFILL_0_OAI21X1_650 gnd vdd FILL
XFILL_1_OAI21X1_810 gnd vdd FILL
XFILL_1_OAI21X1_821 gnd vdd FILL
XFILL_0_OR2X2_18 gnd vdd FILL
XFILL_1_OAI21X1_832 gnd vdd FILL
XFILL_1_OAI21X1_843 gnd vdd FILL
XFILL_1_OAI21X1_854 gnd vdd FILL
XFILL_0_OAI21X1_683 gnd vdd FILL
XFILL_0_OAI21X1_672 gnd vdd FILL
XFILL_0_OAI21X1_661 gnd vdd FILL
XNAND3X1_26 INVX4_28/A NOR2X1_99/Y NOR2X1_97/Y gnd OR2X2_14/A vdd NAND3X1
XNAND3X1_37 bundleStartMajId_i[3] INVX4_28/A NOR3X1_10/Y gnd NOR2X1_120/B vdd NAND3X1
XFILL_1_OAI21X1_876 gnd vdd FILL
XFILL_0_OAI21X1_694 gnd vdd FILL
XNAND3X1_48 bundleAddress_i[9] INVX4_48/A AND2X2_24/Y gnd NAND3X1_48/Y vdd NAND3X1
XFILL_1_OAI21X1_887 gnd vdd FILL
XFILL_1_OAI21X1_865 gnd vdd FILL
XNAND3X1_15 bundleStartMajId_i[48] bundleStartMajId_i[47] AND2X2_12/Y gnd NOR2X1_62/B
+ vdd NAND3X1
XFILL_1_OAI21X1_898 gnd vdd FILL
XNAND3X1_59 AND2X2_33/Y AND2X2_26/Y INVX1_210/Y gnd NOR2X1_211/B vdd NAND3X1
XFILL_3_DFFPOSX1_13 gnd vdd FILL
XBUFX2_719 BUFX2_719/A gnd pid3_o[17] vdd BUFX2
XFILL_28_6_0 gnd vdd FILL
XFILL_3_DFFPOSX1_24 gnd vdd FILL
XBUFX2_708 BUFX2_708/A gnd pid2_o[26] vdd BUFX2
XNOR2X1_37 bundleStartMajId_i[21] NOR2X1_37/B gnd NOR2X1_37/Y vdd NOR2X1
XFILL_3_6_0 gnd vdd FILL
XFILL_3_DFFPOSX1_35 gnd vdd FILL
XNOR2X1_26 INVX2_43/Y INVX1_16/Y gnd NOR2X1_26/Y vdd NOR2X1
XNOR2X1_15 INVX2_20/Y INVX4_8/Y gnd AND2X2_3/B vdd NOR2X1
XFILL_3_DFFPOSX1_68 gnd vdd FILL
XFILL_3_DFFPOSX1_57 gnd vdd FILL
XFILL_3_DFFPOSX1_46 gnd vdd FILL
XNOR2X1_48 INVX4_24/Y INVX1_3/Y gnd INVX2_46/A vdd NOR2X1
XNOR2X1_59 INVX1_24/A NOR2X1_59/B gnd NOR2X1_59/Y vdd NOR2X1
XFILL_3_DFFPOSX1_79 gnd vdd FILL
XFILL_0_OAI21X1_1460 gnd vdd FILL
XFILL_29_11_1 gnd vdd FILL
XFILL_0_OAI21X1_1471 gnd vdd FILL
XFILL_0_OAI21X1_1482 gnd vdd FILL
XFILL_0_OAI21X1_1493 gnd vdd FILL
XFILL_11_5_0 gnd vdd FILL
XFILL_0_BUFX2_2 gnd vdd FILL
XFILL_0_BUFX2_404 gnd vdd FILL
XFILL_0_BUFX2_448 gnd vdd FILL
XFILL_0_BUFX2_437 gnd vdd FILL
XFILL_0_BUFX2_426 gnd vdd FILL
XFILL_0_BUFX2_415 gnd vdd FILL
XFILL_0_BUFX2_459 gnd vdd FILL
XFILL_19_6_0 gnd vdd FILL
XFILL_2_OAI21X1_1510 gnd vdd FILL
XFILL_0_NAND2X1_13 gnd vdd FILL
XFILL_4_12_1 gnd vdd FILL
XFILL_0_NAND2X1_35 gnd vdd FILL
XFILL_0_NAND2X1_46 gnd vdd FILL
XFILL_0_NAND2X1_24 gnd vdd FILL
XNOR2X1_105 NOR2X1_105/A NOR2X1_11/B gnd NOR2X1_105/Y vdd NOR2X1
XFILL_2_OAI21X1_1598 gnd vdd FILL
XNOR2X1_127 NOR2X1_216/A NOR2X1_127/B gnd INVX2_94/A vdd NOR2X1
XNOR2X1_149 bundleAddress_i[31] NOR2X1_149/B gnd NOR2X1_149/Y vdd NOR2X1
XFILL_0_NAND2X1_57 gnd vdd FILL
XNOR2X1_116 INVX1_43/Y XNOR2X1_55/A gnd NOR2X1_117/B vdd NOR2X1
XFILL_0_NAND2X1_68 gnd vdd FILL
XFILL_0_NAND2X1_79 gnd vdd FILL
XNOR2X1_138 bundleAddress_i[42] NOR2X1_138/B gnd NOR2X1_138/Y vdd NOR2X1
XFILL_0_INVX2_2 gnd vdd FILL
XFILL_16_3 gnd vdd FILL
XFILL_1_OAI21X1_1111 gnd vdd FILL
XFILL_1_OAI21X1_1100 gnd vdd FILL
XFILL_1_OAI21X1_1122 gnd vdd FILL
XDFFPOSX1_503 BUFX2_532/A CLKBUF1_88/Y OAI21X1_556/Y gnd vdd DFFPOSX1
XDFFPOSX1_514 BUFX2_545/A CLKBUF1_63/Y OAI21X1_581/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_701 gnd vdd FILL
XFILL_1_OAI21X1_1155 gnd vdd FILL
XFILL_1_OAI21X1_1144 gnd vdd FILL
XDFFPOSX1_547 BUFX2_581/A CLKBUF1_29/Y AOI21X1_28/Y gnd vdd DFFPOSX1
XDFFPOSX1_525 BUFX2_557/A CLKBUF1_91/Y OAI21X1_606/Y gnd vdd DFFPOSX1
XDFFPOSX1_536 BUFX2_569/A CLKBUF1_100/Y OAI21X1_633/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_712 gnd vdd FILL
XFILL_1_DFFPOSX1_723 gnd vdd FILL
XFILL_0_BUFX2_960 gnd vdd FILL
XFILL_1_OAI21X1_1133 gnd vdd FILL
XFILL_0_BUFX2_993 gnd vdd FILL
XFILL_1_OAI21X1_106 gnd vdd FILL
XFILL_1_DFFPOSX1_756 gnd vdd FILL
XFILL_0_BUFX2_982 gnd vdd FILL
XFILL_1_OAI21X1_1177 gnd vdd FILL
XFILL_1_OAI21X1_117 gnd vdd FILL
XFILL_1_DFFPOSX1_745 gnd vdd FILL
XFILL_1_OAI21X1_1199 gnd vdd FILL
XFILL_1_DFFPOSX1_734 gnd vdd FILL
XDFFPOSX1_569 BUFX2_599/A CLKBUF1_24/Y OAI21X1_720/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1188 gnd vdd FILL
XFILL_1_DFFPOSX1_767 gnd vdd FILL
XFILL_1_OAI21X1_1166 gnd vdd FILL
XDFFPOSX1_558 BUFX2_587/A CLKBUF1_46/Y OAI21X1_688/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_971 gnd vdd FILL
XFILL_1_OAI21X1_139 gnd vdd FILL
XFILL_1_DFFPOSX1_789 gnd vdd FILL
XNAND2X1_617 bundleAddress_i[18] bundleAddress_i[17] gnd NOR2X1_204/B vdd NAND2X1
XNAND2X1_606 INVX1_207/Y NOR2X1_193/Y gnd NAND2X1_606/Y vdd NAND2X1
XFILL_1_DFFPOSX1_778 gnd vdd FILL
XFILL_1_OAI21X1_128 gnd vdd FILL
XNAND2X1_628 NAND2X1_628/A NOR2X1_222/B gnd NAND2X1_628/Y vdd NAND2X1
XNAND2X1_639 NAND2X1_639/A INVX2_110/Y gnd NAND2X1_639/Y vdd NAND2X1
XINVX1_18 NOR3X1_3/C gnd INVX1_18/Y vdd INVX1
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XFILL_6_DFFPOSX1_360 gnd vdd FILL
XFILL_6_DFFPOSX1_371 gnd vdd FILL
XFILL_9_11_1 gnd vdd FILL
XFILL_6_DFFPOSX1_382 gnd vdd FILL
XFILL_6_DFFPOSX1_393 gnd vdd FILL
XNAND2X1_70 BUFX2_900/A BUFX4_217/Y gnd OAI21X1_70/C vdd NAND2X1
XNAND2X1_81 BUFX2_456/A BUFX4_387/Y gnd NAND2X1_81/Y vdd NAND2X1
XNAND2X1_92 BUFX2_406/A BUFX4_383/Y gnd NAND2X1_92/Y vdd NAND2X1
XFILL_1_NAND2X1_112 gnd vdd FILL
XFILL_10_18_1 gnd vdd FILL
XFILL_1_NAND2X1_101 gnd vdd FILL
XFILL_0_XNOR2X1_103 gnd vdd FILL
XFILL_1_NAND2X1_134 gnd vdd FILL
XFILL_0_DFFPOSX1_313 gnd vdd FILL
XFILL_0_DFFPOSX1_302 gnd vdd FILL
XFILL_0_DFFPOSX1_324 gnd vdd FILL
XFILL_0_DFFPOSX1_346 gnd vdd FILL
XFILL_0_DFFPOSX1_335 gnd vdd FILL
XFILL_1_NAND2X1_189 gnd vdd FILL
XFILL_0_DFFPOSX1_357 gnd vdd FILL
XFILL_1_NAND2X1_178 gnd vdd FILL
XFILL_1_NAND2X1_167 gnd vdd FILL
XFILL_0_DFFPOSX1_368 gnd vdd FILL
XFILL_0_DFFPOSX1_379 gnd vdd FILL
XFILL_3_DFFPOSX1_839 gnd vdd FILL
XFILL_3_DFFPOSX1_806 gnd vdd FILL
XFILL_3_DFFPOSX1_817 gnd vdd FILL
XFILL_3_DFFPOSX1_828 gnd vdd FILL
XOAI21X1_1480 BUFX4_170/Y BUFX4_35/Y BUFX2_220/A gnd OAI21X1_1482/C vdd OAI21X1
XOAI21X1_1491 BUFX4_160/Y BUFX4_66/A BUFX2_223/A gnd OAI21X1_1492/C vdd OAI21X1
XFILL_1_NOR2X1_212 gnd vdd FILL
XFILL_1_NOR2X1_201 gnd vdd FILL
XFILL_1_OAI21X1_651 gnd vdd FILL
XFILL_0_OAI21X1_491 gnd vdd FILL
XFILL_1_OAI21X1_640 gnd vdd FILL
XFILL_3_NOR3X1_2 gnd vdd FILL
XFILL_1_OAI21X1_662 gnd vdd FILL
XFILL_0_OAI21X1_480 gnd vdd FILL
XFILL_2_OAI21X1_855 gnd vdd FILL
XFILL_1_OAI21X1_695 gnd vdd FILL
XFILL_1_OAI21X1_684 gnd vdd FILL
XFILL_1_OAI21X1_673 gnd vdd FILL
XFILL_15_17_1 gnd vdd FILL
XBUFX2_516 BUFX2_516/A gnd majID2_o[1] vdd BUFX2
XFILL_4_DFFPOSX1_14 gnd vdd FILL
XFILL_2_DFFPOSX1_418 gnd vdd FILL
XFILL_2_DFFPOSX1_407 gnd vdd FILL
XBUFX2_505 BUFX2_505/A gnd majID2_o[11] vdd BUFX2
XBUFX2_527 BUFX2_527/A gnd majID3_o[49] vdd BUFX2
XFILL_2_DFFPOSX1_429 gnd vdd FILL
XFILL_4_DFFPOSX1_36 gnd vdd FILL
XFILL_4_DFFPOSX1_47 gnd vdd FILL
XFILL_4_DFFPOSX1_25 gnd vdd FILL
XBUFX2_538 BUFX2_538/A gnd majID3_o[39] vdd BUFX2
XBUFX2_549 BUFX2_549/A gnd majID3_o[29] vdd BUFX2
XFILL_4_DFFPOSX1_69 gnd vdd FILL
XFILL_4_DFFPOSX1_58 gnd vdd FILL
XFILL_1_NAND2X1_690 gnd vdd FILL
XFILL_0_OAI21X1_1290 gnd vdd FILL
XFILL_0_DFFPOSX1_880 gnd vdd FILL
XFILL_0_DFFPOSX1_891 gnd vdd FILL
XDFFPOSX1_1010 BUFX2_677/A CLKBUF1_41/Y OAI21X1_1587/Y gnd vdd DFFPOSX1
XDFFPOSX1_1032 BUFX2_670/A CLKBUF1_101/Y OAI21X1_1609/Y gnd vdd DFFPOSX1
XDFFPOSX1_1021 BUFX2_658/A CLKBUF1_95/Y OAI21X1_1598/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_201 gnd vdd FILL
XFILL_0_BUFX2_212 gnd vdd FILL
XFILL_0_BUFX2_223 gnd vdd FILL
XFILL_0_BUFX2_234 gnd vdd FILL
XFILL_0_BUFX2_256 gnd vdd FILL
XFILL_0_BUFX2_245 gnd vdd FILL
XFILL_0_BUFX2_278 gnd vdd FILL
XFILL_0_BUFX2_267 gnd vdd FILL
XFILL_0_BUFX2_289 gnd vdd FILL
XFILL_33_18_1 gnd vdd FILL
XFILL_14_12_0 gnd vdd FILL
XFILL_35_9_1 gnd vdd FILL
XFILL_2_DFFPOSX1_941 gnd vdd FILL
XFILL_2_OAI21X1_1373 gnd vdd FILL
XFILL_2_DFFPOSX1_930 gnd vdd FILL
XFILL_2_OAI21X1_1362 gnd vdd FILL
XFILL_34_4_0 gnd vdd FILL
XFILL_2_DFFPOSX1_952 gnd vdd FILL
XFILL_2_DFFPOSX1_985 gnd vdd FILL
XFILL_2_DFFPOSX1_963 gnd vdd FILL
XFILL_2_DFFPOSX1_974 gnd vdd FILL
XFILL_21_1 gnd vdd FILL
XFILL_2_DFFPOSX1_996 gnd vdd FILL
XFILL_0_NAND3X1_8 gnd vdd FILL
XOAI21X1_419 OAI21X1_419/A BUFX4_181/Y OAI21X1_419/C gnd OAI21X1_419/Y vdd OAI21X1
XOAI21X1_408 INVX1_8/A NOR2X1_60/A INVX2_13/Y gnd OAI21X1_408/Y vdd OAI21X1
XFILL_3_XNOR2X1_21 gnd vdd FILL
XFILL_3_XNOR2X1_32 gnd vdd FILL
XFILL_3_XNOR2X1_10 gnd vdd FILL
XDFFPOSX1_322 BUFX2_993/A CLKBUF1_102/Y OAI21X1_261/Y gnd vdd DFFPOSX1
XDFFPOSX1_311 BUFX2_980/A CLKBUF1_72/Y OAI21X1_239/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_65 gnd vdd FILL
XFILL_3_XNOR2X1_43 gnd vdd FILL
XFILL_3_XNOR2X1_54 gnd vdd FILL
XDFFPOSX1_300 BUFX2_1031/A CLKBUF1_4/Y OAI21X1_217/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_76 gnd vdd FILL
XFILL_1_DFFPOSX1_542 gnd vdd FILL
XDFFPOSX1_333 BUFX2_1005/A CLKBUF1_21/Y OAI21X1_283/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_98 gnd vdd FILL
XFILL_1_DFFPOSX1_520 gnd vdd FILL
XFILL_1_DFFPOSX1_531 gnd vdd FILL
XFILL_3_XNOR2X1_87 gnd vdd FILL
XDFFPOSX1_355 BUFX2_1029/A CLKBUF1_58/Y OAI21X1_327/Y gnd vdd DFFPOSX1
XDFFPOSX1_344 BUFX2_1017/A CLKBUF1_15/Y OAI21X1_305/Y gnd vdd DFFPOSX1
XFILL_38_17_1 gnd vdd FILL
XFILL_1_DFFPOSX1_575 gnd vdd FILL
XDFFPOSX1_388 BUFX2_419/A CLKBUF1_79/Y OAI21X1_360/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_564 gnd vdd FILL
XFILL_0_BUFX2_790 gnd vdd FILL
XDFFPOSX1_377 BUFX2_407/A CLKBUF1_18/Y OAI21X1_349/Y gnd vdd DFFPOSX1
XDFFPOSX1_366 BUFX2_395/A CLKBUF1_75/Y OAI21X1_338/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_553 gnd vdd FILL
XNAND2X1_414 BUFX2_5/A BUFX4_386/Y gnd NAND2X1_414/Y vdd NAND2X1
XDFFPOSX1_399 BUFX2_431/A CLKBUF1_100/Y OAI21X1_371/Y gnd vdd DFFPOSX1
XNAND2X1_403 BUFX2_2/A BUFX4_376/Y gnd NAND2X1_403/Y vdd NAND2X1
XFILL_19_11_0 gnd vdd FILL
XNAND2X1_436 BUFX2_29/A BUFX4_324/Y gnd NAND2X1_436/Y vdd NAND2X1
XFILL_1_DFFPOSX1_586 gnd vdd FILL
XFILL_1_DFFPOSX1_597 gnd vdd FILL
XFILL_2_OAI21X1_129 gnd vdd FILL
XNAND2X1_425 BUFX2_17/A BUFX4_326/Y gnd NAND2X1_425/Y vdd NAND2X1
XNAND2X1_469 BUFX4_238/Y NOR2X1_123/Y gnd NAND2X1_469/Y vdd NAND2X1
XNAND2X1_447 BUFX2_41/A BUFX4_381/Y gnd NAND2X1_447/Y vdd NAND2X1
XNAND2X1_458 BUFX2_53/A BUFX4_343/Y gnd NAND2X1_458/Y vdd NAND2X1
XFILL_32_13_0 gnd vdd FILL
XFILL_26_9_1 gnd vdd FILL
XFILL_25_4_0 gnd vdd FILL
XFILL_1_9_1 gnd vdd FILL
XFILL_0_4_0 gnd vdd FILL
XFILL_0_DFFPOSX1_121 gnd vdd FILL
XFILL_1_XNOR2X1_104 gnd vdd FILL
XFILL_0_DFFPOSX1_110 gnd vdd FILL
XFILL_0_DFFPOSX1_132 gnd vdd FILL
XFILL_0_DFFPOSX1_154 gnd vdd FILL
XFILL_0_DFFPOSX1_143 gnd vdd FILL
XFILL_1_BUFX2_903 gnd vdd FILL
XFILL_0_DFFPOSX1_165 gnd vdd FILL
XFILL_0_DFFPOSX1_198 gnd vdd FILL
XFILL_1_BUFX2_947 gnd vdd FILL
XFILL_1_BUFX2_925 gnd vdd FILL
XFILL_1_BUFX2_936 gnd vdd FILL
XFILL_0_DFFPOSX1_176 gnd vdd FILL
XFILL_0_DFFPOSX1_187 gnd vdd FILL
XOAI21X1_931 BUFX4_123/Y INVX1_120/Y OAI21X1_931/C gnd OAI21X1_931/Y vdd OAI21X1
XFILL_4_CLKBUF1_100 gnd vdd FILL
XFILL_3_DFFPOSX1_603 gnd vdd FILL
XOAI21X1_942 BUFX4_104/Y BUFX4_326/Y BUFX2_334/A gnd OAI21X1_943/C vdd OAI21X1
XOAI21X1_920 BUFX4_6/Y OAI21X1_7/A BUFX2_353/A gnd OAI21X1_921/C vdd OAI21X1
XOAI21X1_975 BUFX4_293/Y INVX1_142/Y OAI21X1_975/C gnd OAI21X1_975/Y vdd OAI21X1
XFILL_3_DFFPOSX1_636 gnd vdd FILL
XOAI21X1_953 BUFX4_141/Y INVX1_131/Y OAI21X1_953/C gnd OAI21X1_953/Y vdd OAI21X1
XOAI21X1_964 BUFX4_10/A BUFX4_335/Y BUFX2_346/A gnd OAI21X1_965/C vdd OAI21X1
XFILL_3_DFFPOSX1_647 gnd vdd FILL
XFILL_3_DFFPOSX1_625 gnd vdd FILL
XFILL_3_DFFPOSX1_614 gnd vdd FILL
XFILL_3_DFFPOSX1_658 gnd vdd FILL
XFILL_3_DFFPOSX1_669 gnd vdd FILL
XOAI21X1_986 BUFX4_158/Y BUFX4_28/Y BUFX2_386/A gnd OAI21X1_987/C vdd OAI21X1
XOAI21X1_997 BUFX4_303/Y INVX1_153/Y OAI21X1_997/C gnd OAI21X1_997/Y vdd OAI21X1
XFILL_37_12_0 gnd vdd FILL
XFILL_8_5_0 gnd vdd FILL
XINVX2_61 bundleAddress_i[55] gnd INVX2_61/Y vdd INVX2
XINVX2_72 bundleAddress_i[36] gnd INVX2_72/Y vdd INVX2
XINVX2_50 INVX2_50/A gnd INVX2_50/Y vdd INVX2
XFILL_1_OAI21X1_481 gnd vdd FILL
XFILL_1_OAI21X1_470 gnd vdd FILL
XINVX2_94 INVX2_94/A gnd INVX2_94/Y vdd INVX2
XFILL_1_OAI21X1_492 gnd vdd FILL
XINVX2_83 bundleAddress_i[14] gnd INVX2_83/Y vdd INVX2
XFILL_0_AOI21X1_2 gnd vdd FILL
XFILL_2_OAI21X1_696 gnd vdd FILL
XFILL_2_DFFPOSX1_204 gnd vdd FILL
XBUFX2_302 BUFX2_302/A gnd instr2_o[14] vdd BUFX2
XFILL_2_DFFPOSX1_237 gnd vdd FILL
XBUFX2_335 BUFX2_335/A gnd instr3_o[13] vdd BUFX2
XFILL_2_DFFPOSX1_215 gnd vdd FILL
XFILL_2_DFFPOSX1_226 gnd vdd FILL
XBUFX2_313 BUFX2_313/A gnd instr2_o[4] vdd BUFX2
XBUFX2_324 BUFX2_324/A gnd instr2_o[22] vdd BUFX2
XFILL_5_DFFPOSX1_37 gnd vdd FILL
XFILL_5_DFFPOSX1_26 gnd vdd FILL
XFILL_2_DFFPOSX1_248 gnd vdd FILL
XFILL_5_DFFPOSX1_15 gnd vdd FILL
XFILL_2_DFFPOSX1_259 gnd vdd FILL
XFILL_17_9_1 gnd vdd FILL
XFILL_16_4_0 gnd vdd FILL
XBUFX2_368 BUFX2_368/A gnd instr4_o[12] vdd BUFX2
XBUFX2_357 BUFX2_357/A gnd instr4_o[31] vdd BUFX2
XBUFX2_346 BUFX2_346/A gnd instr3_o[3] vdd BUFX2
XBUFX2_379 BUFX2_379/A gnd instr4_o[2] vdd BUFX2
XFILL_5_DFFPOSX1_59 gnd vdd FILL
XFILL_1_INVX4_50 gnd vdd FILL
XFILL_5_DFFPOSX1_48 gnd vdd FILL
XOAI21X1_35 INVX2_173/Y BUFX4_234/Y OAI21X1_35/C gnd OAI21X1_35/Y vdd OAI21X1
XOAI21X1_24 INVX2_162/Y BUFX4_223/Y OAI21X1_24/C gnd OAI21X1_24/Y vdd OAI21X1
XFILL_1_NOR3X1_18 gnd vdd FILL
XFILL_1_BUFX4_240 gnd vdd FILL
XFILL_5_DFFPOSX1_719 gnd vdd FILL
XFILL_5_DFFPOSX1_708 gnd vdd FILL
XOAI21X1_13 INVX2_151/Y BUFX4_196/Y OAI21X1_13/C gnd OAI21X1_13/Y vdd OAI21X1
XOAI21X1_46 INVX2_184/Y BUFX4_227/Y OAI21X1_46/C gnd OAI21X1_46/Y vdd OAI21X1
XFILL_1_BUFX4_251 gnd vdd FILL
XFILL_1_BUFX4_273 gnd vdd FILL
XOAI21X1_57 INVX2_195/Y BUFX4_195/Y OAI21X1_57/C gnd OAI21X1_57/Y vdd OAI21X1
XFILL_1_BUFX4_262 gnd vdd FILL
XOAI21X1_68 INVX2_4/Y BUFX4_186/Y OAI21X1_68/C gnd OAI21X1_68/Y vdd OAI21X1
XFILL_1_BUFX4_295 gnd vdd FILL
XFILL_1_BUFX4_284 gnd vdd FILL
XOAI21X1_79 BUFX4_135/Y INVX2_149/Y OAI21X1_79/C gnd OAI21X1_79/Y vdd OAI21X1
XFILL_0_DFFPOSX1_11 gnd vdd FILL
XFILL_4_DFFPOSX1_309 gnd vdd FILL
XFILL_0_DFFPOSX1_44 gnd vdd FILL
XFILL_0_DFFPOSX1_22 gnd vdd FILL
XFILL_0_DFFPOSX1_33 gnd vdd FILL
XFILL_0_DFFPOSX1_77 gnd vdd FILL
XFILL_0_DFFPOSX1_55 gnd vdd FILL
XFILL_0_DFFPOSX1_66 gnd vdd FILL
XFILL_0_DFFPOSX1_88 gnd vdd FILL
XFILL_0_DFFPOSX1_99 gnd vdd FILL
XFILL_2_DFFPOSX1_760 gnd vdd FILL
XFILL_2_OAI21X1_1181 gnd vdd FILL
XFILL_2_OAI21X1_1192 gnd vdd FILL
XBUFX2_880 BUFX2_880/A gnd tid2_o[19] vdd BUFX2
XBUFX2_891 BUFX2_891/A gnd tid2_o[9] vdd BUFX2
XFILL_2_DFFPOSX1_771 gnd vdd FILL
XFILL_2_DFFPOSX1_793 gnd vdd FILL
XFILL_2_DFFPOSX1_782 gnd vdd FILL
XFILL_0_NOR2X1_220 gnd vdd FILL
XFILL_0_NOR2X1_231 gnd vdd FILL
XOAI21X1_238 BUFX4_161/Y BUFX4_63/Y BUFX2_980/A gnd OAI21X1_239/C vdd OAI21X1
XOAI21X1_216 BUFX4_135/Y BUFX4_49/Y BUFX2_1031/A gnd OAI21X1_217/C vdd OAI21X1
XOAI21X1_205 INVX2_148/Y BUFX4_300/Y OAI21X1_205/C gnd OAI21X1_205/Y vdd OAI21X1
XOAI21X1_227 INVX2_159/Y BUFX4_302/Y OAI21X1_227/C gnd OAI21X1_227/Y vdd OAI21X1
XFILL_6_DFFPOSX1_7 gnd vdd FILL
XOAI21X1_249 INVX2_170/Y BUFX4_291/Y OAI21X1_249/C gnd OAI21X1_249/Y vdd OAI21X1
XFILL_21_10_1 gnd vdd FILL
XDFFPOSX1_130 BUFX2_801/A CLKBUF1_93/Y OAI21X1_1804/Y gnd vdd DFFPOSX1
XAND2X2_16 NOR2X1_97/Y INVX1_43/A gnd NOR2X1_98/B vdd AND2X2
XAND2X2_27 AND2X2_27/A INVX4_37/Y gnd AND2X2_27/Y vdd AND2X2
XDFFPOSX1_163 NAND2X1_7/A CLKBUF1_38/Y OAI21X1_7/Y gnd vdd DFFPOSX1
XDFFPOSX1_152 BUFX2_825/A CLKBUF1_15/Y OAI21X1_1826/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_350 gnd vdd FILL
XDFFPOSX1_141 BUFX2_813/A CLKBUF1_81/Y OAI21X1_1815/Y gnd vdd DFFPOSX1
XDFFPOSX1_185 BUFX2_855/A CLKBUF1_64/Y OAI21X1_29/Y gnd vdd DFFPOSX1
XNAND2X1_200 BUFX2_481/A BUFX4_209/Y gnd OAI21X1_445/C vdd NAND2X1
XNAND2X1_211 BUFX2_488/A BUFX4_221/Y gnd OAI21X1_455/C vdd NAND2X1
XFILL_0_NOR3X1_6 gnd vdd FILL
XDFFPOSX1_196 BUFX2_867/A CLKBUF1_6/Y OAI21X1_40/Y gnd vdd DFFPOSX1
XDFFPOSX1_174 BUFX2_843/A CLKBUF1_51/Y OAI21X1_18/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_361 gnd vdd FILL
XFILL_1_DFFPOSX1_372 gnd vdd FILL
XFILL_1_DFFPOSX1_383 gnd vdd FILL
XFILL_1_DFFPOSX1_394 gnd vdd FILL
XNAND2X1_222 BUFX2_494/A BUFX4_204/Y gnd OAI21X1_463/C vdd NAND2X1
XNAND2X1_233 INVX1_18/Y NOR2X1_41/Y gnd NOR2X1_42/B vdd NAND2X1
XNAND2X1_244 bundleStartMajId_i[11] NOR2X1_47/Y gnd INVX1_20/A vdd NAND2X1
XFILL_4_DFFPOSX1_821 gnd vdd FILL
XFILL_4_DFFPOSX1_810 gnd vdd FILL
XNAND2X1_255 BUFX2_510/A BUFX4_221/Y gnd OAI21X1_489/C vdd NAND2X1
XNAND2X1_266 INVX2_8/Y INVX2_9/Y gnd OAI21X1_663/A vdd NAND2X1
XNAND2X1_277 AND2X2_3/B NOR2X1_64/B gnd MUX2X1_1/A vdd NAND2X1
XFILL_4_DFFPOSX1_832 gnd vdd FILL
XNAND2X1_299 INVX2_51/A NOR2X1_51/Y gnd OR2X2_13/B vdd NAND2X1
XFILL_4_DFFPOSX1_854 gnd vdd FILL
XNAND2X1_288 NOR2X1_67/Y NOR2X1_74/Y gnd NOR2X1_76/B vdd NAND2X1
XFILL_4_DFFPOSX1_843 gnd vdd FILL
XFILL_4_DFFPOSX1_865 gnd vdd FILL
XFILL_4_DFFPOSX1_887 gnd vdd FILL
XFILL_4_DFFPOSX1_876 gnd vdd FILL
XFILL_4_DFFPOSX1_898 gnd vdd FILL
XFILL_0_OAI21X1_5 gnd vdd FILL
XFILL_0_BUFX2_70 gnd vdd FILL
XFILL_1_BUFX2_700 gnd vdd FILL
XFILL_0_BUFX2_81 gnd vdd FILL
XFILL_0_BUFX2_92 gnd vdd FILL
XFILL_1_BUFX2_733 gnd vdd FILL
XFILL_1_BUFX2_744 gnd vdd FILL
XFILL_0_BUFX4_307 gnd vdd FILL
XFILL_1_NOR2X1_40 gnd vdd FILL
XFILL_1_BUFX2_788 gnd vdd FILL
XFILL_0_BUFX4_329 gnd vdd FILL
XFILL_1_BUFX2_777 gnd vdd FILL
XFILL_0_BUFX4_318 gnd vdd FILL
XFILL_23_18_0 gnd vdd FILL
XOAI21X1_750 OAI21X1_750/A BUFX4_299/Y OAI21X1_750/C gnd OAI21X1_750/Y vdd OAI21X1
XFILL_1_NOR2X1_84 gnd vdd FILL
XFILL_3_DFFPOSX1_422 gnd vdd FILL
XFILL_3_DFFPOSX1_400 gnd vdd FILL
XFILL_3_DFFPOSX1_411 gnd vdd FILL
XOAI21X1_772 OAI21X1_772/A BUFX4_300/Y OAI21X1_772/C gnd OAI21X1_772/Y vdd OAI21X1
XOAI21X1_761 INVX2_48/Y OR2X2_15/Y OAI21X1_761/C gnd OAI21X1_763/A vdd OAI21X1
XOAI21X1_794 NOR3X1_9/B OR2X2_15/A OAI21X1_794/C gnd OAI21X1_796/A vdd OAI21X1
XOAI21X1_783 NOR2X1_114/B NOR3X1_2/B NOR3X1_2/A gnd OAI21X1_784/C vdd OAI21X1
XFILL_1_BUFX2_799 gnd vdd FILL
XFILL_3_DFFPOSX1_433 gnd vdd FILL
XFILL_3_DFFPOSX1_455 gnd vdd FILL
XFILL_3_DFFPOSX1_444 gnd vdd FILL
XFILL_3_DFFPOSX1_477 gnd vdd FILL
XFILL_3_DFFPOSX1_466 gnd vdd FILL
XFILL_3_DFFPOSX1_488 gnd vdd FILL
XFILL_3_DFFPOSX1_499 gnd vdd FILL
XFILL_6_DFFPOSX1_904 gnd vdd FILL
XFILL_6_DFFPOSX1_915 gnd vdd FILL
XFILL_6_DFFPOSX1_926 gnd vdd FILL
XFILL_2_OAI21X1_482 gnd vdd FILL
XBUFX2_110 BUFX2_110/A gnd addr2_o[58] vdd BUFX2
XFILL_2_XNOR2X1_40 gnd vdd FILL
XFILL_0_NAND2X1_507 gnd vdd FILL
XBUFX2_121 BUFX2_121/A gnd addr2_o[57] vdd BUFX2
XBUFX2_132 BUFX2_132/A gnd addr3_o[52] vdd BUFX2
XFILL_0_NAND2X1_529 gnd vdd FILL
XFILL_2_XNOR2X1_73 gnd vdd FILL
XFILL_2_XNOR2X1_62 gnd vdd FILL
XFILL_0_NAND2X1_518 gnd vdd FILL
XFILL_2_XNOR2X1_51 gnd vdd FILL
XBUFX2_143 BUFX2_143/A gnd addr3_o[42] vdd BUFX2
XFILL_1_10_1 gnd vdd FILL
XBUFX2_154 BUFX2_154/A gnd addr3_o[32] vdd BUFX2
XFILL_6_DFFPOSX1_16 gnd vdd FILL
XBUFX2_187 BUFX2_187/A gnd addr3_o[2] vdd BUFX2
XFILL_2_XNOR2X1_95 gnd vdd FILL
XBUFX2_176 BUFX2_176/A gnd addr3_o[12] vdd BUFX2
XBUFX2_165 BUFX2_165/A gnd addr3_o[22] vdd BUFX2
XFILL_2_XNOR2X1_84 gnd vdd FILL
XBUFX2_198 BUFX2_198/A gnd addr4_o[50] vdd BUFX2
XFILL_32_7_1 gnd vdd FILL
XFILL_31_2_0 gnd vdd FILL
XFILL_28_17_0 gnd vdd FILL
XFILL_5_DFFPOSX1_516 gnd vdd FILL
XFILL_5_DFFPOSX1_527 gnd vdd FILL
XFILL_5_DFFPOSX1_505 gnd vdd FILL
XFILL_5_DFFPOSX1_538 gnd vdd FILL
XFILL_5_DFFPOSX1_549 gnd vdd FILL
XBUFX2_1002 BUFX2_1002/A gnd tid4_o[24] vdd BUFX2
XBUFX2_1013 BUFX2_1013/A gnd tid4_o[14] vdd BUFX2
XBUFX2_1024 BUFX2_1024/A gnd tid4_o[4] vdd BUFX2
XCLKBUF1_14 BUFX4_92/Y gnd CLKBUF1_14/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_117 gnd vdd FILL
XCLKBUF1_25 BUFX4_87/Y gnd CLKBUF1_25/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_12 gnd vdd FILL
XCLKBUF1_47 BUFX4_86/Y gnd CLKBUF1_47/Y vdd CLKBUF1
XCLKBUF1_36 BUFX4_92/Y gnd CLKBUF1_36/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_106 gnd vdd FILL
XFILL_1_DFFPOSX1_23 gnd vdd FILL
XFILL_1_DFFPOSX1_45 gnd vdd FILL
XFILL_1_DFFPOSX1_56 gnd vdd FILL
XFILL_4_DFFPOSX1_139 gnd vdd FILL
XCLKBUF1_69 BUFX4_89/Y gnd CLKBUF1_69/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_34 gnd vdd FILL
XFILL_4_DFFPOSX1_128 gnd vdd FILL
XCLKBUF1_58 BUFX4_89/Y gnd CLKBUF1_58/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_78 gnd vdd FILL
XFILL_1_DFFPOSX1_89 gnd vdd FILL
XFILL_3_18_0 gnd vdd FILL
XFILL_1_DFFPOSX1_67 gnd vdd FILL
XFILL_0_OAI21X1_1801 gnd vdd FILL
XBUFX4_90 clock_i gnd BUFX4_90/Y vdd BUFX4
XFILL_0_OAI21X1_1812 gnd vdd FILL
XFILL_0_OAI21X1_1823 gnd vdd FILL
XFILL_23_7_1 gnd vdd FILL
XFILL_2_DFFPOSX1_590 gnd vdd FILL
XFILL_22_2_0 gnd vdd FILL
XFILL_2_AOI21X1_51 gnd vdd FILL
XFILL_1_DFFPOSX1_191 gnd vdd FILL
XFILL_1_DFFPOSX1_180 gnd vdd FILL
XFILL_8_17_0 gnd vdd FILL
XFILL_4_DFFPOSX1_640 gnd vdd FILL
XFILL_5_3_0 gnd vdd FILL
XFILL_6_8_1 gnd vdd FILL
XFILL_4_DFFPOSX1_662 gnd vdd FILL
XFILL_4_DFFPOSX1_651 gnd vdd FILL
XFILL_4_DFFPOSX1_673 gnd vdd FILL
XFILL_4_DFFPOSX1_695 gnd vdd FILL
XFILL_12_15_1 gnd vdd FILL
XFILL_4_DFFPOSX1_684 gnd vdd FILL
XFILL_14_7_1 gnd vdd FILL
XFILL_4_CLKBUF1_9 gnd vdd FILL
XFILL_13_2_0 gnd vdd FILL
XFILL_1_BUFX2_530 gnd vdd FILL
XFILL_0_BUFX4_115 gnd vdd FILL
XFILL_0_BUFX4_104 gnd vdd FILL
XFILL_1_INVX1_51 gnd vdd FILL
XFILL_1_BUFX2_552 gnd vdd FILL
XFILL_1_BUFX2_541 gnd vdd FILL
XFILL_0_BUFX4_137 gnd vdd FILL
XFILL_1_BUFX2_574 gnd vdd FILL
XFILL_0_BUFX4_126 gnd vdd FILL
XFILL_0_BUFX4_148 gnd vdd FILL
XFILL_1_BUFX2_596 gnd vdd FILL
XFILL_1_BUFX2_585 gnd vdd FILL
XFILL_3_DFFPOSX1_230 gnd vdd FILL
XOAI21X1_1309 OAI21X1_1309/A BUFX4_169/Y OAI21X1_1309/C gnd OAI21X1_1309/Y vdd OAI21X1
XFILL_3_DFFPOSX1_252 gnd vdd FILL
XFILL_1_BUFX2_26 gnd vdd FILL
XFILL_0_BUFX4_159 gnd vdd FILL
XFILL_1_OAI21X1_1529 gnd vdd FILL
XFILL_1_OAI21X1_1518 gnd vdd FILL
XFILL_3_DFFPOSX1_263 gnd vdd FILL
XOAI21X1_580 OR2X2_6/Y NOR2X1_74/A INVX8_6/A gnd OAI21X1_581/A vdd OAI21X1
XFILL_1_OAI21X1_1507 gnd vdd FILL
XOAI21X1_591 OR2X2_9/A OR2X2_8/A OR2X2_8/B gnd OAI21X1_592/C vdd OAI21X1
XFILL_3_DFFPOSX1_241 gnd vdd FILL
XFILL_1_BUFX2_15 gnd vdd FILL
XFILL_3_DFFPOSX1_296 gnd vdd FILL
XFILL_3_DFFPOSX1_285 gnd vdd FILL
XFILL_0_OAI21X1_309 gnd vdd FILL
XFILL_3_DFFPOSX1_274 gnd vdd FILL
XFILL_1_BUFX2_37 gnd vdd FILL
XFILL_5_DFFPOSX1_4 gnd vdd FILL
XFILL_17_14_1 gnd vdd FILL
XFILL_6_DFFPOSX1_778 gnd vdd FILL
XFILL_4_3 gnd vdd FILL
XFILL_6_DFFPOSX1_767 gnd vdd FILL
XFILL_6_DFFPOSX1_789 gnd vdd FILL
XFILL_30_16_1 gnd vdd FILL
XFILL_0_NAND2X1_304 gnd vdd FILL
XFILL_0_NAND2X1_326 gnd vdd FILL
XFILL_0_NAND2X1_315 gnd vdd FILL
XFILL_0_OAI21X1_1108 gnd vdd FILL
XFILL_0_NAND2X1_337 gnd vdd FILL
XFILL_0_OAI21X1_1119 gnd vdd FILL
XFILL_11_10_0 gnd vdd FILL
XFILL_0_NAND2X1_348 gnd vdd FILL
XFILL_0_NAND2X1_359 gnd vdd FILL
XFILL_1_NOR2X1_6 gnd vdd FILL
XFILL_39_2 gnd vdd FILL
XFILL_0_DFFPOSX1_709 gnd vdd FILL
XFILL_1_DFFPOSX1_1021 gnd vdd FILL
XFILL_5_DFFPOSX1_302 gnd vdd FILL
XFILL_1_DFFPOSX1_1010 gnd vdd FILL
XFILL_1_DFFPOSX1_1032 gnd vdd FILL
XFILL_5_DFFPOSX1_335 gnd vdd FILL
XFILL_5_DFFPOSX1_313 gnd vdd FILL
XFILL_5_DFFPOSX1_324 gnd vdd FILL
XFILL_5_DFFPOSX1_346 gnd vdd FILL
XFILL_5_DFFPOSX1_357 gnd vdd FILL
XFILL_5_DFFPOSX1_368 gnd vdd FILL
XFILL_5_DFFPOSX1_379 gnd vdd FILL
XOAI21X1_1821 BUFX4_361/Y INVX2_193/Y NAND2X1_762/Y gnd OAI21X1_1821/Y vdd OAI21X1
XOAI21X1_1810 BUFX4_311/Y INVX2_182/Y NAND2X1_751/Y gnd OAI21X1_1810/Y vdd OAI21X1
XFILL_1_NAND2X1_17 gnd vdd FILL
XFILL_1_NAND2X1_39 gnd vdd FILL
XINVX4_18 bundleStartMajId_i[24] gnd INVX4_18/Y vdd INVX4
XINVX4_29 INVX4_29/A gnd INVX4_29/Y vdd INVX4
XFILL_0_OAI21X1_832 gnd vdd FILL
XFILL_0_OAI21X1_810 gnd vdd FILL
XFILL_0_OAI21X1_821 gnd vdd FILL
XFILL_0_OAI21X1_843 gnd vdd FILL
XFILL_0_OAI21X1_854 gnd vdd FILL
XFILL_0_OAI21X1_865 gnd vdd FILL
XFILL_0_OAI21X1_898 gnd vdd FILL
XFILL_0_OAI21X1_876 gnd vdd FILL
XFILL_0_OAI21X1_887 gnd vdd FILL
XFILL_35_15_1 gnd vdd FILL
XFILL_2_DFFPOSX1_13 gnd vdd FILL
XFILL_2_DFFPOSX1_46 gnd vdd FILL
XFILL_2_DFFPOSX1_24 gnd vdd FILL
XFILL_2_DFFPOSX1_35 gnd vdd FILL
XFILL_2_DFFPOSX1_68 gnd vdd FILL
XFILL_2_DFFPOSX1_57 gnd vdd FILL
XFILL_2_DFFPOSX1_79 gnd vdd FILL
XFILL_0_OAI21X1_1642 gnd vdd FILL
XFILL_0_OAI21X1_1631 gnd vdd FILL
XFILL_0_OAI21X1_1620 gnd vdd FILL
XFILL_0_OAI21X1_1675 gnd vdd FILL
XFILL_0_OAI21X1_1653 gnd vdd FILL
XFILL_0_OAI21X1_1664 gnd vdd FILL
XFILL_0_OAI21X1_1686 gnd vdd FILL
XFILL_0_OAI21X1_1697 gnd vdd FILL
XFILL_0_BUFX4_6 gnd vdd FILL
XFILL_5_DFFPOSX1_880 gnd vdd FILL
XFILL_5_DFFPOSX1_891 gnd vdd FILL
XFILL_0_BUFX2_608 gnd vdd FILL
XFILL_0_BUFX2_619 gnd vdd FILL
XFILL_4_DFFPOSX1_1014 gnd vdd FILL
XFILL_1_XNOR2X1_81 gnd vdd FILL
XFILL_4_DFFPOSX1_1003 gnd vdd FILL
XFILL_1_XNOR2X1_70 gnd vdd FILL
XFILL_4_DFFPOSX1_1025 gnd vdd FILL
XFILL_1_XNOR2X1_92 gnd vdd FILL
XFILL_34_10_0 gnd vdd FILL
XBUFX4_216 BUFX4_24/Y gnd BUFX4_216/Y vdd BUFX4
XBUFX4_205 BUFX4_23/Y gnd BUFX4_205/Y vdd BUFX4
XBUFX4_227 BUFX4_23/Y gnd BUFX4_227/Y vdd BUFX4
XFILL_0_INVX2_126 gnd vdd FILL
XBUFX4_249 INVX8_5/Y gnd BUFX4_8/A vdd BUFX4
XFILL_2_OAI21X1_1736 gnd vdd FILL
XFILL_4_DFFPOSX1_470 gnd vdd FILL
XFILL_4_DFFPOSX1_481 gnd vdd FILL
XBUFX4_238 INVX8_1/Y gnd BUFX4_238/Y vdd BUFX4
XFILL_0_INVX2_104 gnd vdd FILL
XFILL_0_INVX2_115 gnd vdd FILL
XFILL_0_INVX2_137 gnd vdd FILL
XFILL_0_INVX2_148 gnd vdd FILL
XFILL_0_INVX2_159 gnd vdd FILL
XFILL_4_DFFPOSX1_492 gnd vdd FILL
XFILL_0_INVX4_6 gnd vdd FILL
XOAI21X1_1106 OAI21X1_1106/A BUFX4_216/Y NAND2X1_471/Y gnd OAI21X1_1106/Y vdd OAI21X1
XOAI21X1_1128 OAI21X1_1128/A BUFX4_235/Y NAND2X1_493/Y gnd OAI21X1_1128/Y vdd OAI21X1
XOAI21X1_1117 INVX2_93/Y INVX4_32/Y INVX2_62/Y gnd OAI21X1_1118/C vdd OAI21X1
XFILL_1_BUFX2_382 gnd vdd FILL
XFILL_1_BUFX2_393 gnd vdd FILL
XFILL_1_OAI21X1_1304 gnd vdd FILL
XDFFPOSX1_718 BUFX2_385/A CLKBUF1_17/Y OAI21X1_985/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1337 gnd vdd FILL
XDFFPOSX1_729 BUFX2_366/A CLKBUF1_78/Y OAI21X1_1007/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_905 gnd vdd FILL
XFILL_1_DFFPOSX1_916 gnd vdd FILL
XFILL_1_OAI21X1_1326 gnd vdd FILL
XFILL_1_OAI21X1_1348 gnd vdd FILL
XDFFPOSX1_707 BUFX2_345/A CLKBUF1_54/Y OAI21X1_963/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1315 gnd vdd FILL
XOAI21X1_1139 NAND2X1_507/Y OR2X2_18/B INVX2_70/Y gnd OAI21X1_1140/C vdd OAI21X1
XFILL_0_OAI21X1_106 gnd vdd FILL
XFILL_1_DFFPOSX1_949 gnd vdd FILL
XFILL_1_DFFPOSX1_938 gnd vdd FILL
XFILL_0_OAI21X1_117 gnd vdd FILL
XFILL_1_DFFPOSX1_927 gnd vdd FILL
XFILL_1_OAI21X1_1359 gnd vdd FILL
XFILL_0_OAI21X1_128 gnd vdd FILL
XFILL_0_OAI21X1_139 gnd vdd FILL
XFILL_6_DFFPOSX1_520 gnd vdd FILL
XFILL_6_DFFPOSX1_542 gnd vdd FILL
XFILL_6_DFFPOSX1_531 gnd vdd FILL
XFILL_6_DFFPOSX1_553 gnd vdd FILL
XFILL_6_DFFPOSX1_575 gnd vdd FILL
XFILL_6_DFFPOSX1_564 gnd vdd FILL
XFILL_37_6_1 gnd vdd FILL
XFILL_0_BUFX4_16 gnd vdd FILL
XFILL_0_BUFX4_27 gnd vdd FILL
XFILL_36_1_0 gnd vdd FILL
XFILL_1_NAND2X1_305 gnd vdd FILL
XFILL_0_NAND2X1_134 gnd vdd FILL
XFILL_0_NAND2X1_123 gnd vdd FILL
XFILL_0_BUFX4_38 gnd vdd FILL
XFILL_0_BUFX4_49 gnd vdd FILL
XFILL_0_NAND2X1_112 gnd vdd FILL
XFILL_0_NAND2X1_101 gnd vdd FILL
XFILL_1_NAND2X1_327 gnd vdd FILL
XFILL_1_NAND2X1_316 gnd vdd FILL
XFILL_0_NAND2X1_156 gnd vdd FILL
XFILL_1_NAND2X1_338 gnd vdd FILL
XFILL_0_DFFPOSX1_506 gnd vdd FILL
XFILL_0_NAND2X1_145 gnd vdd FILL
XFILL_0_NAND2X1_167 gnd vdd FILL
XFILL_0_INVX1_170 gnd vdd FILL
XFILL_0_NAND2X1_189 gnd vdd FILL
XFILL_0_DFFPOSX1_539 gnd vdd FILL
XFILL_0_DFFPOSX1_528 gnd vdd FILL
XFILL_0_INVX1_181 gnd vdd FILL
XFILL_0_NAND2X1_178 gnd vdd FILL
XFILL_0_DFFPOSX1_517 gnd vdd FILL
XFILL_0_INVX1_192 gnd vdd FILL
XFILL_5_DFFPOSX1_110 gnd vdd FILL
XFILL_5_DFFPOSX1_121 gnd vdd FILL
XFILL_5_DFFPOSX1_143 gnd vdd FILL
XFILL_20_5_1 gnd vdd FILL
XFILL_5_DFFPOSX1_132 gnd vdd FILL
XFILL_5_DFFPOSX1_154 gnd vdd FILL
XFILL_5_DFFPOSX1_176 gnd vdd FILL
XFILL_5_DFFPOSX1_187 gnd vdd FILL
XFILL_5_DFFPOSX1_165 gnd vdd FILL
XFILL_5_DFFPOSX1_198 gnd vdd FILL
XOAI21X1_1651 BUFX4_123/Y INVX2_119/Y OAI21X1_1651/C gnd DFFPOSX1_38/D vdd OAI21X1
XOAI21X1_1640 INVX2_143/Y BUFX4_227/Y NAND2X1_708/Y gnd DFFPOSX1_30/D vdd OAI21X1
XOAI21X1_1662 BUFX4_11/A BUFX4_349/Y BUFX2_743/A gnd OAI21X1_1663/C vdd OAI21X1
XOAI21X1_1684 BUFX4_2/A BUFX4_362/Y BUFX2_724/A gnd OAI21X1_1685/C vdd OAI21X1
XOAI21X1_1673 BUFX4_157/Y INVX2_130/Y OAI21X1_1673/C gnd DFFPOSX1_49/D vdd OAI21X1
XOAI21X1_1695 BUFX4_149/Y INVX2_141/Y OAI21X1_1695/C gnd DFFPOSX1_60/D vdd OAI21X1
XFILL_1_OAI21X1_811 gnd vdd FILL
XFILL_0_OR2X2_19 gnd vdd FILL
XFILL_0_OAI21X1_640 gnd vdd FILL
XFILL_1_OAI21X1_800 gnd vdd FILL
XFILL_0_OAI21X1_651 gnd vdd FILL
XFILL_1_OAI21X1_855 gnd vdd FILL
XFILL_1_OAI21X1_822 gnd vdd FILL
XFILL_0_OAI21X1_662 gnd vdd FILL
XFILL_1_OAI21X1_844 gnd vdd FILL
XFILL_0_OAI21X1_673 gnd vdd FILL
XFILL_1_OAI21X1_833 gnd vdd FILL
XFILL_1_OAI21X1_888 gnd vdd FILL
XNAND3X1_38 INVX1_184/A INVX1_185/Y INVX2_94/A gnd INVX1_186/A vdd NAND3X1
XFILL_1_OAI21X1_877 gnd vdd FILL
XNAND3X1_16 INVX8_6/A OR2X2_6/Y NAND3X1_16/C gnd NAND3X1_16/Y vdd NAND3X1
XFILL_0_OAI21X1_695 gnd vdd FILL
XFILL_1_OAI21X1_866 gnd vdd FILL
XFILL_0_OAI21X1_684 gnd vdd FILL
XNAND3X1_27 bundleStartMajId_i[41] AND2X2_3/B NOR2X1_107/Y gnd XNOR2X1_45/A vdd NAND3X1
XFILL_1_AND2X2_30 gnd vdd FILL
XNAND3X1_49 NOR2X1_172/Y INVX1_196/Y INVX1_197/Y gnd OR2X2_21/B vdd NAND3X1
XFILL_1_OAI21X1_899 gnd vdd FILL
XFILL_3_DFFPOSX1_25 gnd vdd FILL
XFILL_3_DFFPOSX1_14 gnd vdd FILL
XFILL_28_6_1 gnd vdd FILL
XNOR2X1_27 OR2X2_5/A OR2X2_3/B gnd NOR2X1_27/Y vdd NOR2X1
XNOR2X1_16 NOR2X1_16/A OR2X2_3/Y gnd NOR2X1_16/Y vdd NOR2X1
XBUFX2_709 BUFX2_709/A gnd pid2_o[25] vdd BUFX2
XFILL_3_DFFPOSX1_58 gnd vdd FILL
XFILL_3_DFFPOSX1_36 gnd vdd FILL
XFILL_3_DFFPOSX1_47 gnd vdd FILL
XFILL_27_1_0 gnd vdd FILL
XNOR2X1_38 INVX4_21/Y NOR3X1_3/A gnd INVX2_44/A vdd NOR2X1
XNOR2X1_49 INVX2_46/Y INVX1_20/A gnd NOR2X1_49/Y vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XFILL_3_6_1 gnd vdd FILL
XFILL_3_DFFPOSX1_69 gnd vdd FILL
XFILL_0_NAND2X1_690 gnd vdd FILL
XFILL_0_OAI21X1_1461 gnd vdd FILL
XFILL_0_OAI21X1_1450 gnd vdd FILL
XFILL_0_OAI21X1_1472 gnd vdd FILL
XFILL_0_OAI21X1_1483 gnd vdd FILL
XFILL_0_OAI21X1_1494 gnd vdd FILL
XFILL_11_5_1 gnd vdd FILL
XFILL_4_DFFPOSX1_1 gnd vdd FILL
XFILL_0_BUFX2_3 gnd vdd FILL
XFILL_10_0_0 gnd vdd FILL
XFILL_0_BUFX2_405 gnd vdd FILL
XFILL_20_16_0 gnd vdd FILL
XFILL_0_BUFX2_416 gnd vdd FILL
XFILL_0_BUFX2_427 gnd vdd FILL
XFILL_0_BUFX2_438 gnd vdd FILL
XFILL_0_BUFX2_449 gnd vdd FILL
XFILL_19_6_1 gnd vdd FILL
XFILL_0_NAND2X1_25 gnd vdd FILL
XFILL_0_NAND2X1_14 gnd vdd FILL
XFILL_18_1_0 gnd vdd FILL
XFILL_2_OAI21X1_1566 gnd vdd FILL
XNOR2X1_106 OR2X2_5/Y INVX1_36/A gnd NOR2X1_106/Y vdd NOR2X1
XFILL_0_NAND2X1_47 gnd vdd FILL
XFILL_0_NAND2X1_36 gnd vdd FILL
XFILL_0_NAND2X1_58 gnd vdd FILL
XNOR2X1_128 INVX2_63/Y INVX1_186/A gnd INVX2_95/A vdd NOR2X1
XFILL_0_NAND2X1_69 gnd vdd FILL
XNOR2X1_117 bundleStartMajId_i[4] NOR2X1_117/B gnd NOR2X1_117/Y vdd NOR2X1
XNOR2X1_139 OR2X2_17/Y INVX1_187/A gnd XNOR2X1_61/A vdd NOR2X1
XFILL_0_INVX2_3 gnd vdd FILL
XFILL_25_15_0 gnd vdd FILL
XFILL_1_BUFX2_190 gnd vdd FILL
XFILL_1_OAI21X1_1123 gnd vdd FILL
XFILL_1_OAI21X1_1112 gnd vdd FILL
XFILL_1_OAI21X1_1101 gnd vdd FILL
XDFFPOSX1_504 BUFX2_534/A CLKBUF1_88/Y OAI21X1_559/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_713 gnd vdd FILL
XFILL_0_BUFX2_961 gnd vdd FILL
XFILL_1_OAI21X1_1156 gnd vdd FILL
XFILL_1_OAI21X1_1145 gnd vdd FILL
XDFFPOSX1_515 BUFX2_546/A CLKBUF1_47/Y OAI21X1_584/Y gnd vdd DFFPOSX1
XDFFPOSX1_537 BUFX2_570/A CLKBUF1_91/Y OAI21X1_635/Y gnd vdd DFFPOSX1
XDFFPOSX1_526 BUFX2_558/A CLKBUF1_100/Y OAI21X1_608/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_702 gnd vdd FILL
XFILL_1_DFFPOSX1_724 gnd vdd FILL
XFILL_0_BUFX2_950 gnd vdd FILL
XFILL_1_OAI21X1_1134 gnd vdd FILL
XFILL_1_OAI21X1_107 gnd vdd FILL
XFILL_1_DFFPOSX1_746 gnd vdd FILL
XFILL_0_BUFX2_972 gnd vdd FILL
XFILL_1_DFFPOSX1_757 gnd vdd FILL
XFILL_0_BUFX2_994 gnd vdd FILL
XFILL_1_OAI21X1_1178 gnd vdd FILL
XFILL_0_BUFX2_983 gnd vdd FILL
XDFFPOSX1_548 BUFX2_585/A CLKBUF1_22/Y OAI21X1_659/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_735 gnd vdd FILL
XDFFPOSX1_559 BUFX2_588/A CLKBUF1_45/Y OAI21X1_692/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1167 gnd vdd FILL
XFILL_1_OAI21X1_1189 gnd vdd FILL
XFILL_1_OAI21X1_118 gnd vdd FILL
XNAND2X1_607 BUFX4_310/Y AND2X2_30/A gnd NAND2X1_607/Y vdd NAND2X1
XNAND2X1_618 INVX1_211/A NOR3X1_17/Y gnd INVX1_212/A vdd NAND2X1
XFILL_1_DFFPOSX1_779 gnd vdd FILL
XFILL_1_OAI21X1_129 gnd vdd FILL
XFILL_1_DFFPOSX1_768 gnd vdd FILL
XINVX1_19 NOR3X1_4/C gnd INVX1_19/Y vdd INVX1
XNAND2X1_629 bundleAddress_i[43] NOR2X1_221/Y gnd INVX1_222/A vdd NAND2X1
XNAND2X1_60 BUFX2_889/A BUFX4_190/Y gnd OAI21X1_60/C vdd NAND2X1
XNAND2X1_93 BUFX2_407/A BUFX4_337/Y gnd NAND2X1_93/Y vdd NAND2X1
XNAND2X1_71 BUFX2_901/A BUFX4_196/Y gnd OAI21X1_71/C vdd NAND2X1
XNAND2X1_82 BUFX2_395/A BUFX4_388/Y gnd NAND2X1_82/Y vdd NAND2X1
XFILL_1_NAND2X1_102 gnd vdd FILL
XFILL_0_DFFPOSX1_303 gnd vdd FILL
XFILL_0_DFFPOSX1_314 gnd vdd FILL
XFILL_0_XNOR2X1_104 gnd vdd FILL
XFILL_1_NAND2X1_124 gnd vdd FILL
XFILL_1_NAND2X1_135 gnd vdd FILL
XFILL_0_16_0 gnd vdd FILL
XFILL_0_DFFPOSX1_336 gnd vdd FILL
XFILL_0_DFFPOSX1_325 gnd vdd FILL
XFILL_0_DFFPOSX1_347 gnd vdd FILL
XFILL_1_NAND2X1_168 gnd vdd FILL
XFILL_1_NAND2X1_157 gnd vdd FILL
XFILL_1_NAND2X1_179 gnd vdd FILL
XFILL_0_DFFPOSX1_358 gnd vdd FILL
XFILL_0_DFFPOSX1_369 gnd vdd FILL
XFILL_3_CLKBUF1_100 gnd vdd FILL
XFILL_3_DFFPOSX1_818 gnd vdd FILL
XFILL_3_DFFPOSX1_807 gnd vdd FILL
XFILL_0_NOR3X1_10 gnd vdd FILL
XFILL_3_DFFPOSX1_829 gnd vdd FILL
XOAI21X1_1481 XNOR2X1_99/A INVX2_99/Y INVX2_75/Y gnd NAND2X1_636/B vdd OAI21X1
XOAI21X1_1470 OAI21X1_1470/A BUFX4_294/Y OAI21X1_1470/C gnd OAI21X1_1470/Y vdd OAI21X1
XOAI21X1_1492 OAI21X1_1492/A BUFX4_294/Y OAI21X1_1492/C gnd OAI21X1_1492/Y vdd OAI21X1
XFILL_1_OAI21X1_1690 gnd vdd FILL
XFILL_1_OAI21X1_630 gnd vdd FILL
XFILL_1_NOR2X1_213 gnd vdd FILL
XFILL_1_OAI21X1_652 gnd vdd FILL
XFILL_1_OAI21X1_641 gnd vdd FILL
XFILL_0_OAI21X1_492 gnd vdd FILL
XFILL_1_NOR2X1_224 gnd vdd FILL
XFILL_3_NOR3X1_3 gnd vdd FILL
XFILL_1_OAI21X1_663 gnd vdd FILL
XFILL_2_OAI21X1_834 gnd vdd FILL
XFILL_0_OAI21X1_481 gnd vdd FILL
XFILL_0_OAI21X1_470 gnd vdd FILL
XFILL_1_OAI21X1_696 gnd vdd FILL
XFILL_1_OAI21X1_685 gnd vdd FILL
XFILL_1_OAI21X1_674 gnd vdd FILL
XFILL_5_15_0 gnd vdd FILL
XBUFX2_517 BUFX2_517/A gnd majID2_o[0] vdd BUFX2
XFILL_4_DFFPOSX1_15 gnd vdd FILL
XFILL_2_DFFPOSX1_408 gnd vdd FILL
XFILL_2_DFFPOSX1_419 gnd vdd FILL
XBUFX2_506 BUFX2_506/A gnd majID2_o[10] vdd BUFX2
XFILL_4_DFFPOSX1_37 gnd vdd FILL
XFILL_4_DFFPOSX1_26 gnd vdd FILL
XBUFX2_539 BUFX2_539/A gnd majID3_o[38] vdd BUFX2
XFILL_4_DFFPOSX1_48 gnd vdd FILL
XBUFX2_528 BUFX2_528/A gnd majID3_o[48] vdd BUFX2
XFILL_4_DFFPOSX1_59 gnd vdd FILL
XFILL_1_NAND2X1_691 gnd vdd FILL
XFILL_0_OAI21X1_1291 gnd vdd FILL
XFILL_0_DFFPOSX1_870 gnd vdd FILL
XFILL_0_OAI21X1_1280 gnd vdd FILL
XDFFPOSX1_1011 BUFX2_678/A CLKBUF1_93/Y OAI21X1_1588/Y gnd vdd DFFPOSX1
XFILL_0_DFFPOSX1_881 gnd vdd FILL
XDFFPOSX1_1000 BUFX2_389/A CLKBUF1_5/Y OAI21X1_1575/Y gnd vdd DFFPOSX1
XFILL_0_DFFPOSX1_892 gnd vdd FILL
XDFFPOSX1_1022 BUFX2_659/A CLKBUF1_73/Y OAI21X1_1599/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_202 gnd vdd FILL
XFILL_0_BUFX2_213 gnd vdd FILL
XFILL_0_BUFX2_235 gnd vdd FILL
XFILL_0_BUFX2_224 gnd vdd FILL
XFILL_0_BUFX2_246 gnd vdd FILL
XFILL_0_BUFX2_279 gnd vdd FILL
XFILL_0_BUFX2_268 gnd vdd FILL
XFILL_0_BUFX2_257 gnd vdd FILL
XFILL_14_12_1 gnd vdd FILL
XFILL_2_DFFPOSX1_942 gnd vdd FILL
XFILL_2_DFFPOSX1_920 gnd vdd FILL
XFILL_2_DFFPOSX1_931 gnd vdd FILL
XFILL_34_4_1 gnd vdd FILL
XFILL_2_DFFPOSX1_953 gnd vdd FILL
XFILL_2_DFFPOSX1_964 gnd vdd FILL
XFILL_2_DFFPOSX1_975 gnd vdd FILL
XFILL_21_2 gnd vdd FILL
XFILL_2_DFFPOSX1_997 gnd vdd FILL
XFILL_2_DFFPOSX1_986 gnd vdd FILL
XFILL_0_NAND3X1_9 gnd vdd FILL
XOAI21X1_409 OAI21X1_409/A BUFX4_199/Y OAI21X1_409/C gnd OAI21X1_409/Y vdd OAI21X1
XFILL_3_XNOR2X1_33 gnd vdd FILL
XFILL_3_XNOR2X1_22 gnd vdd FILL
XFILL_3_XNOR2X1_11 gnd vdd FILL
XDFFPOSX1_301 BUFX2_1032/A CLKBUF1_29/Y OAI21X1_219/Y gnd vdd DFFPOSX1
XDFFPOSX1_312 BUFX2_982/A CLKBUF1_5/Y OAI21X1_241/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_66 gnd vdd FILL
XFILL_3_XNOR2X1_55 gnd vdd FILL
XFILL_3_XNOR2X1_44 gnd vdd FILL
XDFFPOSX1_345 BUFX2_1018/A CLKBUF1_95/Y OAI21X1_307/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_77 gnd vdd FILL
XDFFPOSX1_323 BUFX2_994/A CLKBUF1_64/Y OAI21X1_263/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_99 gnd vdd FILL
XFILL_1_DFFPOSX1_510 gnd vdd FILL
XDFFPOSX1_356 BUFX2_393/A CLKBUF1_45/Y OAI21X1_328/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_521 gnd vdd FILL
XFILL_1_DFFPOSX1_532 gnd vdd FILL
XDFFPOSX1_334 BUFX2_1006/A CLKBUF1_83/Y OAI21X1_285/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_780 gnd vdd FILL
XFILL_0_BUFX2_791 gnd vdd FILL
XFILL_1_DFFPOSX1_543 gnd vdd FILL
XFILL_1_DFFPOSX1_565 gnd vdd FILL
XDFFPOSX1_378 BUFX2_408/A CLKBUF1_18/Y OAI21X1_350/Y gnd vdd DFFPOSX1
XDFFPOSX1_367 BUFX2_396/A CLKBUF1_6/Y OAI21X1_339/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_554 gnd vdd FILL
XDFFPOSX1_389 BUFX2_420/A CLKBUF1_44/Y OAI21X1_361/Y gnd vdd DFFPOSX1
XNAND2X1_404 BUFX2_13/A BUFX4_353/Y gnd NAND2X1_404/Y vdd NAND2X1
XNAND2X1_415 BUFX2_6/A BUFX4_340/Y gnd NAND2X1_415/Y vdd NAND2X1
XFILL_1_DFFPOSX1_598 gnd vdd FILL
XFILL_19_11_1 gnd vdd FILL
XFILL_1_DFFPOSX1_587 gnd vdd FILL
XFILL_1_DFFPOSX1_576 gnd vdd FILL
XNAND2X1_426 BUFX2_18/A BUFX4_354/Y gnd NAND2X1_426/Y vdd NAND2X1
XFILL_6_DFFPOSX1_180 gnd vdd FILL
XNAND2X1_448 BUFX2_42/A BUFX4_360/Y gnd NAND2X1_448/Y vdd NAND2X1
XNAND2X1_437 BUFX2_30/A BUFX4_384/Y gnd NAND2X1_437/Y vdd NAND2X1
XNAND2X1_459 BUFX2_54/A BUFX4_374/Y gnd NAND2X1_459/Y vdd NAND2X1
XFILL_6_DFFPOSX1_191 gnd vdd FILL
XFILL_32_13_1 gnd vdd FILL
XFILL_25_4_1 gnd vdd FILL
XFILL_0_4_1 gnd vdd FILL
XFILL_0_DFFPOSX1_111 gnd vdd FILL
XFILL_0_DFFPOSX1_100 gnd vdd FILL
XFILL_0_DFFPOSX1_122 gnd vdd FILL
XFILL_0_DFFPOSX1_133 gnd vdd FILL
XFILL_0_DFFPOSX1_144 gnd vdd FILL
XFILL_0_DFFPOSX1_155 gnd vdd FILL
XFILL_0_DFFPOSX1_166 gnd vdd FILL
XFILL_1_BUFX2_915 gnd vdd FILL
XFILL_0_DFFPOSX1_188 gnd vdd FILL
XFILL_0_DFFPOSX1_199 gnd vdd FILL
XFILL_1_BUFX2_926 gnd vdd FILL
XFILL_0_DFFPOSX1_177 gnd vdd FILL
XOAI21X1_932 BUFX4_2/A BUFX4_352/Y BUFX2_329/A gnd OAI21X1_933/C vdd OAI21X1
XOAI21X1_910 BUFX4_105/Y BUFX4_375/Y BUFX2_326/A gnd OAI21X1_911/C vdd OAI21X1
XFILL_3_DFFPOSX1_604 gnd vdd FILL
XFILL_1_BUFX2_959 gnd vdd FILL
XOAI21X1_943 BUFX4_124/Y INVX1_126/Y OAI21X1_943/C gnd OAI21X1_943/Y vdd OAI21X1
XOAI21X1_921 BUFX4_154/Y INVX1_115/Y OAI21X1_921/C gnd OAI21X1_921/Y vdd OAI21X1
XFILL_3_DFFPOSX1_615 gnd vdd FILL
XOAI21X1_976 BUFX4_162/Y BUFX4_47/Y BUFX2_369/A gnd OAI21X1_977/C vdd OAI21X1
XOAI21X1_965 BUFX4_131/Y INVX1_137/Y OAI21X1_965/C gnd OAI21X1_965/Y vdd OAI21X1
XFILL_3_DFFPOSX1_626 gnd vdd FILL
XFILL_3_DFFPOSX1_637 gnd vdd FILL
XOAI21X1_954 BUFX4_4/A BUFX4_326/Y BUFX2_341/A gnd OAI21X1_955/C vdd OAI21X1
XOAI21X1_998 BUFX4_149/Y BUFX4_65/Y BUFX2_362/A gnd OAI21X1_999/C vdd OAI21X1
XFILL_3_DFFPOSX1_648 gnd vdd FILL
XOAI21X1_987 BUFX4_303/Y INVX1_148/Y OAI21X1_987/C gnd OAI21X1_987/Y vdd OAI21X1
XFILL_3_DFFPOSX1_659 gnd vdd FILL
XFILL_37_12_1 gnd vdd FILL
XDFFPOSX1_890 BUFX2_139/A CLKBUF1_23/Y OAI21X1_1261/Y gnd vdd DFFPOSX1
XFILL_8_5_1 gnd vdd FILL
XINVX2_62 bundleAddress_i[54] gnd INVX2_62/Y vdd INVX2
XINVX2_73 bundleAddress_i[33] gnd INVX2_73/Y vdd INVX2
XINVX2_51 INVX2_51/A gnd INVX2_51/Y vdd INVX2
XFILL_2_OAI21X1_631 gnd vdd FILL
XFILL_1_OAI21X1_460 gnd vdd FILL
XFILL_7_0_0 gnd vdd FILL
XINVX2_40 NOR2X1_3/Y gnd INVX2_40/Y vdd INVX2
XFILL_1_OAI21X1_471 gnd vdd FILL
XINVX2_95 INVX2_95/A gnd INVX2_95/Y vdd INVX2
XFILL_1_OAI21X1_493 gnd vdd FILL
XFILL_1_OAI21X1_482 gnd vdd FILL
XINVX2_84 bundleAddress_i[12] gnd INVX2_84/Y vdd INVX2
XFILL_2_OAI21X1_675 gnd vdd FILL
XFILL_0_AOI21X1_3 gnd vdd FILL
XBUFX2_325 BUFX2_325/A gnd instr3_o[31] vdd BUFX2
XBUFX2_336 BUFX2_336/A gnd instr3_o[12] vdd BUFX2
XFILL_2_DFFPOSX1_205 gnd vdd FILL
XBUFX2_314 BUFX2_314/A gnd instr2_o[3] vdd BUFX2
XFILL_2_DFFPOSX1_216 gnd vdd FILL
XFILL_2_DFFPOSX1_227 gnd vdd FILL
XBUFX2_303 BUFX2_303/A gnd instr2_o[13] vdd BUFX2
XBUFX2_358 BUFX2_358/A gnd instr4_o[30] vdd BUFX2
XFILL_5_DFFPOSX1_27 gnd vdd FILL
XFILL_2_DFFPOSX1_249 gnd vdd FILL
XBUFX2_369 BUFX2_369/A gnd instr4_o[29] vdd BUFX2
XFILL_2_DFFPOSX1_238 gnd vdd FILL
XFILL_5_DFFPOSX1_16 gnd vdd FILL
XFILL_16_4_1 gnd vdd FILL
XBUFX2_347 BUFX2_347/A gnd instr3_o[2] vdd BUFX2
XFILL_5_DFFPOSX1_38 gnd vdd FILL
XFILL_5_DFFPOSX1_49 gnd vdd FILL
XFILL_1_INVX4_40 gnd vdd FILL
XOAI21X1_25 INVX2_163/Y BUFX4_198/Y OAI21X1_25/C gnd OAI21X1_25/Y vdd OAI21X1
XFILL_1_BUFX4_230 gnd vdd FILL
XOAI21X1_14 INVX2_152/Y BUFX4_219/Y OAI21X1_14/C gnd OAI21X1_14/Y vdd OAI21X1
XFILL_5_DFFPOSX1_709 gnd vdd FILL
XOAI21X1_58 INVX2_196/Y BUFX4_218/Y OAI21X1_58/C gnd OAI21X1_58/Y vdd OAI21X1
XOAI21X1_69 INVX2_5/Y BUFX4_230/Y OAI21X1_69/C gnd OAI21X1_69/Y vdd OAI21X1
XFILL_1_BUFX4_263 gnd vdd FILL
XFILL_1_BUFX4_252 gnd vdd FILL
XFILL_1_BUFX4_241 gnd vdd FILL
XOAI21X1_47 INVX2_185/Y BUFX4_188/Y OAI21X1_47/C gnd OAI21X1_47/Y vdd OAI21X1
XOAI21X1_36 INVX2_174/Y BUFX4_196/Y OAI21X1_36/C gnd OAI21X1_36/Y vdd OAI21X1
XFILL_1_BUFX4_296 gnd vdd FILL
XFILL_1_BUFX4_274 gnd vdd FILL
XFILL_1_BUFX4_285 gnd vdd FILL
XFILL_0_DFFPOSX1_12 gnd vdd FILL
XFILL_2_XNOR2X1_1 gnd vdd FILL
XFILL_0_DFFPOSX1_23 gnd vdd FILL
XFILL_0_DFFPOSX1_34 gnd vdd FILL
XFILL_0_DFFPOSX1_45 gnd vdd FILL
XFILL_0_DFFPOSX1_56 gnd vdd FILL
XFILL_0_DFFPOSX1_67 gnd vdd FILL
XFILL_0_DFFPOSX1_78 gnd vdd FILL
XFILL_0_DFFPOSX1_89 gnd vdd FILL
XFILL_2_DFFPOSX1_750 gnd vdd FILL
XBUFX2_881 BUFX2_881/A gnd tid2_o[18] vdd BUFX2
XFILL_2_DFFPOSX1_761 gnd vdd FILL
XFILL_2_DFFPOSX1_772 gnd vdd FILL
XBUFX2_870 BUFX2_870/A gnd tid2_o[28] vdd BUFX2
XFILL_2_DFFPOSX1_783 gnd vdd FILL
XBUFX2_892 BUFX2_892/A gnd tid2_o[8] vdd BUFX2
XFILL_0_NOR2X1_221 gnd vdd FILL
XFILL_0_NOR2X1_210 gnd vdd FILL
XFILL_2_DFFPOSX1_794 gnd vdd FILL
XFILL_0_NOR2X1_232 gnd vdd FILL
XOAI21X1_228 BUFX4_165/Y BUFX4_60/A BUFX2_975/A gnd OAI21X1_229/C vdd OAI21X1
XOAI21X1_206 BUFX4_175/Y BUFX4_67/Y BUFX2_992/A gnd OAI21X1_207/C vdd OAI21X1
XOAI21X1_217 INVX2_154/Y BUFX4_302/Y OAI21X1_217/C gnd OAI21X1_217/Y vdd OAI21X1
XOAI21X1_239 INVX2_165/Y BUFX4_289/Y OAI21X1_239/C gnd OAI21X1_239/Y vdd OAI21X1
XFILL_3_CLKBUF1_1 gnd vdd FILL
XAND2X2_17 NOR2X1_97/Y NOR2X1_99/Y gnd AND2X2_17/Y vdd AND2X2
XAND2X2_28 AND2X2_28/A INVX1_207/Y gnd AND2X2_29/B vdd AND2X2
XDFFPOSX1_120 BUFX2_790/A CLKBUF1_15/Y OAI21X1_1794/Y gnd vdd DFFPOSX1
XDFFPOSX1_153 BUFX2_826/A CLKBUF1_95/Y OAI21X1_1827/Y gnd vdd DFFPOSX1
XDFFPOSX1_164 NAND2X1_8/A CLKBUF1_59/Y OAI21X1_8/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_340 gnd vdd FILL
XDFFPOSX1_131 BUFX2_802/A CLKBUF1_78/Y OAI21X1_1805/Y gnd vdd DFFPOSX1
XDFFPOSX1_142 BUFX2_814/A CLKBUF1_53/Y OAI21X1_1816/Y gnd vdd DFFPOSX1
XDFFPOSX1_175 BUFX2_844/A CLKBUF1_14/Y OAI21X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_197 BUFX2_868/A CLKBUF1_98/Y OAI21X1_41/Y gnd vdd DFFPOSX1
XDFFPOSX1_186 BUFX2_856/A CLKBUF1_42/Y OAI21X1_30/Y gnd vdd DFFPOSX1
XFILL_0_NOR3X1_7 gnd vdd FILL
XNAND2X1_201 bundleStartMajId_i[33] NOR3X1_1/Y gnd NOR2X1_21/B vdd NAND2X1
XFILL_1_DFFPOSX1_384 gnd vdd FILL
XFILL_1_DFFPOSX1_373 gnd vdd FILL
XFILL_1_DFFPOSX1_362 gnd vdd FILL
XFILL_1_DFFPOSX1_351 gnd vdd FILL
XNAND2X1_234 BUFX2_500/A BUFX4_204/Y gnd OAI21X1_473/C vdd NAND2X1
XFILL_1_DFFPOSX1_395 gnd vdd FILL
XNAND2X1_223 BUFX2_495/A BUFX4_183/Y gnd OAI21X1_464/C vdd NAND2X1
XNAND2X1_212 bundleStartMajId_i[27] bundleStartMajId_i[26] gnd NOR3X1_6/B vdd NAND2X1
XFILL_4_DFFPOSX1_822 gnd vdd FILL
XNAND2X1_256 BUFX2_511/A BUFX4_231/Y gnd OAI21X1_490/C vdd NAND2X1
XFILL_4_DFFPOSX1_811 gnd vdd FILL
XNAND2X1_267 INVX1_24/A OAI21X1_663/A gnd OAI21X1_505/A vdd NAND2X1
XNAND2X1_278 bundleStartMajId_i[42] bundleStartMajId_i[41] gnd NOR2X1_69/A vdd NAND2X1
XFILL_4_DFFPOSX1_800 gnd vdd FILL
XNAND2X1_245 BUFX2_505/A BUFX4_182/Y gnd OAI21X1_480/C vdd NAND2X1
XFILL_4_DFFPOSX1_855 gnd vdd FILL
XFILL_4_DFFPOSX1_833 gnd vdd FILL
XNAND2X1_289 NOR2X1_76/Y AND2X2_13/Y gnd OR2X2_9/A vdd NAND2X1
XFILL_4_DFFPOSX1_844 gnd vdd FILL
XFILL_4_DFFPOSX1_888 gnd vdd FILL
XFILL_4_DFFPOSX1_877 gnd vdd FILL
XFILL_4_DFFPOSX1_899 gnd vdd FILL
XFILL_4_DFFPOSX1_866 gnd vdd FILL
XFILL_0_OAI21X1_6 gnd vdd FILL
XFILL_1_BUFX2_712 gnd vdd FILL
XFILL_0_BUFX2_71 gnd vdd FILL
XFILL_0_BUFX2_60 gnd vdd FILL
XFILL_0_BUFX2_82 gnd vdd FILL
XFILL_1_BUFX2_734 gnd vdd FILL
XFILL_1_BUFX2_723 gnd vdd FILL
XFILL_1_NOR2X1_52 gnd vdd FILL
XFILL_1_NOR2X1_63 gnd vdd FILL
XFILL_1_NOR2X1_41 gnd vdd FILL
XFILL_0_BUFX2_93 gnd vdd FILL
XFILL_23_18_1 gnd vdd FILL
XFILL_1_BUFX2_756 gnd vdd FILL
XFILL_0_BUFX4_319 gnd vdd FILL
XFILL_3_DFFPOSX1_412 gnd vdd FILL
XFILL_1_BUFX2_767 gnd vdd FILL
XFILL_1_NOR2X1_85 gnd vdd FILL
XFILL_0_BUFX4_308 gnd vdd FILL
XFILL_1_NOR2X1_74 gnd vdd FILL
XOAI21X1_740 BUFX4_175/Y BUFX4_71/Y BUFX2_606/A gnd OAI21X1_741/C vdd OAI21X1
XFILL_3_DFFPOSX1_401 gnd vdd FILL
XOAI21X1_751 OR2X2_15/A OR2X2_15/B INVX4_15/Y gnd OAI21X1_752/C vdd OAI21X1
XFILL_1_BUFX2_778 gnd vdd FILL
XFILL_3_DFFPOSX1_445 gnd vdd FILL
XOAI21X1_762 BUFX4_142/Y BUFX4_43/Y BUFX2_615/A gnd OAI21X1_763/C vdd OAI21X1
XOAI21X1_784 INVX4_31/Y INVX2_49/Y OAI21X1_784/C gnd OAI21X1_786/A vdd OAI21X1
XOAI21X1_773 BUFX4_122/Y BUFX4_29/Y BUFX2_621/A gnd OAI21X1_774/C vdd OAI21X1
XFILL_3_DFFPOSX1_423 gnd vdd FILL
XFILL_3_DFFPOSX1_434 gnd vdd FILL
XFILL_3_DFFPOSX1_478 gnd vdd FILL
XOAI21X1_795 BUFX4_161/Y BUFX4_63/Y BUFX2_627/A gnd OAI21X1_796/C vdd OAI21X1
XFILL_3_DFFPOSX1_456 gnd vdd FILL
XFILL_3_DFFPOSX1_489 gnd vdd FILL
XFILL_3_DFFPOSX1_467 gnd vdd FILL
XFILL_6_DFFPOSX1_949 gnd vdd FILL
XFILL_1_OAI21X1_290 gnd vdd FILL
XBUFX2_111 BUFX2_111/A gnd addr2_o[13] vdd BUFX2
XFILL_2_XNOR2X1_41 gnd vdd FILL
XBUFX2_100 BUFX2_100/A gnd addr2_o[23] vdd BUFX2
XFILL_0_NAND2X1_508 gnd vdd FILL
XFILL_2_XNOR2X1_30 gnd vdd FILL
XBUFX2_133 BUFX2_133/A gnd addr3_o[51] vdd BUFX2
XFILL_2_XNOR2X1_74 gnd vdd FILL
XFILL_2_XNOR2X1_63 gnd vdd FILL
XFILL_0_NAND2X1_519 gnd vdd FILL
XFILL_2_XNOR2X1_52 gnd vdd FILL
XBUFX2_122 BUFX2_122/A gnd addr2_o[3] vdd BUFX2
XBUFX2_144 BUFX2_144/A gnd addr3_o[41] vdd BUFX2
XBUFX2_155 BUFX2_155/A gnd addr3_o[31] vdd BUFX2
XFILL_2_XNOR2X1_85 gnd vdd FILL
XFILL_2_XNOR2X1_96 gnd vdd FILL
XBUFX2_166 INVX1_209/A gnd addr3_o[21] vdd BUFX2
XBUFX2_177 BUFX2_177/A gnd addr3_o[11] vdd BUFX2
XBUFX2_199 BUFX2_199/A gnd addr4_o[49] vdd BUFX2
XFILL_6_DFFPOSX1_39 gnd vdd FILL
XBUFX2_188 BUFX2_188/A gnd addr3_o[1] vdd BUFX2
XFILL_31_2_1 gnd vdd FILL
XFILL_28_17_1 gnd vdd FILL
XFILL_5_DFFPOSX1_506 gnd vdd FILL
XFILL_5_DFFPOSX1_517 gnd vdd FILL
XFILL_5_DFFPOSX1_539 gnd vdd FILL
XFILL_5_DFFPOSX1_528 gnd vdd FILL
XBUFX2_1003 BUFX2_1003/A gnd tid4_o[59] vdd BUFX2
XFILL_22_13_0 gnd vdd FILL
XBUFX2_1025 BUFX2_1025/A gnd tid4_o[57] vdd BUFX2
XBUFX2_1014 BUFX2_1014/A gnd tid4_o[58] vdd BUFX2
XFILL_3_DFFPOSX1_990 gnd vdd FILL
XCLKBUF1_15 BUFX4_88/Y gnd CLKBUF1_15/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_13 gnd vdd FILL
XFILL_4_DFFPOSX1_118 gnd vdd FILL
XCLKBUF1_26 BUFX4_87/Y gnd CLKBUF1_26/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_107 gnd vdd FILL
XCLKBUF1_48 BUFX4_84/Y gnd CLKBUF1_48/Y vdd CLKBUF1
XCLKBUF1_37 BUFX4_89/Y gnd CLKBUF1_37/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_57 gnd vdd FILL
XFILL_1_DFFPOSX1_46 gnd vdd FILL
XCLKBUF1_59 BUFX4_91/Y gnd CLKBUF1_59/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_24 gnd vdd FILL
XFILL_4_DFFPOSX1_129 gnd vdd FILL
XFILL_1_DFFPOSX1_35 gnd vdd FILL
XFILL_1_DFFPOSX1_68 gnd vdd FILL
XFILL_1_DFFPOSX1_79 gnd vdd FILL
XBUFX4_80 BUFX4_80/A gnd BUFX4_80/Y vdd BUFX4
XBUFX4_91 clock_i gnd BUFX4_91/Y vdd BUFX4
XFILL_3_18_1 gnd vdd FILL
XFILL_2_BUFX4_228 gnd vdd FILL
XFILL_0_OAI21X1_1824 gnd vdd FILL
XFILL_0_OAI21X1_1813 gnd vdd FILL
XFILL_0_OAI21X1_1802 gnd vdd FILL
XFILL_2_DFFPOSX1_591 gnd vdd FILL
XFILL_2_DFFPOSX1_580 gnd vdd FILL
XFILL_22_2_1 gnd vdd FILL
XFILL_27_12_0 gnd vdd FILL
XFILL_1_DFFPOSX1_181 gnd vdd FILL
XFILL_1_DFFPOSX1_170 gnd vdd FILL
XXNOR2X1_1 NOR2X1_5/Y bundleStartMajId_i[54] gnd XNOR2X1_1/Y vdd XNOR2X1
XFILL_1_DFFPOSX1_192 gnd vdd FILL
XFILL_8_17_1 gnd vdd FILL
XFILL_4_DFFPOSX1_630 gnd vdd FILL
XFILL_5_3_1 gnd vdd FILL
XFILL_4_DFFPOSX1_652 gnd vdd FILL
XFILL_4_DFFPOSX1_663 gnd vdd FILL
XFILL_4_DFFPOSX1_641 gnd vdd FILL
XFILL_4_DFFPOSX1_696 gnd vdd FILL
XFILL_4_DFFPOSX1_674 gnd vdd FILL
XFILL_2_13_0 gnd vdd FILL
XFILL_4_DFFPOSX1_685 gnd vdd FILL
XFILL_13_2_1 gnd vdd FILL
XFILL_1_BUFX2_520 gnd vdd FILL
XFILL_0_BUFX4_105 gnd vdd FILL
XINVX1_1 bundleStartMajId_i[50] gnd INVX1_1/Y vdd INVX1
XFILL_1_BUFX2_531 gnd vdd FILL
XFILL_1_BUFX2_564 gnd vdd FILL
XFILL_3_DFFPOSX1_220 gnd vdd FILL
XFILL_1_BUFX2_575 gnd vdd FILL
XFILL_0_BUFX4_149 gnd vdd FILL
XFILL_0_BUFX4_138 gnd vdd FILL
XFILL_0_BUFX4_127 gnd vdd FILL
XFILL_0_BUFX4_116 gnd vdd FILL
XFILL_3_DFFPOSX1_242 gnd vdd FILL
XFILL_1_OAI21X1_1519 gnd vdd FILL
XFILL_3_DFFPOSX1_253 gnd vdd FILL
XFILL_3_DFFPOSX1_264 gnd vdd FILL
XOAI21X1_570 OR2X2_4/A NOR2X1_70/B OAI21X1_570/C gnd OAI21X1_571/A vdd OAI21X1
XOAI21X1_581 OAI21X1_581/A AOI21X1_7/Y OAI21X1_581/C gnd OAI21X1_581/Y vdd OAI21X1
XFILL_3_DFFPOSX1_231 gnd vdd FILL
XFILL_1_OAI21X1_1508 gnd vdd FILL
XOAI21X1_592 OR2X2_9/B OR2X2_9/A OAI21X1_592/C gnd OAI21X1_594/A vdd OAI21X1
XFILL_1_BUFX2_16 gnd vdd FILL
XFILL_3_DFFPOSX1_275 gnd vdd FILL
XFILL_1_BUFX2_49 gnd vdd FILL
XFILL_3_DFFPOSX1_297 gnd vdd FILL
XFILL_3_DFFPOSX1_286 gnd vdd FILL
XFILL_6_DFFPOSX1_702 gnd vdd FILL
XFILL_6_DFFPOSX1_713 gnd vdd FILL
XFILL_6_DFFPOSX1_735 gnd vdd FILL
XFILL_6_DFFPOSX1_724 gnd vdd FILL
XFILL_5_DFFPOSX1_5 gnd vdd FILL
XFILL_6_DFFPOSX1_746 gnd vdd FILL
XFILL_6_DFFPOSX1_757 gnd vdd FILL
XFILL_7_12_0 gnd vdd FILL
XFILL_0_NAND2X1_305 gnd vdd FILL
XFILL_0_NAND2X1_316 gnd vdd FILL
XFILL_0_OAI21X1_1109 gnd vdd FILL
XFILL_0_NAND2X1_349 gnd vdd FILL
XFILL_0_NAND2X1_327 gnd vdd FILL
XFILL_11_10_1 gnd vdd FILL
XFILL_0_NAND2X1_338 gnd vdd FILL
XFILL_39_3 gnd vdd FILL
XFILL_1_NOR2X1_7 gnd vdd FILL
XFILL_1_DFFPOSX1_1011 gnd vdd FILL
XFILL_1_DFFPOSX1_1000 gnd vdd FILL
XFILL_1_DFFPOSX1_1022 gnd vdd FILL
XFILL_5_DFFPOSX1_336 gnd vdd FILL
XFILL_5_DFFPOSX1_325 gnd vdd FILL
XFILL_5_DFFPOSX1_303 gnd vdd FILL
XFILL_5_DFFPOSX1_314 gnd vdd FILL
XFILL_5_DFFPOSX1_358 gnd vdd FILL
XFILL_5_DFFPOSX1_347 gnd vdd FILL
XFILL_5_DFFPOSX1_369 gnd vdd FILL
XOAI21X1_1800 BUFX4_363/Y INVX2_172/Y NAND2X1_741/Y gnd OAI21X1_1800/Y vdd OAI21X1
XOAI21X1_1811 BUFX4_352/Y INVX2_183/Y NAND2X1_752/Y gnd OAI21X1_1811/Y vdd OAI21X1
XOAI21X1_1822 BUFX4_377/Y INVX2_194/Y NAND2X1_763/Y gnd OAI21X1_1822/Y vdd OAI21X1
XFILL_1_NAND2X1_18 gnd vdd FILL
XINVX4_19 bundleStartMajId_i[23] gnd INVX4_19/Y vdd INVX4
XFILL_0_OAI21X1_822 gnd vdd FILL
XFILL_0_OAI21X1_811 gnd vdd FILL
XFILL_0_OAI21X1_800 gnd vdd FILL
XFILL_0_OAI21X1_855 gnd vdd FILL
XFILL_0_OAI21X1_866 gnd vdd FILL
XFILL_0_OAI21X1_844 gnd vdd FILL
XFILL_0_OAI21X1_833 gnd vdd FILL
XFILL_0_OAI21X1_888 gnd vdd FILL
XFILL_0_OAI21X1_877 gnd vdd FILL
XFILL_0_OAI21X1_899 gnd vdd FILL
XFILL_2_DFFPOSX1_36 gnd vdd FILL
XFILL_2_DFFPOSX1_25 gnd vdd FILL
XFILL_2_DFFPOSX1_14 gnd vdd FILL
XFILL_2_DFFPOSX1_69 gnd vdd FILL
XFILL_2_DFFPOSX1_58 gnd vdd FILL
XFILL_2_DFFPOSX1_47 gnd vdd FILL
XFILL_13_18_0 gnd vdd FILL
XFILL_0_OAI21X1_1621 gnd vdd FILL
XFILL_0_OAI21X1_1632 gnd vdd FILL
XFILL_0_OAI21X1_1643 gnd vdd FILL
XFILL_0_OAI21X1_1610 gnd vdd FILL
XFILL_0_OAI21X1_1676 gnd vdd FILL
XFILL_0_OAI21X1_1665 gnd vdd FILL
XFILL_0_OAI21X1_1654 gnd vdd FILL
XFILL_0_OAI21X1_1698 gnd vdd FILL
XFILL_0_OAI21X1_1687 gnd vdd FILL
XFILL_0_BUFX4_7 gnd vdd FILL
XFILL_5_DFFPOSX1_881 gnd vdd FILL
XFILL_5_DFFPOSX1_870 gnd vdd FILL
XFILL_0_BUFX2_609 gnd vdd FILL
XFILL_5_DFFPOSX1_892 gnd vdd FILL
XFILL_4_DFFPOSX1_1004 gnd vdd FILL
XFILL_4_DFFPOSX1_1015 gnd vdd FILL
XFILL_1_XNOR2X1_82 gnd vdd FILL
XFILL_1_XNOR2X1_71 gnd vdd FILL
XFILL_1_XNOR2X1_60 gnd vdd FILL
XFILL_4_DFFPOSX1_1026 gnd vdd FILL
XFILL_1_XNOR2X1_93 gnd vdd FILL
XFILL_18_17_0 gnd vdd FILL
XFILL_34_10_1 gnd vdd FILL
XBUFX4_206 BUFX4_21/Y gnd BUFX4_206/Y vdd BUFX4
XBUFX4_228 BUFX4_26/Y gnd BUFX4_228/Y vdd BUFX4
XBUFX4_217 BUFX4_20/Y gnd BUFX4_217/Y vdd BUFX4
XFILL_0_INVX2_105 gnd vdd FILL
XFILL_4_DFFPOSX1_471 gnd vdd FILL
XFILL_4_DFFPOSX1_482 gnd vdd FILL
XFILL_4_DFFPOSX1_460 gnd vdd FILL
XBUFX4_239 INVX8_1/Y gnd BUFX4_239/Y vdd BUFX4
XFILL_0_INVX2_116 gnd vdd FILL
XFILL_0_INVX2_127 gnd vdd FILL
XFILL_0_INVX2_138 gnd vdd FILL
XFILL_4_DFFPOSX1_493 gnd vdd FILL
XFILL_0_INVX2_149 gnd vdd FILL
XFILL_0_INVX4_7 gnd vdd FILL
XFILL_1_BUFX2_372 gnd vdd FILL
XFILL_1_BUFX2_361 gnd vdd FILL
XOAI21X1_1107 INVX1_184/Y INVX1_185/A BUFX4_241/Y gnd OAI21X1_1108/A vdd OAI21X1
XOAI21X1_1118 NAND2X1_476/Y INVX2_94/Y OAI21X1_1118/C gnd OAI21X1_1119/A vdd OAI21X1
XOAI21X1_1129 XNOR2X1_57/Y BUFX4_224/Y NAND2X1_496/Y gnd OAI21X1_1129/Y vdd OAI21X1
XFILL_1_BUFX2_383 gnd vdd FILL
XFILL_1_OAI21X1_1305 gnd vdd FILL
XAND2X2_1 NOR2X1_3/Y NOR2X1_4/Y gnd AND2X2_1/Y vdd AND2X2
XFILL_1_OAI21X1_1338 gnd vdd FILL
XFILL_1_DFFPOSX1_906 gnd vdd FILL
XFILL_1_OAI21X1_1327 gnd vdd FILL
XDFFPOSX1_719 BUFX2_386/A CLKBUF1_71/Y OAI21X1_987/Y gnd vdd DFFPOSX1
XDFFPOSX1_708 BUFX2_346/A CLKBUF1_6/Y OAI21X1_965/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1316 gnd vdd FILL
XFILL_0_OAI21X1_107 gnd vdd FILL
XFILL_0_OAI21X1_118 gnd vdd FILL
XFILL_1_DFFPOSX1_939 gnd vdd FILL
XFILL_1_DFFPOSX1_917 gnd vdd FILL
XFILL_1_OAI21X1_1349 gnd vdd FILL
XFILL_1_DFFPOSX1_928 gnd vdd FILL
XFILL_6_DFFPOSX1_510 gnd vdd FILL
XFILL_0_OAI21X1_129 gnd vdd FILL
XFILL_36_18_0 gnd vdd FILL
XFILL_2_1 gnd vdd FILL
XFILL_6_DFFPOSX1_598 gnd vdd FILL
XFILL_0_BUFX4_17 gnd vdd FILL
XFILL_36_1_1 gnd vdd FILL
XFILL_0_NAND2X1_113 gnd vdd FILL
XFILL_0_NAND2X1_124 gnd vdd FILL
XFILL_0_BUFX4_39 gnd vdd FILL
XFILL_0_NAND2X1_102 gnd vdd FILL
XFILL_0_BUFX4_28 gnd vdd FILL
XFILL_1_NAND2X1_306 gnd vdd FILL
XFILL_1_NAND2X1_328 gnd vdd FILL
XFILL_1_NAND2X1_317 gnd vdd FILL
XFILL_0_NAND2X1_168 gnd vdd FILL
XFILL_0_NAND2X1_135 gnd vdd FILL
XFILL_1_NAND2X1_339 gnd vdd FILL
XFILL_0_NAND2X1_157 gnd vdd FILL
XFILL_0_NAND2X1_146 gnd vdd FILL
XFILL_0_INVX1_171 gnd vdd FILL
XFILL_1_AOI21X1_60 gnd vdd FILL
XFILL_0_INVX1_182 gnd vdd FILL
XFILL_0_DFFPOSX1_529 gnd vdd FILL
XFILL_0_DFFPOSX1_507 gnd vdd FILL
XFILL_0_INVX1_160 gnd vdd FILL
XFILL_0_NAND2X1_179 gnd vdd FILL
XFILL_0_DFFPOSX1_518 gnd vdd FILL
XFILL_5_DFFPOSX1_111 gnd vdd FILL
XFILL_5_DFFPOSX1_100 gnd vdd FILL
XFILL_2_CLKBUF1_100 gnd vdd FILL
XFILL_0_INVX1_193 gnd vdd FILL
XFILL_5_DFFPOSX1_133 gnd vdd FILL
XFILL_5_DFFPOSX1_144 gnd vdd FILL
XFILL_5_DFFPOSX1_122 gnd vdd FILL
XFILL_5_DFFPOSX1_155 gnd vdd FILL
XFILL_5_DFFPOSX1_166 gnd vdd FILL
XFILL_5_DFFPOSX1_177 gnd vdd FILL
XFILL_5_DFFPOSX1_188 gnd vdd FILL
XFILL_5_DFFPOSX1_199 gnd vdd FILL
XOAI21X1_1630 INVX2_133/Y BUFX4_198/Y NAND2X1_698/Y gnd DFFPOSX1_20/D vdd OAI21X1
XOAI21X1_1641 INVX2_144/Y BUFX4_190/Y NAND2X1_709/Y gnd DFFPOSX1_31/D vdd OAI21X1
XOAI21X1_1674 BUFX4_11/Y BUFX4_341/Y BUFX2_719/A gnd OAI21X1_1675/C vdd OAI21X1
XOAI21X1_1663 BUFX4_140/Y INVX2_125/Y OAI21X1_1663/C gnd DFFPOSX1_44/D vdd OAI21X1
XOAI21X1_1652 BUFX4_4/A BUFX4_377/Y BUFX2_736/A gnd OAI21X1_1653/C vdd OAI21X1
XFILL_0_OAI21X1_641 gnd vdd FILL
XFILL_1_OAI21X1_812 gnd vdd FILL
XOAI21X1_1696 BUFX4_108/Y BUFX4_334/Y BUFX2_731/A gnd OAI21X1_1697/C vdd OAI21X1
XFILL_0_OAI21X1_630 gnd vdd FILL
XOAI21X1_1685 BUFX4_176/Y INVX2_136/Y OAI21X1_1685/C gnd DFFPOSX1_55/D vdd OAI21X1
XFILL_1_OAI21X1_801 gnd vdd FILL
XFILL_0_OAI21X1_652 gnd vdd FILL
XFILL_1_OAI21X1_823 gnd vdd FILL
XFILL_1_OAI21X1_845 gnd vdd FILL
XFILL_0_OAI21X1_663 gnd vdd FILL
XFILL_1_OAI21X1_834 gnd vdd FILL
XFILL_0_OAI21X1_674 gnd vdd FILL
XFILL_1_OAI21X1_867 gnd vdd FILL
XNAND3X1_39 bundleAddress_i[50] bundleAddress_i[49] INVX2_96/Y gnd NOR2X1_185/A vdd
+ NAND3X1
XFILL_1_OAI21X1_878 gnd vdd FILL
XNAND3X1_17 bundleStartMajId_i[32] AND2X2_6/Y NOR2X1_72/Y gnd OR2X2_7/A vdd NAND3X1
XNAND3X1_28 NOR2X1_28/Y INVX1_13/A NOR2X1_109/Y gnd NOR3X1_7/C vdd NAND3X1
XFILL_0_OAI21X1_696 gnd vdd FILL
XFILL_1_OAI21X1_856 gnd vdd FILL
XFILL_0_OAI21X1_685 gnd vdd FILL
XFILL_1_OAI21X1_889 gnd vdd FILL
XFILL_1_AND2X2_31 gnd vdd FILL
XFILL_1_AND2X2_20 gnd vdd FILL
XFILL_3_DFFPOSX1_26 gnd vdd FILL
XFILL_3_DFFPOSX1_15 gnd vdd FILL
XNOR2X1_28 OR2X2_4/A OR2X2_4/B gnd NOR2X1_28/Y vdd NOR2X1
XNOR2X1_17 INVX4_10/Y NOR3X1_1/C gnd NOR2X1_17/Y vdd NOR2X1
XFILL_3_DFFPOSX1_59 gnd vdd FILL
XFILL_3_DFFPOSX1_37 gnd vdd FILL
XFILL_27_1_1 gnd vdd FILL
XFILL_3_DFFPOSX1_48 gnd vdd FILL
XNOR2X1_39 INVX2_30/Y INVX2_31/Y gnd INVX1_33/A vdd NOR2X1
XFILL_2_1_1 gnd vdd FILL
XFILL_0_OAI21X1_1440 gnd vdd FILL
XFILL_0_OAI21X1_1451 gnd vdd FILL
XFILL_0_NAND2X1_680 gnd vdd FILL
XFILL_0_NAND2X1_691 gnd vdd FILL
XFILL_0_OAI21X1_1473 gnd vdd FILL
XFILL_0_OAI21X1_1462 gnd vdd FILL
XFILL_0_OAI21X1_1484 gnd vdd FILL
XFILL_0_OAI21X1_1495 gnd vdd FILL
XFILL_4_DFFPOSX1_2 gnd vdd FILL
XFILL_0_BUFX2_4 gnd vdd FILL
XFILL_10_0_1 gnd vdd FILL
XFILL_0_BUFX2_439 gnd vdd FILL
XFILL_0_BUFX2_428 gnd vdd FILL
XFILL_0_BUFX2_406 gnd vdd FILL
XFILL_0_BUFX2_417 gnd vdd FILL
XFILL_20_16_1 gnd vdd FILL
XFILL_2_OAI21X1_1512 gnd vdd FILL
XFILL_0_NAND2X1_15 gnd vdd FILL
XFILL_0_NAND2X1_26 gnd vdd FILL
XFILL_18_1_1 gnd vdd FILL
XFILL_4_DFFPOSX1_290 gnd vdd FILL
XFILL_0_NAND2X1_37 gnd vdd FILL
XFILL_2_OAI21X1_1545 gnd vdd FILL
XNOR2X1_129 INVX2_96/A INVX2_95/Y gnd NOR2X1_129/Y vdd NOR2X1
XNOR2X1_118 INVX2_38/Y NOR3X1_11/C gnd NOR2X1_119/B vdd NOR2X1
XFILL_0_NAND2X1_59 gnd vdd FILL
XFILL_0_NAND2X1_48 gnd vdd FILL
XNOR2X1_107 OR2X2_3/Y NOR3X1_9/A gnd NOR2X1_107/Y vdd NOR2X1
XFILL_0_INVX2_4 gnd vdd FILL
XFILL_30_8_0 gnd vdd FILL
XFILL_25_15_1 gnd vdd FILL
XFILL_1_BUFX2_180 gnd vdd FILL
XFILL_1_OAI21X1_1102 gnd vdd FILL
XFILL_1_OAI21X1_1113 gnd vdd FILL
XDFFPOSX1_505 MUX2X1_1/B CLKBUF1_18/Y NOR2X1_66/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_951 gnd vdd FILL
XFILL_1_OAI21X1_1124 gnd vdd FILL
XFILL_1_OAI21X1_1146 gnd vdd FILL
XFILL_1_DFFPOSX1_714 gnd vdd FILL
XDFFPOSX1_516 NOR2X1_73/A CLKBUF1_88/Y AOI21X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_527 BUFX2_559/A CLKBUF1_84/Y OAI21X1_611/Y gnd vdd DFFPOSX1
XDFFPOSX1_538 BUFX2_571/A CLKBUF1_79/Y OAI21X1_637/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_940 gnd vdd FILL
XFILL_1_DFFPOSX1_703 gnd vdd FILL
XFILL_1_OAI21X1_1135 gnd vdd FILL
XFILL_0_BUFX2_973 gnd vdd FILL
XFILL_1_DFFPOSX1_747 gnd vdd FILL
XFILL_1_DFFPOSX1_725 gnd vdd FILL
XFILL_1_DFFPOSX1_758 gnd vdd FILL
XFILL_1_DFFPOSX1_736 gnd vdd FILL
XFILL_1_OAI21X1_108 gnd vdd FILL
XFILL_0_BUFX2_984 gnd vdd FILL
XFILL_1_OAI21X1_1168 gnd vdd FILL
XFILL_1_OAI21X1_1179 gnd vdd FILL
XFILL_1_OAI21X1_1157 gnd vdd FILL
XFILL_0_BUFX2_995 gnd vdd FILL
XFILL_0_BUFX2_962 gnd vdd FILL
XDFFPOSX1_549 BUFX2_586/A CLKBUF1_48/Y OAI21X1_661/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_119 gnd vdd FILL
XFILL_1_DFFPOSX1_769 gnd vdd FILL
XNAND2X1_608 INVX1_208/Y INVX2_106/A gnd XNOR2X1_83/A vdd NAND2X1
XNAND2X1_619 bundleAddress_i[14] bundleAddress_i[13] gnd NOR2X1_207/B vdd NAND2X1
XFILL_6_DFFPOSX1_362 gnd vdd FILL
XFILL_6_DFFPOSX1_351 gnd vdd FILL
XFILL_6_DFFPOSX1_395 gnd vdd FILL
XFILL_6_DFFPOSX1_384 gnd vdd FILL
XFILL_6_DFFPOSX1_373 gnd vdd FILL
XFILL_38_9_0 gnd vdd FILL
XNAND2X1_61 BUFX2_890/A BUFX4_220/Y gnd OAI21X1_61/C vdd NAND2X1
XNAND2X1_50 BUFX2_878/A BUFX4_228/Y gnd OAI21X1_50/C vdd NAND2X1
XNAND2X1_72 BUFX2_393/A BUFX4_321/Y gnd NAND2X1_72/Y vdd NAND2X1
XNAND2X1_83 BUFX2_396/A BUFX4_387/Y gnd NAND2X1_83/Y vdd NAND2X1
XNAND2X1_94 BUFX2_408/A BUFX4_383/Y gnd NAND2X1_94/Y vdd NAND2X1
XFILL_0_XNOR2X1_90 gnd vdd FILL
XFILL_1_NAND2X1_114 gnd vdd FILL
XFILL_0_DFFPOSX1_304 gnd vdd FILL
XFILL_0_DFFPOSX1_315 gnd vdd FILL
XFILL_0_16_1 gnd vdd FILL
XFILL_1_NAND2X1_147 gnd vdd FILL
XFILL_0_DFFPOSX1_337 gnd vdd FILL
XFILL_0_DFFPOSX1_348 gnd vdd FILL
XFILL_0_DFFPOSX1_326 gnd vdd FILL
XFILL_1_NAND2X1_169 gnd vdd FILL
XFILL_21_8_0 gnd vdd FILL
XFILL_0_DFFPOSX1_359 gnd vdd FILL
XFILL_3_CLKBUF1_101 gnd vdd FILL
XFILL_3_DFFPOSX1_808 gnd vdd FILL
XFILL_3_DFFPOSX1_819 gnd vdd FILL
XFILL_24_10_0 gnd vdd FILL
XFILL_0_NOR3X1_11 gnd vdd FILL
XOAI21X1_1460 NAND2X1_633/Y BUFX4_292/Y OAI21X1_1460/C gnd OAI21X1_1460/Y vdd OAI21X1
XOAI21X1_1471 INVX2_109/Y NOR2X1_145/A INVX2_73/Y gnd NAND2X1_634/B vdd OAI21X1
XOAI21X1_1482 NAND2X1_636/Y BUFX4_297/Y OAI21X1_1482/C gnd OAI21X1_1482/Y vdd OAI21X1
XOAI21X1_1493 INVX1_223/A NAND2X1_637/Y INVX4_41/Y gnd OAI21X1_1494/C vdd OAI21X1
XFILL_1_OAI21X1_1691 gnd vdd FILL
XFILL_1_OAI21X1_1680 gnd vdd FILL
XFILL_1_NOR2X1_203 gnd vdd FILL
XFILL_1_NOR2X1_214 gnd vdd FILL
XFILL_1_OAI21X1_620 gnd vdd FILL
XFILL_1_OAI21X1_653 gnd vdd FILL
XFILL_1_OAI21X1_642 gnd vdd FILL
XFILL_1_OAI21X1_631 gnd vdd FILL
XFILL_3_NOR3X1_4 gnd vdd FILL
XFILL_0_OAI21X1_460 gnd vdd FILL
XFILL_0_OAI21X1_482 gnd vdd FILL
XFILL_0_OAI21X1_471 gnd vdd FILL
XFILL_2_OAI21X1_868 gnd vdd FILL
XFILL_0_OAI21X1_493 gnd vdd FILL
XFILL_1_OAI21X1_664 gnd vdd FILL
XFILL_1_OAI21X1_697 gnd vdd FILL
XFILL_1_INVX1_103 gnd vdd FILL
XFILL_1_INVX1_114 gnd vdd FILL
XFILL_1_OAI21X1_686 gnd vdd FILL
XFILL_1_OAI21X1_675 gnd vdd FILL
XFILL_29_9_0 gnd vdd FILL
XFILL_5_15_1 gnd vdd FILL
XFILL_2_DFFPOSX1_409 gnd vdd FILL
XBUFX2_518 BUFX2_518/A gnd majID2_o[56] vdd BUFX2
XFILL_4_9_0 gnd vdd FILL
XBUFX2_507 BUFX2_507/A gnd majID2_o[9] vdd BUFX2
XFILL_4_DFFPOSX1_27 gnd vdd FILL
XFILL_4_DFFPOSX1_38 gnd vdd FILL
XFILL_4_DFFPOSX1_16 gnd vdd FILL
XBUFX2_529 BUFX2_529/A gnd majID3_o[47] vdd BUFX2
XFILL_4_DFFPOSX1_49 gnd vdd FILL
XFILL_2_OR2X2_1 gnd vdd FILL
XFILL_1_NAND2X1_692 gnd vdd FILL
XFILL_1_NAND2X1_670 gnd vdd FILL
XFILL_0_OAI21X1_1292 gnd vdd FILL
XFILL_0_OAI21X1_1281 gnd vdd FILL
XFILL_0_OAI21X1_1270 gnd vdd FILL
XFILL_0_DFFPOSX1_860 gnd vdd FILL
XFILL_0_DFFPOSX1_882 gnd vdd FILL
XDFFPOSX1_1001 BUFX2_390/A CLKBUF1_5/Y OAI21X1_1576/Y gnd vdd DFFPOSX1
XFILL_0_DFFPOSX1_871 gnd vdd FILL
XFILL_0_DFFPOSX1_893 gnd vdd FILL
XFILL_12_8_0 gnd vdd FILL
XDFFPOSX1_1012 BUFX2_679/A CLKBUF1_8/Y OAI21X1_1589/Y gnd vdd DFFPOSX1
XDFFPOSX1_1023 BUFX2_660/A CLKBUF1_45/Y OAI21X1_1600/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_203 gnd vdd FILL
XFILL_0_BUFX2_214 gnd vdd FILL
XFILL_0_BUFX2_236 gnd vdd FILL
XFILL_0_BUFX2_247 gnd vdd FILL
XFILL_0_BUFX2_225 gnd vdd FILL
XFILL_0_BUFX2_269 gnd vdd FILL
XFILL_0_BUFX2_258 gnd vdd FILL
XFILL_4_10_0 gnd vdd FILL
XFILL_2_DFFPOSX1_932 gnd vdd FILL
XFILL_2_DFFPOSX1_921 gnd vdd FILL
XFILL_2_OAI21X1_1353 gnd vdd FILL
XFILL_2_DFFPOSX1_910 gnd vdd FILL
XFILL_2_DFFPOSX1_954 gnd vdd FILL
XFILL_2_DFFPOSX1_943 gnd vdd FILL
XFILL_2_OAI21X1_1386 gnd vdd FILL
XFILL_2_DFFPOSX1_965 gnd vdd FILL
XFILL_2_DFFPOSX1_976 gnd vdd FILL
XFILL_2_DFFPOSX1_998 gnd vdd FILL
XFILL_2_DFFPOSX1_987 gnd vdd FILL
XFILL_21_3 gnd vdd FILL
XFILL_3_XNOR2X1_23 gnd vdd FILL
XFILL_3_XNOR2X1_56 gnd vdd FILL
XDFFPOSX1_313 BUFX2_983/A CLKBUF1_22/Y OAI21X1_243/Y gnd vdd DFFPOSX1
XDFFPOSX1_302 BUFX2_971/A CLKBUF1_83/Y OAI21X1_221/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_34 gnd vdd FILL
XDFFPOSX1_346 BUFX2_1019/A CLKBUF1_98/Y OAI21X1_309/Y gnd vdd DFFPOSX1
XDFFPOSX1_335 BUFX2_1007/A CLKBUF1_27/Y OAI21X1_287/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_89 gnd vdd FILL
XFILL_3_XNOR2X1_78 gnd vdd FILL
XFILL_1_DFFPOSX1_533 gnd vdd FILL
XDFFPOSX1_324 BUFX2_995/A CLKBUF1_56/Y OAI21X1_265/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_67 gnd vdd FILL
XFILL_1_DFFPOSX1_500 gnd vdd FILL
XFILL_1_DFFPOSX1_522 gnd vdd FILL
XFILL_1_DFFPOSX1_511 gnd vdd FILL
XFILL_0_BUFX2_781 gnd vdd FILL
XFILL_1_DFFPOSX1_544 gnd vdd FILL
XFILL_0_BUFX2_792 gnd vdd FILL
XFILL_1_DFFPOSX1_555 gnd vdd FILL
XFILL_1_DFFPOSX1_566 gnd vdd FILL
XDFFPOSX1_357 BUFX2_394/A CLKBUF1_45/Y OAI21X1_329/Y gnd vdd DFFPOSX1
XDFFPOSX1_368 BUFX2_397/A CLKBUF1_94/Y OAI21X1_340/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_770 gnd vdd FILL
XDFFPOSX1_379 BUFX2_409/A CLKBUF1_18/Y OAI21X1_351/Y gnd vdd DFFPOSX1
XNAND2X1_405 BUFX2_24/A BUFX4_312/Y gnd NAND2X1_405/Y vdd NAND2X1
XNAND2X1_416 BUFX2_7/A BUFX4_340/Y gnd NAND2X1_416/Y vdd NAND2X1
XFILL_1_DFFPOSX1_599 gnd vdd FILL
XFILL_1_DFFPOSX1_588 gnd vdd FILL
XNAND2X1_427 BUFX2_19/A OAI21X1_5/A gnd NAND2X1_427/Y vdd NAND2X1
XFILL_1_DFFPOSX1_577 gnd vdd FILL
XNAND2X1_449 BUFX2_43/A BUFX4_339/Y gnd NAND2X1_449/Y vdd NAND2X1
XNAND2X1_438 BUFX2_31/A BUFX4_350/Y gnd NAND2X1_438/Y vdd NAND2X1
XFILL_10_16_0 gnd vdd FILL
XFILL_0_DFFPOSX1_112 gnd vdd FILL
XFILL_0_DFFPOSX1_123 gnd vdd FILL
XFILL_0_DFFPOSX1_101 gnd vdd FILL
XFILL_0_DFFPOSX1_134 gnd vdd FILL
XFILL_0_DFFPOSX1_156 gnd vdd FILL
XFILL_0_DFFPOSX1_145 gnd vdd FILL
XOAI21X1_900 INVX1_101/Y BUFX4_197/Y OAI21X1_900/C gnd OAI21X1_900/Y vdd OAI21X1
XFILL_0_DFFPOSX1_178 gnd vdd FILL
XFILL_0_DFFPOSX1_189 gnd vdd FILL
XFILL_1_BUFX2_916 gnd vdd FILL
XFILL_1_BUFX2_905 gnd vdd FILL
XFILL_1_BUFX2_938 gnd vdd FILL
XFILL_0_DFFPOSX1_167 gnd vdd FILL
XOAI21X1_933 BUFX4_136/Y INVX1_121/Y OAI21X1_933/C gnd OAI21X1_933/Y vdd OAI21X1
XOAI21X1_911 BUFX4_140/Y INVX1_110/Y OAI21X1_911/C gnd OAI21X1_911/Y vdd OAI21X1
XFILL_4_CLKBUF1_102 gnd vdd FILL
XOAI21X1_922 BUFX4_1/Y BUFX4_330/Y BUFX2_354/A gnd OAI21X1_923/C vdd OAI21X1
XFILL_1_BUFX2_949 gnd vdd FILL
XOAI21X1_944 BUFX4_100/Y BUFX4_352/Y BUFX2_335/A gnd OAI21X1_945/C vdd OAI21X1
XFILL_3_DFFPOSX1_627 gnd vdd FILL
XFILL_3_DFFPOSX1_605 gnd vdd FILL
XFILL_3_DFFPOSX1_616 gnd vdd FILL
XFILL_3_DFFPOSX1_638 gnd vdd FILL
XOAI21X1_955 BUFX4_124/Y INVX1_132/Y OAI21X1_955/C gnd OAI21X1_955/Y vdd OAI21X1
XOAI21X1_966 BUFX4_7/A BUFX4_315/Y BUFX2_347/A gnd OAI21X1_967/C vdd OAI21X1
XOAI21X1_999 BUFX4_291/Y INVX1_154/Y OAI21X1_999/C gnd OAI21X1_999/Y vdd OAI21X1
XFILL_3_DFFPOSX1_649 gnd vdd FILL
XOAI21X1_977 BUFX4_297/Y INVX1_143/Y OAI21X1_977/C gnd OAI21X1_977/Y vdd OAI21X1
XOAI21X1_988 BUFX4_130/Y BUFX4_82/A BUFX2_387/A gnd OAI21X1_989/C vdd OAI21X1
XOAI21X1_1290 OAI21X1_1290/A NOR2X1_195/Y OAI21X1_1290/C gnd OAI21X1_1290/Y vdd OAI21X1
XDFFPOSX1_880 BUFX2_191/A CLKBUF1_12/Y OAI21X1_1231/Y gnd vdd DFFPOSX1
XDFFPOSX1_891 BUFX2_140/A CLKBUF1_35/Y OAI21X1_1263/Y gnd vdd DFFPOSX1
XINVX2_30 bundleStartMajId_i[18] gnd INVX2_30/Y vdd INVX2
XFILL_0_OAI21X1_290 gnd vdd FILL
XINVX2_63 bundleAddress_i[53] gnd INVX2_63/Y vdd INVX2
XFILL_1_OAI21X1_472 gnd vdd FILL
XFILL_1_OAI21X1_461 gnd vdd FILL
XINVX2_41 NOR2X1_5/Y gnd NOR2X1_6/B vdd INVX2
XFILL_1_OAI21X1_450 gnd vdd FILL
XFILL_7_0_1 gnd vdd FILL
XINVX2_52 INVX2_52/A gnd INVX2_52/Y vdd INVX2
XINVX2_96 INVX2_96/A gnd INVX2_96/Y vdd INVX2
XINVX2_74 bundleAddress_i[31] gnd INVX2_74/Y vdd INVX2
XFILL_1_OAI21X1_494 gnd vdd FILL
XINVX2_85 bundleAddress_i[11] gnd INVX2_85/Y vdd INVX2
XFILL_1_OAI21X1_483 gnd vdd FILL
XFILL_0_AOI21X1_4 gnd vdd FILL
XFILL_15_15_0 gnd vdd FILL
XFILL_2_OAI21X1_687 gnd vdd FILL
XFILL_2_OAI21X1_698 gnd vdd FILL
XFILL_2_DFFPOSX1_217 gnd vdd FILL
XFILL_2_DFFPOSX1_228 gnd vdd FILL
XBUFX2_326 BUFX2_326/A gnd instr3_o[30] vdd BUFX2
XBUFX2_315 BUFX2_315/A gnd instr2_o[2] vdd BUFX2
XBUFX2_304 BUFX2_304/A gnd instr2_o[12] vdd BUFX2
XFILL_2_DFFPOSX1_206 gnd vdd FILL
XBUFX2_348 BUFX2_348/A gnd instr3_o[28] vdd BUFX2
XFILL_2_DFFPOSX1_239 gnd vdd FILL
XBUFX2_359 BUFX2_359/A gnd instr4_o[21] vdd BUFX2
XFILL_5_DFFPOSX1_17 gnd vdd FILL
XBUFX2_337 BUFX2_337/A gnd instr3_o[29] vdd BUFX2
XFILL_5_DFFPOSX1_28 gnd vdd FILL
XFILL_5_DFFPOSX1_39 gnd vdd FILL
XFILL_1_INVX4_41 gnd vdd FILL
XFILL_1_BUFX4_220 gnd vdd FILL
XFILL_1_BUFX4_231 gnd vdd FILL
XOAI21X1_15 INVX2_153/Y BUFX4_219/Y OAI21X1_15/C gnd OAI21X1_15/Y vdd OAI21X1
XOAI21X1_26 INVX2_164/Y BUFX4_187/Y OAI21X1_26/C gnd OAI21X1_26/Y vdd OAI21X1
XFILL_1_BUFX4_253 gnd vdd FILL
XOAI21X1_59 INVX2_197/Y BUFX4_219/Y OAI21X1_59/C gnd OAI21X1_59/Y vdd OAI21X1
XFILL_1_BUFX4_242 gnd vdd FILL
XFILL_1_BUFX4_264 gnd vdd FILL
XOAI21X1_48 INVX2_186/Y BUFX4_190/Y OAI21X1_48/C gnd OAI21X1_48/Y vdd OAI21X1
XOAI21X1_37 INVX2_175/Y BUFX4_201/Y OAI21X1_37/C gnd OAI21X1_37/Y vdd OAI21X1
XFILL_0_DFFPOSX1_690 gnd vdd FILL
XFILL_1_BUFX4_297 gnd vdd FILL
XFILL_1_BUFX4_286 gnd vdd FILL
XFILL_1_BUFX4_275 gnd vdd FILL
XFILL_0_DFFPOSX1_13 gnd vdd FILL
XFILL_0_DFFPOSX1_24 gnd vdd FILL
XFILL_2_XNOR2X1_2 gnd vdd FILL
XFILL_0_DFFPOSX1_35 gnd vdd FILL
XFILL_0_DFFPOSX1_68 gnd vdd FILL
XFILL_0_DFFPOSX1_57 gnd vdd FILL
XFILL_0_DFFPOSX1_46 gnd vdd FILL
XFILL_33_16_0 gnd vdd FILL
XFILL_0_DFFPOSX1_79 gnd vdd FILL
XFILL_2_DFFPOSX1_751 gnd vdd FILL
XFILL_2_DFFPOSX1_740 gnd vdd FILL
XFILL_35_7_0 gnd vdd FILL
XFILL_2_OAI21X1_1172 gnd vdd FILL
XBUFX2_860 BUFX2_860/A gnd tid2_o[37] vdd BUFX2
XBUFX2_871 BUFX2_871/A gnd tid2_o[27] vdd BUFX2
XFILL_2_DFFPOSX1_773 gnd vdd FILL
XFILL_2_DFFPOSX1_762 gnd vdd FILL
XBUFX2_882 BUFX2_882/A gnd tid2_o[17] vdd BUFX2
XFILL_2_DFFPOSX1_784 gnd vdd FILL
XBUFX2_893 BUFX2_893/A gnd tid2_o[7] vdd BUFX2
XFILL_0_NOR2X1_211 gnd vdd FILL
XFILL_0_NOR2X1_222 gnd vdd FILL
XFILL_0_NOR2X1_200 gnd vdd FILL
XFILL_2_DFFPOSX1_795 gnd vdd FILL
XFILL_0_NOR2X1_233 gnd vdd FILL
XOAI21X1_229 INVX2_160/Y BUFX4_293/Y OAI21X1_229/C gnd OAI21X1_229/Y vdd OAI21X1
XOAI21X1_218 BUFX4_156/Y BUFX4_43/Y BUFX2_1032/A gnd OAI21X1_219/C vdd OAI21X1
XOAI21X1_207 INVX2_149/Y BUFX4_300/Y OAI21X1_207/C gnd OAI21X1_207/Y vdd OAI21X1
XFILL_6_DFFPOSX1_9 gnd vdd FILL
XFILL_3_CLKBUF1_2 gnd vdd FILL
XDFFPOSX1_121 BUFX2_791/A CLKBUF1_39/Y OAI21X1_1795/Y gnd vdd DFFPOSX1
XAND2X2_29 AND2X2_29/A AND2X2_29/B gnd OR2X2_20/A vdd AND2X2
XDFFPOSX1_110 BUFX2_779/A CLKBUF1_2/Y OAI21X1_1784/Y gnd vdd DFFPOSX1
XAND2X2_18 NOR2X1_4/Y INVX2_52/A gnd AND2X2_18/Y vdd AND2X2
XFILL_1_DFFPOSX1_330 gnd vdd FILL
XDFFPOSX1_154 BUFX2_827/A CLKBUF1_98/Y OAI21X1_1828/Y gnd vdd DFFPOSX1
XDFFPOSX1_143 BUFX2_815/A CLKBUF1_8/Y OAI21X1_1817/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_341 gnd vdd FILL
XDFFPOSX1_132 BUFX2_803/A CLKBUF1_66/Y OAI21X1_1806/Y gnd vdd DFFPOSX1
XFILL_38_15_0 gnd vdd FILL
XDFFPOSX1_198 BUFX2_869/A CLKBUF1_57/Y OAI21X1_42/Y gnd vdd DFFPOSX1
XDFFPOSX1_176 BUFX2_845/A CLKBUF1_99/Y OAI21X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_187 BUFX2_857/A CLKBUF1_42/Y OAI21X1_31/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_374 gnd vdd FILL
XFILL_0_NOR3X1_8 gnd vdd FILL
XFILL_1_DFFPOSX1_352 gnd vdd FILL
XNAND2X1_202 NOR2X1_16/Y NOR2X1_22/Y gnd NOR3X1_9/C vdd NAND2X1
XDFFPOSX1_165 NAND2X1_9/A CLKBUF1_62/Y OAI21X1_9/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_363 gnd vdd FILL
XNAND2X1_213 BUFX2_489/A BUFX4_213/Y gnd OAI21X1_456/C vdd NAND2X1
XNAND2X1_235 bundleStartMajId_i[14] NOR2X1_43/Y gnd OAI21X1_476/A vdd NAND2X1
XNAND2X1_224 bundleStartMajId_i[21] NOR2X1_37/B gnd XNOR2X1_19/A vdd NAND2X1
XFILL_1_DFFPOSX1_396 gnd vdd FILL
XFILL_1_DFFPOSX1_385 gnd vdd FILL
XFILL_4_DFFPOSX1_812 gnd vdd FILL
XNAND2X1_257 BUFX2_512/A BUFX4_213/Y gnd OAI21X1_492/C vdd NAND2X1
XNAND2X1_268 bundleStartMajId_i[60] INVX1_24/Y gnd INVX1_25/A vdd NAND2X1
XNAND2X1_246 BUFX2_506/A BUFX4_182/Y gnd OAI21X1_481/C vdd NAND2X1
XFILL_4_DFFPOSX1_801 gnd vdd FILL
XFILL_4_DFFPOSX1_856 gnd vdd FILL
XFILL_4_DFFPOSX1_823 gnd vdd FILL
XFILL_4_DFFPOSX1_834 gnd vdd FILL
XNAND2X1_279 NOR2X1_67/Y AND2X2_13/Y gnd OR2X2_6/A vdd NAND2X1
XFILL_4_DFFPOSX1_845 gnd vdd FILL
XFILL_4_DFFPOSX1_889 gnd vdd FILL
XFILL_4_DFFPOSX1_878 gnd vdd FILL
XFILL_4_DFFPOSX1_867 gnd vdd FILL
XFILL_26_7_0 gnd vdd FILL
XFILL_0_OAI21X1_7 gnd vdd FILL
XFILL_1_7_0 gnd vdd FILL
XFILL_4_CLKBUF1_90 gnd vdd FILL
XFILL_1_BUFX2_702 gnd vdd FILL
XFILL_1_BUFX2_713 gnd vdd FILL
XFILL_0_BUFX2_72 gnd vdd FILL
XFILL_0_BUFX2_61 gnd vdd FILL
XFILL_0_BUFX2_50 gnd vdd FILL
XFILL_1_BUFX2_746 gnd vdd FILL
XFILL_0_BUFX2_83 gnd vdd FILL
XFILL_0_BUFX2_94 gnd vdd FILL
XFILL_1_BUFX2_757 gnd vdd FILL
XFILL_3_DFFPOSX1_413 gnd vdd FILL
XFILL_1_NOR2X1_97 gnd vdd FILL
XFILL_0_BUFX4_309 gnd vdd FILL
XOAI21X1_741 OAI21X1_741/A BUFX4_295/Y OAI21X1_741/C gnd OAI21X1_741/Y vdd OAI21X1
XFILL_1_NOR2X1_75 gnd vdd FILL
XFILL_3_DFFPOSX1_402 gnd vdd FILL
XOAI21X1_730 NOR2X1_108/B INVX4_10/Y INVX4_11/Y gnd OAI21X1_731/C vdd OAI21X1
XOAI21X1_763 OAI21X1_763/A BUFX4_300/Y OAI21X1_763/C gnd OAI21X1_763/Y vdd OAI21X1
XOAI21X1_785 BUFX4_145/Y BUFX4_76/Y BUFX2_624/A gnd OAI21X1_786/C vdd OAI21X1
XOAI21X1_774 XNOR2X1_52/Y BUFX4_299/Y OAI21X1_774/C gnd OAI21X1_774/Y vdd OAI21X1
XOAI21X1_752 INVX2_43/Y OR2X2_15/A OAI21X1_752/C gnd OAI21X1_754/A vdd OAI21X1
XFILL_3_DFFPOSX1_424 gnd vdd FILL
XFILL_3_DFFPOSX1_435 gnd vdd FILL
XFILL_3_DFFPOSX1_446 gnd vdd FILL
XFILL_3_DFFPOSX1_479 gnd vdd FILL
XOAI21X1_796 OAI21X1_796/A BUFX4_289/Y OAI21X1_796/C gnd OAI21X1_796/Y vdd OAI21X1
XFILL_3_DFFPOSX1_468 gnd vdd FILL
XFILL_3_DFFPOSX1_457 gnd vdd FILL
XFILL_6_DFFPOSX1_906 gnd vdd FILL
XFILL_6_DFFPOSX1_917 gnd vdd FILL
XFILL_6_DFFPOSX1_928 gnd vdd FILL
XFILL_6_DFFPOSX1_939 gnd vdd FILL
XFILL_9_8_0 gnd vdd FILL
XFILL_1_OAI21X1_280 gnd vdd FILL
XFILL_1_OAI21X1_291 gnd vdd FILL
XFILL_2_OAI21X1_495 gnd vdd FILL
XBUFX2_101 BUFX2_101/A gnd addr2_o[22] vdd BUFX2
XFILL_2_XNOR2X1_31 gnd vdd FILL
XFILL_2_XNOR2X1_20 gnd vdd FILL
XFILL_2_XNOR2X1_64 gnd vdd FILL
XBUFX2_134 BUFX2_134/A gnd addr3_o[50] vdd BUFX2
XFILL_2_XNOR2X1_53 gnd vdd FILL
XBUFX2_123 BUFX2_123/A gnd addr2_o[2] vdd BUFX2
XFILL_17_7_0 gnd vdd FILL
XFILL_0_NAND2X1_509 gnd vdd FILL
XFILL_2_XNOR2X1_42 gnd vdd FILL
XBUFX2_112 BUFX2_112/A gnd addr2_o[12] vdd BUFX2
XFILL_2_XNOR2X1_75 gnd vdd FILL
XBUFX2_156 BUFX2_156/A gnd addr3_o[30] vdd BUFX2
XBUFX2_167 BUFX2_167/A gnd addr3_o[20] vdd BUFX2
XFILL_2_XNOR2X1_97 gnd vdd FILL
XBUFX2_178 BUFX2_178/A gnd addr3_o[10] vdd BUFX2
XFILL_2_XNOR2X1_86 gnd vdd FILL
XBUFX2_145 MUX2X1_2/B gnd addr3_o[40] vdd BUFX2
XFILL_1_NAND2X1_8 gnd vdd FILL
XFILL_6_DFFPOSX1_18 gnd vdd FILL
XFILL_6_DFFPOSX1_29 gnd vdd FILL
XBUFX2_189 BUFX2_189/A gnd addr3_o[0] vdd BUFX2
XFILL_5_DFFPOSX1_507 gnd vdd FILL
XFILL_5_DFFPOSX1_518 gnd vdd FILL
XFILL_5_DFFPOSX1_529 gnd vdd FILL
XFILL_22_13_1 gnd vdd FILL
XBUFX2_1015 BUFX2_1015/A gnd tid4_o[13] vdd BUFX2
XBUFX2_1026 BUFX2_1026/A gnd tid4_o[3] vdd BUFX2
XBUFX2_1004 BUFX2_1004/A gnd tid4_o[23] vdd BUFX2
XFILL_3_DFFPOSX1_980 gnd vdd FILL
XFILL_3_DFFPOSX1_991 gnd vdd FILL
XFILL_1_DFFPOSX1_14 gnd vdd FILL
XCLKBUF1_16 BUFX4_86/Y gnd CLKBUF1_16/Y vdd CLKBUF1
XCLKBUF1_27 BUFX4_92/Y gnd CLKBUF1_27/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_108 gnd vdd FILL
XCLKBUF1_38 BUFX4_89/Y gnd CLKBUF1_38/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_119 gnd vdd FILL
XFILL_1_DFFPOSX1_36 gnd vdd FILL
XFILL_1_DFFPOSX1_47 gnd vdd FILL
XFILL_1_DFFPOSX1_25 gnd vdd FILL
XCLKBUF1_49 BUFX4_92/Y gnd CLKBUF1_49/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_69 gnd vdd FILL
XFILL_1_DFFPOSX1_58 gnd vdd FILL
XBUFX4_70 BUFX4_75/A gnd BUFX4_70/Y vdd BUFX4
XBUFX4_92 clock_i gnd BUFX4_92/Y vdd BUFX4
XBUFX4_81 BUFX4_81/A gnd BUFX4_81/Y vdd BUFX4
XFILL_0_OAI21X1_1825 gnd vdd FILL
XFILL_0_OAI21X1_1803 gnd vdd FILL
XFILL_0_OAI21X1_1814 gnd vdd FILL
XBUFX2_690 BUFX2_690/A gnd pid2_o[14] vdd BUFX2
XFILL_2_DFFPOSX1_592 gnd vdd FILL
XFILL_2_DFFPOSX1_570 gnd vdd FILL
XFILL_2_DFFPOSX1_581 gnd vdd FILL
XFILL_27_12_1 gnd vdd FILL
XFILL_2_AOI21X1_20 gnd vdd FILL
XFILL_2_AOI21X1_31 gnd vdd FILL
XFILL_1_DFFPOSX1_171 gnd vdd FILL
XFILL_1_DFFPOSX1_182 gnd vdd FILL
XFILL_1_DFFPOSX1_160 gnd vdd FILL
XXNOR2X1_2 XNOR2X1_2/A INVX4_4/Y gnd XNOR2X1_2/Y vdd XNOR2X1
XFILL_2_AOI21X1_64 gnd vdd FILL
XFILL_1_DFFPOSX1_193 gnd vdd FILL
XFILL_4_DFFPOSX1_620 gnd vdd FILL
XFILL_4_DFFPOSX1_631 gnd vdd FILL
XFILL_4_DFFPOSX1_664 gnd vdd FILL
XFILL_4_DFFPOSX1_642 gnd vdd FILL
XFILL_4_DFFPOSX1_653 gnd vdd FILL
XFILL_4_DFFPOSX1_675 gnd vdd FILL
XFILL_2_13_1 gnd vdd FILL
XFILL_4_DFFPOSX1_697 gnd vdd FILL
XFILL_4_DFFPOSX1_686 gnd vdd FILL
XFILL_1_BUFX2_510 gnd vdd FILL
XFILL_0_BUFX4_106 gnd vdd FILL
XFILL_1_BUFX2_543 gnd vdd FILL
XFILL_1_BUFX2_554 gnd vdd FILL
XINVX1_2 bundleStartMajId_i[29] gnd INVX1_2/Y vdd INVX1
XFILL_0_BUFX4_128 gnd vdd FILL
XFILL_3_DFFPOSX1_221 gnd vdd FILL
XFILL_0_BUFX4_117 gnd vdd FILL
XFILL_1_BUFX2_565 gnd vdd FILL
XFILL_3_DFFPOSX1_210 gnd vdd FILL
XFILL_1_BUFX2_587 gnd vdd FILL
XFILL_1_INVX1_64 gnd vdd FILL
XFILL_0_BUFX4_139 gnd vdd FILL
XFILL_3_DFFPOSX1_232 gnd vdd FILL
XFILL_3_DFFPOSX1_254 gnd vdd FILL
XFILL_3_DFFPOSX1_243 gnd vdd FILL
XOAI21X1_571 OAI21X1_571/A BUFX4_147/Y OAI21X1_571/C gnd OAI21X1_571/Y vdd OAI21X1
XFILL_1_BUFX2_598 gnd vdd FILL
XOAI21X1_582 OR2X2_6/Y NOR2X1_74/A INVX2_24/Y gnd OAI21X1_582/Y vdd OAI21X1
XFILL_1_OAI21X1_1509 gnd vdd FILL
XOAI21X1_593 BUFX4_7/Y BUFX4_372/Y BUFX2_550/A gnd OAI21X1_594/C vdd OAI21X1
XOAI21X1_560 BUFX4_10/A BUFX4_337/Y BUFX2_536/A gnd OAI21X1_561/C vdd OAI21X1
XFILL_3_DFFPOSX1_276 gnd vdd FILL
XFILL_1_BUFX2_28 gnd vdd FILL
XFILL_3_DFFPOSX1_265 gnd vdd FILL
XFILL_1_BUFX2_39 gnd vdd FILL
XFILL_3_DFFPOSX1_287 gnd vdd FILL
XFILL_3_DFFPOSX1_298 gnd vdd FILL
XFILL_5_DFFPOSX1_6 gnd vdd FILL
XFILL_7_12_1 gnd vdd FILL
XFILL_2_OAI21X1_292 gnd vdd FILL
XFILL_0_NAND2X1_306 gnd vdd FILL
XFILL_0_NAND2X1_317 gnd vdd FILL
XFILL_0_NAND2X1_328 gnd vdd FILL
XFILL_0_NAND2X1_339 gnd vdd FILL
XFILL_32_5_0 gnd vdd FILL
XFILL_1_DFFPOSX1_1012 gnd vdd FILL
XFILL_1_CLKBUF1_100 gnd vdd FILL
XFILL_1_DFFPOSX1_1001 gnd vdd FILL
XFILL_5_DFFPOSX1_304 gnd vdd FILL
XFILL_5_DFFPOSX1_326 gnd vdd FILL
XFILL_5_DFFPOSX1_315 gnd vdd FILL
XFILL_1_DFFPOSX1_1023 gnd vdd FILL
XFILL_5_DFFPOSX1_337 gnd vdd FILL
XFILL_5_DFFPOSX1_348 gnd vdd FILL
XFILL_5_DFFPOSX1_359 gnd vdd FILL
XOAI21X1_1801 BUFX4_332/Y INVX2_173/Y NAND2X1_742/Y gnd OAI21X1_1801/Y vdd OAI21X1
XOAI21X1_1812 BUFX4_322/Y INVX2_184/Y NAND2X1_753/Y gnd OAI21X1_1812/Y vdd OAI21X1
XOAI21X1_1823 BUFX4_313/Y INVX2_195/Y NAND2X1_764/Y gnd OAI21X1_1823/Y vdd OAI21X1
XFILL_0_OAI21X1_812 gnd vdd FILL
XFILL_0_OAI21X1_823 gnd vdd FILL
XFILL_0_OAI21X1_801 gnd vdd FILL
XFILL_0_OAI21X1_845 gnd vdd FILL
XFILL_0_OAI21X1_834 gnd vdd FILL
XFILL_0_OAI21X1_856 gnd vdd FILL
XFILL_0_OAI21X1_867 gnd vdd FILL
XFILL_0_OAI21X1_889 gnd vdd FILL
XFILL_0_OAI21X1_878 gnd vdd FILL
XFILL_2_DFFPOSX1_37 gnd vdd FILL
XFILL_2_DFFPOSX1_26 gnd vdd FILL
XFILL_2_DFFPOSX1_15 gnd vdd FILL
XFILL_2_DFFPOSX1_59 gnd vdd FILL
XFILL_2_DFFPOSX1_48 gnd vdd FILL
XFILL_13_18_1 gnd vdd FILL
XFILL_0_OAI21X1_1600 gnd vdd FILL
XFILL_0_OAI21X1_1622 gnd vdd FILL
XFILL_0_OAI21X1_1633 gnd vdd FILL
XFILL_0_OAI21X1_1611 gnd vdd FILL
XFILL_0_OAI21X1_1677 gnd vdd FILL
XFILL_0_OAI21X1_1666 gnd vdd FILL
XFILL_23_5_0 gnd vdd FILL
XFILL_0_OAI21X1_1655 gnd vdd FILL
XFILL_0_OAI21X1_1644 gnd vdd FILL
XFILL_0_OAI21X1_1688 gnd vdd FILL
XFILL_0_OAI21X1_1699 gnd vdd FILL
XFILL_0_BUFX4_8 gnd vdd FILL
XFILL_5_DFFPOSX1_882 gnd vdd FILL
XFILL_5_DFFPOSX1_871 gnd vdd FILL
XFILL_5_DFFPOSX1_860 gnd vdd FILL
XFILL_5_DFFPOSX1_893 gnd vdd FILL
XFILL_4_DFFPOSX1_1005 gnd vdd FILL
XFILL_1_XNOR2X1_72 gnd vdd FILL
XFILL_1_XNOR2X1_50 gnd vdd FILL
XFILL_1_XNOR2X1_61 gnd vdd FILL
XFILL_4_DFFPOSX1_1027 gnd vdd FILL
XFILL_4_DFFPOSX1_1016 gnd vdd FILL
XFILL_1_XNOR2X1_83 gnd vdd FILL
XFILL_1_XNOR2X1_94 gnd vdd FILL
XFILL_18_17_1 gnd vdd FILL
XBUFX4_207 BUFX4_26/Y gnd BUFX4_207/Y vdd BUFX4
XBUFX4_218 BUFX4_23/Y gnd BUFX4_218/Y vdd BUFX4
XFILL_2_OAI21X1_1705 gnd vdd FILL
XFILL_6_6_0 gnd vdd FILL
XFILL_0_INVX2_117 gnd vdd FILL
XBUFX4_229 BUFX4_26/Y gnd BUFX4_229/Y vdd BUFX4
XFILL_4_DFFPOSX1_450 gnd vdd FILL
XFILL_2_OAI21X1_1749 gnd vdd FILL
XFILL_2_OAI21X1_1716 gnd vdd FILL
XFILL_4_DFFPOSX1_461 gnd vdd FILL
XFILL_0_INVX2_106 gnd vdd FILL
XFILL_4_DFFPOSX1_472 gnd vdd FILL
XFILL_0_INVX2_139 gnd vdd FILL
XFILL_4_DFFPOSX1_483 gnd vdd FILL
XFILL_0_INVX2_128 gnd vdd FILL
XFILL_12_13_0 gnd vdd FILL
XFILL_4_DFFPOSX1_494 gnd vdd FILL
XFILL_14_5_0 gnd vdd FILL
XFILL_0_INVX4_8 gnd vdd FILL
XFILL_1_BUFX2_362 gnd vdd FILL
XFILL_1_BUFX2_340 gnd vdd FILL
XFILL_1_BUFX2_351 gnd vdd FILL
XOAI21X1_1108 OAI21X1_1108/A AOI21X1_36/Y NAND2X1_473/Y gnd OAI21X1_1108/Y vdd OAI21X1
XOAI21X1_1119 OAI21X1_1119/A BUFX4_204/Y NAND2X1_483/Y gnd OAI21X1_1119/Y vdd OAI21X1
XFILL_1_BUFX2_395 gnd vdd FILL
XOAI21X1_390 BUFX4_356/Y INVX1_5/Y OAI21X1_390/C gnd OAI21X1_390/Y vdd OAI21X1
XFILL_1_OAI21X1_1339 gnd vdd FILL
XFILL_1_OAI21X1_1328 gnd vdd FILL
XFILL_1_OAI21X1_1306 gnd vdd FILL
XDFFPOSX1_709 BUFX2_347/A CLKBUF1_56/Y OAI21X1_967/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1317 gnd vdd FILL
XFILL_1_DFFPOSX1_907 gnd vdd FILL
XAND2X2_2 NOR2X1_7/Y AND2X2_2/B gnd AND2X2_2/Y vdd AND2X2
XFILL_0_OAI21X1_119 gnd vdd FILL
XFILL_0_OAI21X1_108 gnd vdd FILL
XFILL_1_DFFPOSX1_918 gnd vdd FILL
XFILL_1_DFFPOSX1_929 gnd vdd FILL
XFILL_6_DFFPOSX1_544 gnd vdd FILL
XFILL_6_DFFPOSX1_533 gnd vdd FILL
XFILL_36_18_1 gnd vdd FILL
XFILL_6_DFFPOSX1_555 gnd vdd FILL
XFILL_6_DFFPOSX1_566 gnd vdd FILL
XFILL_17_12_0 gnd vdd FILL
XFILL_6_DFFPOSX1_577 gnd vdd FILL
XFILL_6_DFFPOSX1_588 gnd vdd FILL
XFILL_0_BUFX4_18 gnd vdd FILL
XFILL_30_14_0 gnd vdd FILL
XFILL_0_BUFX4_29 gnd vdd FILL
XFILL_0_NAND2X1_125 gnd vdd FILL
XFILL_0_NAND2X1_114 gnd vdd FILL
XFILL_0_NAND2X1_103 gnd vdd FILL
XFILL_1_NAND2X1_307 gnd vdd FILL
XFILL_1_NAND2X1_329 gnd vdd FILL
XFILL_0_NAND2X1_158 gnd vdd FILL
XFILL_0_NAND2X1_136 gnd vdd FILL
XFILL_0_NAND2X1_147 gnd vdd FILL
XFILL_1_NAND2X1_318 gnd vdd FILL
XFILL_37_1 gnd vdd FILL
XFILL_0_INVX1_150 gnd vdd FILL
XFILL_0_DFFPOSX1_519 gnd vdd FILL
XFILL_1_AOI21X1_50 gnd vdd FILL
XFILL_0_INVX1_161 gnd vdd FILL
XFILL_0_DFFPOSX1_508 gnd vdd FILL
XFILL_0_INVX1_172 gnd vdd FILL
XFILL_0_NAND2X1_169 gnd vdd FILL
XFILL_0_INVX1_183 gnd vdd FILL
XFILL_1_AOI21X1_61 gnd vdd FILL
XFILL_0_INVX1_194 gnd vdd FILL
XFILL_5_DFFPOSX1_101 gnd vdd FILL
XFILL_5_DFFPOSX1_134 gnd vdd FILL
XFILL_5_DFFPOSX1_112 gnd vdd FILL
XFILL_2_CLKBUF1_101 gnd vdd FILL
XFILL_5_DFFPOSX1_123 gnd vdd FILL
XFILL_5_DFFPOSX1_178 gnd vdd FILL
XFILL_5_DFFPOSX1_156 gnd vdd FILL
XFILL_5_DFFPOSX1_145 gnd vdd FILL
XFILL_5_DFFPOSX1_167 gnd vdd FILL
XFILL_5_DFFPOSX1_189 gnd vdd FILL
XOAI21X1_1642 INVX2_145/Y BUFX4_197/Y NAND2X1_710/Y gnd DFFPOSX1_32/D vdd OAI21X1
XOAI21X1_1631 INVX2_134/Y BUFX4_220/Y NAND2X1_699/Y gnd DFFPOSX1_21/D vdd OAI21X1
XOAI21X1_1620 INVX2_123/Y BUFX4_217/Y NAND2X1_688/Y gnd DFFPOSX1_10/D vdd OAI21X1
XOAI21X1_1675 BUFX4_172/Y INVX2_131/Y OAI21X1_1675/C gnd DFFPOSX1_50/D vdd OAI21X1
XOAI21X1_1653 BUFX4_138/Y INVX2_120/Y OAI21X1_1653/C gnd DFFPOSX1_39/D vdd OAI21X1
XOAI21X1_1664 BUFX4_111/Y BUFX4_375/Y BUFX2_744/A gnd OAI21X1_1665/C vdd OAI21X1
XOAI21X1_1686 BUFX4_11/A BUFX4_339/Y BUFX2_726/A gnd OAI21X1_1687/C vdd OAI21X1
XFILL_1_OAI21X1_802 gnd vdd FILL
XOAI21X1_1697 BUFX4_147/Y INVX2_142/Y OAI21X1_1697/C gnd DFFPOSX1_61/D vdd OAI21X1
XFILL_0_OAI21X1_631 gnd vdd FILL
XFILL_0_OAI21X1_620 gnd vdd FILL
XFILL_0_OAI21X1_653 gnd vdd FILL
XFILL_1_OAI21X1_835 gnd vdd FILL
XFILL_1_OAI21X1_813 gnd vdd FILL
XFILL_1_OAI21X1_824 gnd vdd FILL
XFILL_0_OAI21X1_642 gnd vdd FILL
XFILL_0_OAI21X1_664 gnd vdd FILL
XFILL_1_OAI21X1_846 gnd vdd FILL
XFILL_1_OAI21X1_879 gnd vdd FILL
XFILL_35_13_0 gnd vdd FILL
XFILL_1_OAI21X1_868 gnd vdd FILL
XNAND3X1_29 AND2X2_7/A NOR2X1_105/Y NOR2X1_30/Y gnd NOR2X1_112/B vdd NAND3X1
XNAND3X1_18 NOR2X1_67/Y NOR2X1_69/Y AND2X2_14/Y gnd OR2X2_10/A vdd NAND3X1
XFILL_0_OAI21X1_697 gnd vdd FILL
XFILL_1_OAI21X1_857 gnd vdd FILL
XFILL_0_OAI21X1_686 gnd vdd FILL
XFILL_0_OAI21X1_675 gnd vdd FILL
XFILL_1_AND2X2_32 gnd vdd FILL
XFILL_1_AND2X2_21 gnd vdd FILL
XFILL_1_AND2X2_10 gnd vdd FILL
XFILL_3_DFFPOSX1_16 gnd vdd FILL
XNOR2X1_18 INVX4_10/Y INVX4_11/Y gnd INVX1_12/A vdd NOR2X1
XFILL_3_DFFPOSX1_27 gnd vdd FILL
XFILL_3_DFFPOSX1_38 gnd vdd FILL
XFILL_3_DFFPOSX1_49 gnd vdd FILL
XNOR2X1_29 INVX4_13/Y INVX2_24/Y gnd NOR2X1_29/Y vdd NOR2X1
XFILL_0_OAI21X1_1430 gnd vdd FILL
XFILL_0_NAND2X1_670 gnd vdd FILL
XFILL_0_OAI21X1_1441 gnd vdd FILL
XFILL_0_NAND2X1_681 gnd vdd FILL
XFILL_0_NAND2X1_692 gnd vdd FILL
XFILL_0_OAI21X1_1474 gnd vdd FILL
XFILL_0_OAI21X1_1463 gnd vdd FILL
XFILL_0_OAI21X1_1485 gnd vdd FILL
XFILL_0_OAI21X1_1452 gnd vdd FILL
XFILL_0_OAI21X1_1496 gnd vdd FILL
XFILL_4_DFFPOSX1_3 gnd vdd FILL
XFILL_0_BUFX2_5 gnd vdd FILL
XFILL_5_DFFPOSX1_690 gnd vdd FILL
XFILL_0_BUFX2_429 gnd vdd FILL
XFILL_0_BUFX2_418 gnd vdd FILL
XFILL_0_BUFX2_407 gnd vdd FILL
XFILL_0_NAND2X1_38 gnd vdd FILL
XFILL_0_NAND2X1_27 gnd vdd FILL
XFILL_2_OAI21X1_1557 gnd vdd FILL
XFILL_0_NAND2X1_16 gnd vdd FILL
XFILL_4_DFFPOSX1_280 gnd vdd FILL
XNOR2X1_119 bundleStartMajId_i[2] NOR2X1_119/B gnd NOR2X1_119/Y vdd NOR2X1
XFILL_2_OAI21X1_1579 gnd vdd FILL
XFILL_4_DFFPOSX1_291 gnd vdd FILL
XNOR2X1_108 INVX4_10/Y NOR2X1_108/B gnd INVX1_38/A vdd NOR2X1
XFILL_0_NAND2X1_49 gnd vdd FILL
XFILL_0_INVX2_5 gnd vdd FILL
XFILL_30_8_1 gnd vdd FILL
XFILL_1_BUFX2_192 gnd vdd FILL
XFILL_1_OAI21X1_1114 gnd vdd FILL
XFILL_1_OAI21X1_1103 gnd vdd FILL
XFILL_1_DFFPOSX1_715 gnd vdd FILL
XFILL_1_DFFPOSX1_704 gnd vdd FILL
XFILL_1_OAI21X1_1125 gnd vdd FILL
XFILL_1_OAI21X1_1147 gnd vdd FILL
XFILL_0_BUFX2_930 gnd vdd FILL
XFILL_0_BUFX2_952 gnd vdd FILL
XDFFPOSX1_528 BUFX2_560/A CLKBUF1_80/Y OAI21X1_614/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_941 gnd vdd FILL
XDFFPOSX1_506 BUFX2_536/A CLKBUF1_44/Y OAI21X1_561/Y gnd vdd DFFPOSX1
XDFFPOSX1_517 BUFX2_548/A CLKBUF1_48/Y OAI21X1_586/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1136 gnd vdd FILL
XFILL_0_BUFX2_985 gnd vdd FILL
XFILL_1_DFFPOSX1_737 gnd vdd FILL
XFILL_0_BUFX2_963 gnd vdd FILL
XFILL_1_DFFPOSX1_748 gnd vdd FILL
XDFFPOSX1_539 BUFX2_572/A CLKBUF1_84/Y OAI21X1_640/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1169 gnd vdd FILL
XFILL_1_OAI21X1_1158 gnd vdd FILL
XFILL_1_DFFPOSX1_726 gnd vdd FILL
XFILL_0_BUFX2_974 gnd vdd FILL
XFILL_0_BUFX2_996 gnd vdd FILL
XFILL_1_DFFPOSX1_759 gnd vdd FILL
XFILL_1_OAI21X1_109 gnd vdd FILL
XNAND2X1_609 bundleAddress_i[26] bundleAddress_i[25] gnd NOR2X1_200/B vdd NAND2X1
XFILL_6_DFFPOSX1_330 gnd vdd FILL
XFILL_6_DFFPOSX1_341 gnd vdd FILL
XNAND2X1_51 BUFX2_879/A BUFX4_193/Y gnd OAI21X1_51/C vdd NAND2X1
XNAND2X1_40 BUFX2_867/A BUFX4_215/Y gnd OAI21X1_40/C vdd NAND2X1
XFILL_38_9_1 gnd vdd FILL
XFILL_37_4_0 gnd vdd FILL
XNAND2X1_62 BUFX2_891/A BUFX4_208/Y gnd OAI21X1_62/C vdd NAND2X1
XNAND2X1_73 BUFX2_394/A BUFX4_321/Y gnd NAND2X1_73/Y vdd NAND2X1
XNAND2X1_84 BUFX2_397/A BUFX4_358/Y gnd NAND2X1_84/Y vdd NAND2X1
XNAND2X1_95 BUFX2_409/A BUFX4_337/Y gnd NAND2X1_95/Y vdd NAND2X1
XFILL_0_XNOR2X1_80 gnd vdd FILL
XFILL_0_XNOR2X1_91 gnd vdd FILL
XFILL_1_NAND2X1_137 gnd vdd FILL
XFILL_0_DFFPOSX1_305 gnd vdd FILL
XFILL_0_DFFPOSX1_316 gnd vdd FILL
XFILL_0_DFFPOSX1_327 gnd vdd FILL
XFILL_0_DFFPOSX1_338 gnd vdd FILL
XFILL_1_NAND2X1_148 gnd vdd FILL
XFILL_0_DFFPOSX1_349 gnd vdd FILL
XFILL_3_CLKBUF1_102 gnd vdd FILL
XFILL_21_8_1 gnd vdd FILL
XFILL_20_3_0 gnd vdd FILL
XFILL_24_10_1 gnd vdd FILL
XFILL_3_DFFPOSX1_809 gnd vdd FILL
XFILL_0_NOR3X1_12 gnd vdd FILL
XOAI21X1_1450 BUFX4_129/Y BUFX4_80/Y BUFX2_208/A gnd OAI21X1_1451/C vdd OAI21X1
XOAI21X1_1472 OR2X2_20/B BUFX4_50/Y BUFX2_217/A gnd OAI21X1_1473/C vdd OAI21X1
XOAI21X1_1461 OR2X2_20/B BUFX4_59/Y BUFX2_213/A gnd OAI21X1_1462/C vdd OAI21X1
XOAI21X1_1483 BUFX4_160/Y BUFX4_32/Y BUFX2_221/A gnd OAI21X1_1484/C vdd OAI21X1
XFILL_1_OAI21X1_1692 gnd vdd FILL
XFILL_1_OAI21X1_1681 gnd vdd FILL
XFILL_1_OAI21X1_1670 gnd vdd FILL
XFILL_1_OAI21X1_610 gnd vdd FILL
XFILL_1_OAI21X1_621 gnd vdd FILL
XOAI21X1_1494 INVX2_100/Y INVX1_223/A OAI21X1_1494/C gnd OAI21X1_1496/A vdd OAI21X1
XFILL_1_OAI21X1_654 gnd vdd FILL
XFILL_1_OAI21X1_643 gnd vdd FILL
XFILL_1_NOR2X1_226 gnd vdd FILL
XFILL_0_OAI21X1_472 gnd vdd FILL
XFILL_1_OAI21X1_632 gnd vdd FILL
XFILL_0_OAI21X1_461 gnd vdd FILL
XFILL_0_OAI21X1_483 gnd vdd FILL
XFILL_0_OAI21X1_450 gnd vdd FILL
XFILL_0_OAI21X1_494 gnd vdd FILL
XFILL_1_OAI21X1_665 gnd vdd FILL
XFILL_3_NOR3X1_5 gnd vdd FILL
XFILL_1_OAI21X1_687 gnd vdd FILL
XFILL_1_OAI21X1_676 gnd vdd FILL
XFILL_1_OAI21X1_698 gnd vdd FILL
XFILL_29_9_1 gnd vdd FILL
XFILL_28_4_0 gnd vdd FILL
XFILL_3_4_0 gnd vdd FILL
XFILL_4_9_1 gnd vdd FILL
XBUFX2_508 BUFX2_508/A gnd majID2_o[8] vdd BUFX2
XFILL_4_DFFPOSX1_39 gnd vdd FILL
XFILL_4_DFFPOSX1_17 gnd vdd FILL
XBUFX2_519 BUFX2_519/A gnd majID2_o[55] vdd BUFX2
XFILL_4_DFFPOSX1_28 gnd vdd FILL
XFILL_1_NAND2X1_660 gnd vdd FILL
XFILL_0_OAI21X1_1260 gnd vdd FILL
XFILL_1_NAND2X1_671 gnd vdd FILL
XFILL_0_OAI21X1_1293 gnd vdd FILL
XFILL_0_OAI21X1_1282 gnd vdd FILL
XFILL_0_DFFPOSX1_850 gnd vdd FILL
XFILL_0_OAI21X1_1271 gnd vdd FILL
XFILL_0_DFFPOSX1_861 gnd vdd FILL
XFILL_0_DFFPOSX1_883 gnd vdd FILL
XFILL_0_DFFPOSX1_872 gnd vdd FILL
XFILL_26_18_0 gnd vdd FILL
XDFFPOSX1_1002 BUFX2_391/A CLKBUF1_35/Y OAI21X1_1578/Y gnd vdd DFFPOSX1
XFILL_0_DFFPOSX1_894 gnd vdd FILL
XFILL_12_8_1 gnd vdd FILL
XFILL_11_3_0 gnd vdd FILL
XDFFPOSX1_1013 BUFX2_680/A CLKBUF1_57/Y OAI21X1_1590/Y gnd vdd DFFPOSX1
XDFFPOSX1_1024 BUFX2_662/A CLKBUF1_42/Y OAI21X1_1601/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_204 gnd vdd FILL
XFILL_0_BUFX2_237 gnd vdd FILL
XFILL_0_BUFX2_215 gnd vdd FILL
XFILL_0_BUFX2_226 gnd vdd FILL
XFILL_0_BUFX2_248 gnd vdd FILL
XFILL_0_BUFX2_259 gnd vdd FILL
XFILL_2_DFFPOSX1_900 gnd vdd FILL
XFILL_19_4_0 gnd vdd FILL
XFILL_4_10_1 gnd vdd FILL
XFILL_2_DFFPOSX1_922 gnd vdd FILL
XFILL_2_DFFPOSX1_933 gnd vdd FILL
XFILL_2_DFFPOSX1_911 gnd vdd FILL
XFILL_2_DFFPOSX1_944 gnd vdd FILL
XFILL_2_DFFPOSX1_966 gnd vdd FILL
XFILL_2_DFFPOSX1_955 gnd vdd FILL
XFILL_2_DFFPOSX1_999 gnd vdd FILL
XFILL_2_DFFPOSX1_977 gnd vdd FILL
XFILL_2_DFFPOSX1_988 gnd vdd FILL
XFILL_3_XNOR2X1_13 gnd vdd FILL
XDFFPOSX1_303 BUFX2_972/A CLKBUF1_14/Y OAI21X1_223/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_57 gnd vdd FILL
XFILL_3_XNOR2X1_46 gnd vdd FILL
XFILL_3_XNOR2X1_35 gnd vdd FILL
XFILL_0_BUFX2_760 gnd vdd FILL
XDFFPOSX1_336 BUFX2_1008/A CLKBUF1_7/Y OAI21X1_289/Y gnd vdd DFFPOSX1
XDFFPOSX1_325 BUFX2_996/A CLKBUF1_98/Y OAI21X1_267/Y gnd vdd DFFPOSX1
XDFFPOSX1_314 BUFX2_984/A CLKBUF1_97/Y OAI21X1_245/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_512 gnd vdd FILL
XDFFPOSX1_347 BUFX2_1020/A CLKBUF1_4/Y OAI21X1_311/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_501 gnd vdd FILL
XFILL_1_DFFPOSX1_523 gnd vdd FILL
XFILL_3_XNOR2X1_68 gnd vdd FILL
XFILL_1_DFFPOSX1_545 gnd vdd FILL
XFILL_0_BUFX2_793 gnd vdd FILL
XFILL_1_DFFPOSX1_534 gnd vdd FILL
XDFFPOSX1_358 BUFX2_405/A CLKBUF1_80/Y OAI21X1_330/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_771 gnd vdd FILL
XFILL_0_BUFX2_782 gnd vdd FILL
XFILL_1_DFFPOSX1_556 gnd vdd FILL
XDFFPOSX1_369 BUFX2_398/A CLKBUF1_46/Y OAI21X1_341/Y gnd vdd DFFPOSX1
XNAND2X1_417 BUFX2_8/A BUFX4_385/Y gnd NAND2X1_417/Y vdd NAND2X1
XNAND2X1_406 BUFX2_35/A BUFX4_347/Y gnd NAND2X1_406/Y vdd NAND2X1
XFILL_1_DFFPOSX1_578 gnd vdd FILL
XFILL_1_DFFPOSX1_567 gnd vdd FILL
XFILL_1_DFFPOSX1_589 gnd vdd FILL
XNAND2X1_428 BUFX2_20/A BUFX4_317/Y gnd NAND2X1_428/Y vdd NAND2X1
XNAND2X1_439 BUFX2_32/A BUFX4_370/Y gnd NAND2X1_439/Y vdd NAND2X1
XFILL_6_DFFPOSX1_182 gnd vdd FILL
XFILL_6_18_0 gnd vdd FILL
XFILL_6_DFFPOSX1_193 gnd vdd FILL
XFILL_10_16_1 gnd vdd FILL
XFILL_0_DFFPOSX1_102 gnd vdd FILL
XFILL_0_DFFPOSX1_113 gnd vdd FILL
XFILL_0_DFFPOSX1_157 gnd vdd FILL
XFILL_0_DFFPOSX1_124 gnd vdd FILL
XFILL_0_DFFPOSX1_135 gnd vdd FILL
XFILL_0_DFFPOSX1_146 gnd vdd FILL
XFILL_0_DFFPOSX1_179 gnd vdd FILL
XFILL_0_DFFPOSX1_168 gnd vdd FILL
XFILL_1_BUFX2_928 gnd vdd FILL
XFILL_1_BUFX2_939 gnd vdd FILL
XOAI21X1_923 BUFX4_141/Y INVX1_116/Y OAI21X1_923/C gnd OAI21X1_923/Y vdd OAI21X1
XOAI21X1_934 BUFX4_7/A BUFX4_315/Y BUFX2_330/A gnd OAI21X1_935/C vdd OAI21X1
XOAI21X1_901 INVX1_102/Y BUFX4_196/Y OAI21X1_901/C gnd OAI21X1_901/Y vdd OAI21X1
XOAI21X1_912 BUFX4_102/Y BUFX4_315/Y BUFX2_337/A gnd OAI21X1_913/C vdd OAI21X1
XOAI21X1_956 BUFX4_247/Y BUFX4_329/Y BUFX2_342/A gnd OAI21X1_957/C vdd OAI21X1
XOAI21X1_945 BUFX4_143/Y INVX1_127/Y OAI21X1_945/C gnd OAI21X1_945/Y vdd OAI21X1
XFILL_3_DFFPOSX1_606 gnd vdd FILL
XFILL_3_DFFPOSX1_617 gnd vdd FILL
XFILL_3_DFFPOSX1_628 gnd vdd FILL
XOAI21X1_967 BUFX4_153/Y INVX1_138/Y OAI21X1_967/C gnd OAI21X1_967/Y vdd OAI21X1
XOAI21X1_978 BUFX4_164/Y BUFX4_44/Y BUFX2_380/A gnd OAI21X1_979/C vdd OAI21X1
XFILL_3_DFFPOSX1_639 gnd vdd FILL
XOAI21X1_989 BUFX4_295/Y INVX1_149/Y OAI21X1_989/C gnd OAI21X1_989/Y vdd OAI21X1
XOAI21X1_1291 BUFX4_106/Y BUFX4_318/Y BUFX2_153/A gnd OAI21X1_1292/C vdd OAI21X1
XOAI21X1_1280 AND2X2_27/Y OAI21X1_1280/B OAI21X1_1280/C gnd OAI21X1_1280/Y vdd OAI21X1
XDFFPOSX1_881 BUFX2_192/A CLKBUF1_74/Y OAI21X1_1233/Y gnd vdd DFFPOSX1
XDFFPOSX1_870 BUFX2_124/A CLKBUF1_97/Y OAI21X1_1205/Y gnd vdd DFFPOSX1
XDFFPOSX1_892 BUFX2_142/A CLKBUF1_34/Y OAI21X1_1267/Y gnd vdd DFFPOSX1
XINVX2_20 bundleStartMajId_i[43] gnd INVX2_20/Y vdd INVX2
XFILL_0_OAI21X1_291 gnd vdd FILL
XFILL_2_OAI21X1_633 gnd vdd FILL
XINVX2_53 INVX2_53/A gnd INVX2_53/Y vdd INVX2
XFILL_1_OAI21X1_462 gnd vdd FILL
XINVX2_31 bundleStartMajId_i[17] gnd INVX2_31/Y vdd INVX2
XINVX2_42 OR2X2_4/A gnd INVX2_42/Y vdd INVX2
XFILL_0_OAI21X1_280 gnd vdd FILL
XFILL_1_OAI21X1_451 gnd vdd FILL
XFILL_1_OAI21X1_440 gnd vdd FILL
XINVX2_64 bundleAddress_i[51] gnd INVX2_64/Y vdd INVX2
XINVX2_75 bundleAddress_i[30] gnd INVX2_75/Y vdd INVX2
XFILL_1_OAI21X1_495 gnd vdd FILL
XFILL_1_OAI21X1_473 gnd vdd FILL
XINVX2_97 INVX2_97/A gnd INVX2_97/Y vdd INVX2
XINVX2_86 bundleAddress_i[10] gnd INVX2_86/Y vdd INVX2
XFILL_1_OAI21X1_484 gnd vdd FILL
XFILL_15_15_1 gnd vdd FILL
XBUFX2_327 BUFX2_327/A gnd instr3_o[21] vdd BUFX2
XFILL_2_DFFPOSX1_218 gnd vdd FILL
XFILL_2_DFFPOSX1_207 gnd vdd FILL
XBUFX2_305 BUFX2_305/A gnd instr2_o[29] vdd BUFX2
XFILL_0_AOI21X1_5 gnd vdd FILL
XBUFX2_316 BUFX2_316/A gnd instr2_o[28] vdd BUFX2
XBUFX2_338 BUFX2_338/A gnd instr3_o[11] vdd BUFX2
XFILL_5_DFFPOSX1_18 gnd vdd FILL
XFILL_2_DFFPOSX1_229 gnd vdd FILL
XBUFX2_349 BUFX2_349/A gnd instr3_o[1] vdd BUFX2
XFILL_1_INVX4_20 gnd vdd FILL
XFILL_5_DFFPOSX1_29 gnd vdd FILL
XFILL_1_INVX4_31 gnd vdd FILL
XFILL_1_BUFX4_210 gnd vdd FILL
XFILL_1_BUFX4_221 gnd vdd FILL
XOAI21X1_16 INVX2_154/Y BUFX4_237/Y OAI21X1_16/C gnd OAI21X1_16/Y vdd OAI21X1
XOAI21X1_38 INVX2_176/Y OAI21X1_8/B OAI21X1_38/C gnd OAI21X1_38/Y vdd OAI21X1
XOAI21X1_27 INVX2_165/Y BUFX4_200/Y OAI21X1_27/C gnd OAI21X1_27/Y vdd OAI21X1
XFILL_1_BUFX4_243 gnd vdd FILL
XFILL_1_BUFX4_254 gnd vdd FILL
XOAI21X1_49 INVX2_187/Y BUFX4_188/Y OAI21X1_49/C gnd OAI21X1_49/Y vdd OAI21X1
XFILL_1_BUFX4_232 gnd vdd FILL
XFILL_0_OAI21X1_1090 gnd vdd FILL
XFILL_0_DFFPOSX1_691 gnd vdd FILL
XFILL_0_DFFPOSX1_680 gnd vdd FILL
XFILL_1_BUFX4_265 gnd vdd FILL
XFILL_1_BUFX4_298 gnd vdd FILL
XFILL_1_BUFX4_287 gnd vdd FILL
XFILL_1_BUFX4_276 gnd vdd FILL
XFILL_0_DFFPOSX1_25 gnd vdd FILL
XFILL_0_DFFPOSX1_14 gnd vdd FILL
XFILL_0_DFFPOSX1_58 gnd vdd FILL
XFILL_0_DFFPOSX1_36 gnd vdd FILL
XFILL_0_DFFPOSX1_47 gnd vdd FILL
XFILL_2_XNOR2X1_3 gnd vdd FILL
XFILL_0_DFFPOSX1_69 gnd vdd FILL
XFILL_33_16_1 gnd vdd FILL
XFILL_2_BUFX4_92 gnd vdd FILL
XFILL_14_10_0 gnd vdd FILL
XFILL_2_OAI21X1_1140 gnd vdd FILL
XFILL_2_DFFPOSX1_741 gnd vdd FILL
XFILL_35_7_1 gnd vdd FILL
XFILL_2_DFFPOSX1_730 gnd vdd FILL
XBUFX2_861 BUFX2_861/A gnd tid2_o[36] vdd BUFX2
XBUFX2_850 BUFX2_850/A gnd tid2_o[46] vdd BUFX2
XFILL_2_DFFPOSX1_752 gnd vdd FILL
XFILL_34_2_0 gnd vdd FILL
XFILL_2_DFFPOSX1_774 gnd vdd FILL
XBUFX2_872 BUFX2_872/A gnd tid2_o[26] vdd BUFX2
XFILL_2_DFFPOSX1_763 gnd vdd FILL
XFILL_2_OAI21X1_1184 gnd vdd FILL
XBUFX2_883 BUFX2_883/A gnd tid2_o[16] vdd BUFX2
XBUFX2_894 BUFX2_894/A gnd tid2_o[6] vdd BUFX2
XFILL_0_NOR2X1_212 gnd vdd FILL
XFILL_0_NOR2X1_201 gnd vdd FILL
XFILL_2_DFFPOSX1_785 gnd vdd FILL
XFILL_2_DFFPOSX1_796 gnd vdd FILL
XFILL_0_NOR2X1_223 gnd vdd FILL
XOAI21X1_208 BUFX4_164/Y BUFX4_64/Y BUFX2_1003/A gnd OAI21X1_209/C vdd OAI21X1
XOAI21X1_219 INVX2_155/Y BUFX4_289/Y OAI21X1_219/C gnd OAI21X1_219/Y vdd OAI21X1
XFILL_3_CLKBUF1_3 gnd vdd FILL
XDFFPOSX1_111 BUFX2_780/A CLKBUF1_14/Y OAI21X1_1785/Y gnd vdd DFFPOSX1
XDFFPOSX1_100 BUFX2_777/A CLKBUF1_47/Y OAI21X1_1774/Y gnd vdd DFFPOSX1
XAND2X2_19 AND2X2_19/A bundleStartMajId_i[51] gnd AND2X2_20/A vdd AND2X2
XDFFPOSX1_133 BUFX2_804/A CLKBUF1_39/Y OAI21X1_1807/Y gnd vdd DFFPOSX1
XDFFPOSX1_144 BUFX2_816/A CLKBUF1_7/Y OAI21X1_1818/Y gnd vdd DFFPOSX1
XDFFPOSX1_122 BUFX2_792/A CLKBUF1_67/Y OAI21X1_1796/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_331 gnd vdd FILL
XDFFPOSX1_155 BUFX2_828/A CLKBUF1_87/Y OAI21X1_1829/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_320 gnd vdd FILL
XFILL_38_15_1 gnd vdd FILL
XFILL_1_DFFPOSX1_342 gnd vdd FILL
XDFFPOSX1_188 BUFX2_858/A CLKBUF1_93/Y OAI21X1_32/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_353 gnd vdd FILL
XFILL_1_DFFPOSX1_375 gnd vdd FILL
XFILL_0_NOR3X1_9 gnd vdd FILL
XFILL_1_DFFPOSX1_364 gnd vdd FILL
XDFFPOSX1_166 BUFX2_853/A CLKBUF1_92/Y OAI21X1_10/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_590 gnd vdd FILL
XDFFPOSX1_177 BUFX2_846/A CLKBUF1_10/Y OAI21X1_21/Y gnd vdd DFFPOSX1
XNAND2X1_214 BUFX2_490/A BUFX4_213/Y gnd OAI21X1_457/C vdd NAND2X1
XDFFPOSX1_199 BUFX2_870/A CLKBUF1_73/Y OAI21X1_43/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_397 gnd vdd FILL
XNAND2X1_225 BUFX4_244/Y OAI21X1_465/Y gnd OAI21X1_466/A vdd NAND2X1
XFILL_1_DFFPOSX1_386 gnd vdd FILL
XNAND2X1_203 bundleStartMajId_i[31] INVX1_16/A gnd INVX1_15/A vdd NAND2X1
XFILL_4_DFFPOSX1_813 gnd vdd FILL
XNAND2X1_258 bundleStartMajId_i[4] INVX1_43/A gnd NOR2X1_99/B vdd NAND2X1
XNAND2X1_236 OAI21X1_474/Y OAI21X1_476/A gnd OAI21X1_475/A vdd NAND2X1
XFILL_4_DFFPOSX1_802 gnd vdd FILL
XNAND2X1_269 bundleStartMajId_i[60] bundleStartMajId_i[59] gnd NOR2X1_59/B vdd NAND2X1
XNAND2X1_247 BUFX2_507/A BUFX4_182/Y gnd OAI21X1_483/C vdd NAND2X1
XFILL_4_DFFPOSX1_835 gnd vdd FILL
XFILL_4_DFFPOSX1_824 gnd vdd FILL
XFILL_4_DFFPOSX1_846 gnd vdd FILL
XFILL_4_DFFPOSX1_879 gnd vdd FILL
XFILL_32_11_0 gnd vdd FILL
XFILL_4_DFFPOSX1_868 gnd vdd FILL
XFILL_4_DFFPOSX1_857 gnd vdd FILL
XFILL_0_OAI21X1_8 gnd vdd FILL
XFILL_26_7_1 gnd vdd FILL
XFILL_25_2_0 gnd vdd FILL
XFILL_1_7_1 gnd vdd FILL
XFILL_0_2_0 gnd vdd FILL
XFILL_4_CLKBUF1_91 gnd vdd FILL
XFILL_4_CLKBUF1_80 gnd vdd FILL
XFILL_0_BUFX2_62 gnd vdd FILL
XFILL_0_BUFX2_40 gnd vdd FILL
XFILL_1_NOR2X1_21 gnd vdd FILL
XFILL_0_BUFX2_51 gnd vdd FILL
XFILL_1_BUFX2_736 gnd vdd FILL
XFILL_1_BUFX2_725 gnd vdd FILL
XFILL_0_BUFX2_73 gnd vdd FILL
XFILL_0_BUFX2_84 gnd vdd FILL
XFILL_1_NOR2X1_54 gnd vdd FILL
XFILL_1_NOR2X1_43 gnd vdd FILL
XFILL_1_NOR2X1_32 gnd vdd FILL
XFILL_0_BUFX2_95 gnd vdd FILL
XFILL_1_BUFX2_747 gnd vdd FILL
XFILL_3_DFFPOSX1_403 gnd vdd FILL
XOAI21X1_731 INVX1_12/Y NOR2X1_108/B OAI21X1_731/C gnd OAI21X1_733/A vdd OAI21X1
XOAI21X1_742 BUFX4_130/Y BUFX4_67/Y BUFX2_607/A gnd OAI21X1_743/C vdd OAI21X1
XOAI21X1_720 XNOR2X1_44/Y BUFX4_300/Y OAI21X1_720/C gnd OAI21X1_720/Y vdd OAI21X1
XFILL_1_BUFX2_769 gnd vdd FILL
XFILL_3_DFFPOSX1_414 gnd vdd FILL
XOAI21X1_764 BUFX4_127/Y BUFX4_41/Y BUFX2_616/A gnd OAI21X1_765/C vdd OAI21X1
XOAI21X1_775 INVX4_31/Y INVX4_20/Y INVX2_28/Y gnd OAI21X1_776/C vdd OAI21X1
XOAI21X1_753 BUFX4_177/Y BUFX4_56/Y BUFX2_612/A gnd OAI21X1_754/C vdd OAI21X1
XFILL_3_DFFPOSX1_425 gnd vdd FILL
XFILL_3_DFFPOSX1_436 gnd vdd FILL
XFILL_3_DFFPOSX1_458 gnd vdd FILL
XFILL_3_DFFPOSX1_469 gnd vdd FILL
XOAI21X1_786 OAI21X1_786/A BUFX4_299/Y OAI21X1_786/C gnd OAI21X1_786/Y vdd OAI21X1
XOAI21X1_797 OR2X2_15/A NOR3X1_9/B INVX4_22/Y gnd OAI21X1_797/Y vdd OAI21X1
XFILL_3_DFFPOSX1_447 gnd vdd FILL
XFILL_37_10_0 gnd vdd FILL
XFILL_8_3_0 gnd vdd FILL
XFILL_9_8_1 gnd vdd FILL
XFILL_1_OAI21X1_270 gnd vdd FILL
XNAND2X1_770 BUFX2_828/A BUFX4_367/Y gnd NAND2X1_770/Y vdd NAND2X1
XFILL_1_OAI21X1_292 gnd vdd FILL
XFILL_1_OAI21X1_281 gnd vdd FILL
XFILL_2_XNOR2X1_21 gnd vdd FILL
XFILL_2_XNOR2X1_32 gnd vdd FILL
XFILL_2_XNOR2X1_10 gnd vdd FILL
XBUFX2_102 BUFX2_102/A gnd addr2_o[21] vdd BUFX2
XBUFX2_135 BUFX2_135/A gnd addr3_o[49] vdd BUFX2
XFILL_2_XNOR2X1_65 gnd vdd FILL
XBUFX2_124 BUFX2_124/A gnd addr2_o[1] vdd BUFX2
XFILL_2_XNOR2X1_43 gnd vdd FILL
XFILL_2_XNOR2X1_54 gnd vdd FILL
XBUFX2_113 BUFX2_113/A gnd addr2_o[11] vdd BUFX2
XFILL_2_XNOR2X1_76 gnd vdd FILL
XBUFX2_157 BUFX2_157/A gnd addr3_o[29] vdd BUFX2
XFILL_2_XNOR2X1_98 gnd vdd FILL
XBUFX2_168 BUFX2_168/A gnd addr3_o[19] vdd BUFX2
XFILL_17_7_1 gnd vdd FILL
XFILL_16_2_0 gnd vdd FILL
XBUFX2_146 BUFX2_146/A gnd addr3_o[39] vdd BUFX2
XFILL_2_XNOR2X1_87 gnd vdd FILL
XFILL_0_CLKBUF1_100 gnd vdd FILL
XFILL_1_NAND2X1_9 gnd vdd FILL
XBUFX2_179 BUFX2_179/A gnd addr3_o[9] vdd BUFX2
XFILL_5_DFFPOSX1_508 gnd vdd FILL
XFILL_5_DFFPOSX1_519 gnd vdd FILL
XBUFX2_1005 BUFX2_1005/A gnd tid4_o[22] vdd BUFX2
XBUFX2_1027 BUFX2_1027/A gnd tid4_o[2] vdd BUFX2
XBUFX2_1016 BUFX2_1016/A gnd tid4_o[12] vdd BUFX2
XFILL_3_DFFPOSX1_981 gnd vdd FILL
XFILL_3_DFFPOSX1_970 gnd vdd FILL
XFILL_3_DFFPOSX1_992 gnd vdd FILL
XCLKBUF1_39 BUFX4_85/Y gnd CLKBUF1_39/Y vdd CLKBUF1
XCLKBUF1_17 BUFX4_87/Y gnd CLKBUF1_17/Y vdd CLKBUF1
XFILL_4_DFFPOSX1_109 gnd vdd FILL
XCLKBUF1_28 BUFX4_88/Y gnd CLKBUF1_28/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_37 gnd vdd FILL
XFILL_1_DFFPOSX1_26 gnd vdd FILL
XFILL_1_DFFPOSX1_15 gnd vdd FILL
XFILL_1_DFFPOSX1_48 gnd vdd FILL
XBUFX4_60 BUFX4_60/A gnd BUFX4_60/Y vdd BUFX4
XFILL_1_DFFPOSX1_59 gnd vdd FILL
XBUFX4_71 BUFX4_71/A gnd BUFX4_71/Y vdd BUFX4
XBUFX4_82 BUFX4_82/A gnd BUFX4_82/Y vdd BUFX4
XBUFX4_93 BUFX4_9/A gnd BUFX4_93/Y vdd BUFX4
XFILL_0_OAI21X1_1804 gnd vdd FILL
XFILL_0_OAI21X1_1826 gnd vdd FILL
XFILL_0_OAI21X1_1815 gnd vdd FILL
XBUFX2_680 BUFX2_680/A gnd pid1_o[22] vdd BUFX2
XBUFX2_691 BUFX2_691/A gnd pid2_o[13] vdd BUFX2
XFILL_2_DFFPOSX1_582 gnd vdd FILL
XFILL_2_DFFPOSX1_593 gnd vdd FILL
XFILL_2_DFFPOSX1_560 gnd vdd FILL
XFILL_2_DFFPOSX1_571 gnd vdd FILL
XFILL_2_AOI21X1_43 gnd vdd FILL
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XFILL_1_DFFPOSX1_150 gnd vdd FILL
XFILL_1_DFFPOSX1_183 gnd vdd FILL
XFILL_1_DFFPOSX1_161 gnd vdd FILL
XFILL_1_DFFPOSX1_172 gnd vdd FILL
XXNOR2X1_3 NOR2X1_6/Y bundleStartMajId_i[50] gnd XNOR2X1_3/Y vdd XNOR2X1
XFILL_1_DFFPOSX1_194 gnd vdd FILL
XFILL_4_DFFPOSX1_621 gnd vdd FILL
XFILL_4_DFFPOSX1_610 gnd vdd FILL
XFILL_4_DFFPOSX1_654 gnd vdd FILL
XFILL_4_DFFPOSX1_632 gnd vdd FILL
XFILL_4_DFFPOSX1_643 gnd vdd FILL
XFILL_4_DFFPOSX1_698 gnd vdd FILL
XFILL_4_DFFPOSX1_687 gnd vdd FILL
XFILL_4_DFFPOSX1_665 gnd vdd FILL
XFILL_4_DFFPOSX1_676 gnd vdd FILL
XFILL_1_BUFX2_500 gnd vdd FILL
XFILL_1_INVX1_21 gnd vdd FILL
XFILL_1_BUFX2_533 gnd vdd FILL
XINVX1_3 bundleStartMajId_i[9] gnd INVX1_3/Y vdd INVX1
XFILL_1_BUFX2_544 gnd vdd FILL
XFILL_1_BUFX2_522 gnd vdd FILL
XFILL_3_DFFPOSX1_211 gnd vdd FILL
XFILL_3_DFFPOSX1_200 gnd vdd FILL
XFILL_0_BUFX4_118 gnd vdd FILL
XFILL_0_BUFX4_107 gnd vdd FILL
XFILL_23_16_0 gnd vdd FILL
XFILL_0_BUFX4_129 gnd vdd FILL
XFILL_1_BUFX2_588 gnd vdd FILL
XOAI21X1_550 OR2X2_5/A OR2X2_10/B OAI21X1_550/C gnd OAI21X1_552/A vdd OAI21X1
XFILL_1_BUFX2_577 gnd vdd FILL
XFILL_3_DFFPOSX1_255 gnd vdd FILL
XOAI21X1_583 BUFX4_97/Y BUFX4_334/Y BUFX2_546/A gnd OAI21X1_584/C vdd OAI21X1
XFILL_3_DFFPOSX1_244 gnd vdd FILL
XFILL_3_DFFPOSX1_222 gnd vdd FILL
XFILL_1_BUFX2_18 gnd vdd FILL
XFILL_3_DFFPOSX1_233 gnd vdd FILL
XOAI21X1_561 XNOR2X1_29/Y BUFX4_177/Y OAI21X1_561/C gnd OAI21X1_561/Y vdd OAI21X1
XOAI21X1_572 BUFX4_109/Y BUFX4_314/Y BUFX2_541/A gnd OAI21X1_574/C vdd OAI21X1
XFILL_3_DFFPOSX1_266 gnd vdd FILL
XFILL_3_DFFPOSX1_277 gnd vdd FILL
XFILL_1_BUFX2_29 gnd vdd FILL
XOAI21X1_594 OAI21X1_594/A BUFX4_122/Y OAI21X1_594/C gnd OAI21X1_594/Y vdd OAI21X1
XFILL_3_DFFPOSX1_288 gnd vdd FILL
XFILL_3_DFFPOSX1_299 gnd vdd FILL
XFILL_6_DFFPOSX1_715 gnd vdd FILL
XFILL_6_DFFPOSX1_726 gnd vdd FILL
XFILL_6_DFFPOSX1_759 gnd vdd FILL
XFILL_6_DFFPOSX1_737 gnd vdd FILL
XFILL_6_DFFPOSX1_748 gnd vdd FILL
XFILL_5_DFFPOSX1_7 gnd vdd FILL
XFILL_0_NAND2X1_307 gnd vdd FILL
XFILL_0_NAND2X1_329 gnd vdd FILL
XFILL_0_NAND2X1_318 gnd vdd FILL
XFILL_1_DFFPOSX1_1013 gnd vdd FILL
XFILL_32_5_1 gnd vdd FILL
XFILL_1_CLKBUF1_101 gnd vdd FILL
XFILL_1_DFFPOSX1_1002 gnd vdd FILL
XFILL_5_DFFPOSX1_316 gnd vdd FILL
XFILL_31_0_0 gnd vdd FILL
XFILL_1_DFFPOSX1_1024 gnd vdd FILL
XFILL_28_15_0 gnd vdd FILL
XFILL_5_DFFPOSX1_327 gnd vdd FILL
XFILL_5_DFFPOSX1_305 gnd vdd FILL
XFILL_5_DFFPOSX1_349 gnd vdd FILL
XFILL_5_DFFPOSX1_338 gnd vdd FILL
XOAI21X1_1824 BUFX4_359/Y INVX2_196/Y NAND2X1_765/Y gnd OAI21X1_1824/Y vdd OAI21X1
XOAI21X1_1813 BUFX4_375/Y INVX2_185/Y NAND2X1_754/Y gnd OAI21X1_1813/Y vdd OAI21X1
XOAI21X1_1802 BUFX4_343/Y INVX2_174/Y NAND2X1_743/Y gnd OAI21X1_1802/Y vdd OAI21X1
XFILL_0_OAI21X1_813 gnd vdd FILL
XFILL_0_OAI21X1_802 gnd vdd FILL
XFILL_0_OAI21X1_835 gnd vdd FILL
XFILL_0_OAI21X1_824 gnd vdd FILL
XFILL_0_OAI21X1_857 gnd vdd FILL
XFILL_0_OAI21X1_846 gnd vdd FILL
XFILL_0_OAI21X1_879 gnd vdd FILL
XFILL_0_OAI21X1_868 gnd vdd FILL
XFILL_2_DFFPOSX1_27 gnd vdd FILL
XFILL_2_DFFPOSX1_16 gnd vdd FILL
XFILL_2_DFFPOSX1_38 gnd vdd FILL
XFILL_2_DFFPOSX1_49 gnd vdd FILL
XFILL_3_16_0 gnd vdd FILL
XFILL_0_OAI21X1_1623 gnd vdd FILL
XFILL_0_OAI21X1_1601 gnd vdd FILL
XFILL_0_OAI21X1_1634 gnd vdd FILL
XFILL_0_OAI21X1_1612 gnd vdd FILL
XFILL_0_OAI21X1_1667 gnd vdd FILL
XFILL_0_OAI21X1_1656 gnd vdd FILL
XFILL_2_DFFPOSX1_390 gnd vdd FILL
XFILL_0_OAI21X1_1645 gnd vdd FILL
XFILL_0_OAI21X1_1678 gnd vdd FILL
XFILL_0_OAI21X1_1689 gnd vdd FILL
XFILL_23_5_1 gnd vdd FILL
XFILL_22_0_0 gnd vdd FILL
XFILL_5_DFFPOSX1_872 gnd vdd FILL
XFILL_0_BUFX4_9 gnd vdd FILL
XFILL_5_DFFPOSX1_850 gnd vdd FILL
XFILL_5_DFFPOSX1_861 gnd vdd FILL
XFILL_5_DFFPOSX1_883 gnd vdd FILL
XFILL_5_DFFPOSX1_894 gnd vdd FILL
XFILL_1_XNOR2X1_40 gnd vdd FILL
XFILL_4_DFFPOSX1_1006 gnd vdd FILL
XFILL_1_XNOR2X1_73 gnd vdd FILL
XFILL_1_XNOR2X1_62 gnd vdd FILL
XFILL_1_XNOR2X1_51 gnd vdd FILL
XFILL_4_DFFPOSX1_1017 gnd vdd FILL
XFILL_1_XNOR2X1_95 gnd vdd FILL
XFILL_4_DFFPOSX1_1028 gnd vdd FILL
XFILL_1_XNOR2X1_84 gnd vdd FILL
XFILL_8_15_0 gnd vdd FILL
XBUFX4_208 BUFX4_24/Y gnd BUFX4_208/Y vdd BUFX4
XBUFX4_219 BUFX4_23/Y gnd BUFX4_219/Y vdd BUFX4
XFILL_5_1_0 gnd vdd FILL
XFILL_6_6_1 gnd vdd FILL
XFILL_0_INVX2_107 gnd vdd FILL
XFILL_4_DFFPOSX1_462 gnd vdd FILL
XFILL_4_DFFPOSX1_451 gnd vdd FILL
XFILL_4_DFFPOSX1_473 gnd vdd FILL
XFILL_4_DFFPOSX1_440 gnd vdd FILL
XFILL_0_INVX2_118 gnd vdd FILL
XFILL_0_INVX2_129 gnd vdd FILL
XFILL_4_DFFPOSX1_484 gnd vdd FILL
XFILL_12_13_1 gnd vdd FILL
XFILL_4_DFFPOSX1_495 gnd vdd FILL
XFILL_0_INVX4_9 gnd vdd FILL
XFILL_14_5_1 gnd vdd FILL
XFILL_13_0_0 gnd vdd FILL
XFILL_1_BUFX2_330 gnd vdd FILL
XFILL_1_BUFX2_341 gnd vdd FILL
XFILL_1_BUFX2_385 gnd vdd FILL
XFILL_1_BUFX2_374 gnd vdd FILL
XOAI21X1_1109 INVX1_184/Y INVX1_185/A INVX2_59/Y gnd OAI21X1_1110/C vdd OAI21X1
XFILL_1_BUFX2_396 gnd vdd FILL
XFILL_1_OAI21X1_1329 gnd vdd FILL
XOAI21X1_380 BUFX4_372/Y NOR3X1_8/A OAI21X1_380/C gnd OAI21X1_380/Y vdd OAI21X1
XOAI21X1_391 BUFX4_346/Y INVX2_39/Y OAI21X1_391/C gnd OAI21X1_391/Y vdd OAI21X1
XFILL_1_OAI21X1_1307 gnd vdd FILL
XFILL_1_OAI21X1_1318 gnd vdd FILL
XAND2X2_3 AND2X2_3/A AND2X2_3/B gnd AND2X2_3/Y vdd AND2X2
XFILL_0_OAI21X1_109 gnd vdd FILL
XFILL_1_DFFPOSX1_919 gnd vdd FILL
XFILL_1_DFFPOSX1_908 gnd vdd FILL
XFILL_6_DFFPOSX1_501 gnd vdd FILL
XFILL_6_DFFPOSX1_512 gnd vdd FILL
XFILL_6_DFFPOSX1_523 gnd vdd FILL
XFILL_17_12_1 gnd vdd FILL
XFILL_30_14_1 gnd vdd FILL
XFILL_0_NAND2X1_115 gnd vdd FILL
XFILL_0_BUFX4_19 gnd vdd FILL
XFILL_0_NAND2X1_104 gnd vdd FILL
XFILL_0_INVX1_140 gnd vdd FILL
XFILL_0_NAND2X1_137 gnd vdd FILL
XFILL_0_NAND2X1_126 gnd vdd FILL
XFILL_1_NAND2X1_308 gnd vdd FILL
XFILL_0_NAND2X1_148 gnd vdd FILL
XFILL_0_NAND2X1_159 gnd vdd FILL
XFILL_0_INVX1_151 gnd vdd FILL
XFILL_1_AOI21X1_40 gnd vdd FILL
XFILL_1_AOI21X1_51 gnd vdd FILL
XFILL_0_DFFPOSX1_509 gnd vdd FILL
XFILL_0_INVX1_173 gnd vdd FILL
XFILL_0_INVX1_162 gnd vdd FILL
XFILL_0_INVX1_184 gnd vdd FILL
XFILL_1_AOI21X1_62 gnd vdd FILL
XFILL_0_INVX1_195 gnd vdd FILL
XFILL_5_DFFPOSX1_102 gnd vdd FILL
XFILL_5_DFFPOSX1_124 gnd vdd FILL
XFILL_2_CLKBUF1_102 gnd vdd FILL
XFILL_5_DFFPOSX1_135 gnd vdd FILL
XFILL_5_DFFPOSX1_113 gnd vdd FILL
XFILL_5_DFFPOSX1_157 gnd vdd FILL
XFILL_5_DFFPOSX1_168 gnd vdd FILL
XFILL_5_DFFPOSX1_146 gnd vdd FILL
XFILL_5_DFFPOSX1_179 gnd vdd FILL
XOAI21X1_1621 INVX2_124/Y BUFX4_207/Y NAND2X1_689/Y gnd DFFPOSX1_11/D vdd OAI21X1
XOAI21X1_1632 INVX2_135/Y BUFX4_183/Y NAND2X1_700/Y gnd DFFPOSX1_22/D vdd OAI21X1
XOAI21X1_1610 OAI21X1_7/A INVX2_114/Y NAND2X1_679/Y gnd DFFPOSX1_1/D vdd OAI21X1
XFILL_1_OAI21X1_1830 gnd vdd FILL
XOAI21X1_1665 BUFX4_140/Y INVX2_126/Y OAI21X1_1665/C gnd DFFPOSX1_45/D vdd OAI21X1
XOAI21X1_1654 BUFX4_2/A BUFX4_367/Y BUFX2_739/A gnd OAI21X1_1655/C vdd OAI21X1
XOAI21X1_1643 INVX2_114/Y BUFX4_188/Y NAND2X1_711/Y gnd DFFPOSX1_33/D vdd OAI21X1
XOAI21X1_1676 BUFX4_5/Y BUFX4_341/Y BUFX2_720/A gnd OAI21X1_1677/C vdd OAI21X1
XOAI21X1_1698 BUFX4_103/Y BUFX4_313/Y BUFX2_732/A gnd OAI21X1_1699/C vdd OAI21X1
XOAI21X1_1687 BUFX4_140/Y INVX2_137/Y OAI21X1_1687/C gnd DFFPOSX1_56/D vdd OAI21X1
XFILL_1_OAI21X1_803 gnd vdd FILL
XFILL_0_OAI21X1_632 gnd vdd FILL
XFILL_0_OAI21X1_610 gnd vdd FILL
XFILL_0_OAI21X1_621 gnd vdd FILL
XFILL_2_OAI22X1_1 gnd vdd FILL
XFILL_0_OAI21X1_654 gnd vdd FILL
XFILL_0_OAI21X1_643 gnd vdd FILL
XFILL_1_OAI21X1_836 gnd vdd FILL
XFILL_1_OAI21X1_825 gnd vdd FILL
XFILL_0_OAI21X1_665 gnd vdd FILL
XFILL_1_OAI21X1_814 gnd vdd FILL
XFILL_1_OAI21X1_858 gnd vdd FILL
XNAND3X1_19 bundleStartMajId_i[24] INVX4_19/Y NOR3X1_6/Y gnd NAND3X1_19/Y vdd NAND3X1
XFILL_1_OAI21X1_869 gnd vdd FILL
XFILL_1_OAI21X1_847 gnd vdd FILL
XFILL_0_OAI21X1_687 gnd vdd FILL
XFILL_0_OAI21X1_676 gnd vdd FILL
XFILL_0_OAI21X1_698 gnd vdd FILL
XFILL_35_13_1 gnd vdd FILL
XFILL_1_AND2X2_22 gnd vdd FILL
XFILL_1_AND2X2_11 gnd vdd FILL
XFILL_1_AND2X2_33 gnd vdd FILL
XFILL_3_DFFPOSX1_17 gnd vdd FILL
XNOR2X1_19 OR2X2_4/A NOR2X1_19/B gnd NOR2X1_19/Y vdd NOR2X1
XFILL_3_DFFPOSX1_39 gnd vdd FILL
XFILL_3_DFFPOSX1_28 gnd vdd FILL
XFILL_0_NAND2X1_660 gnd vdd FILL
XFILL_0_OAI21X1_1431 gnd vdd FILL
XFILL_0_OAI21X1_1420 gnd vdd FILL
XFILL_0_NAND2X1_671 gnd vdd FILL
XFILL_0_OAI21X1_1442 gnd vdd FILL
XFILL_0_NAND2X1_682 gnd vdd FILL
XFILL_0_OAI21X1_1475 gnd vdd FILL
XFILL_0_NAND2X1_693 gnd vdd FILL
XFILL_0_OAI21X1_1464 gnd vdd FILL
XFILL_0_OAI21X1_1453 gnd vdd FILL
XFILL_4_DFFPOSX1_4 gnd vdd FILL
XFILL_0_OAI21X1_1486 gnd vdd FILL
XFILL_0_OAI21X1_1497 gnd vdd FILL
XFILL_0_BUFX2_6 gnd vdd FILL
XFILL_5_DFFPOSX1_691 gnd vdd FILL
XFILL_5_DFFPOSX1_680 gnd vdd FILL
XFILL_0_BUFX2_408 gnd vdd FILL
XFILL_0_BUFX2_419 gnd vdd FILL
XFILL_2_OAI21X1_1514 gnd vdd FILL
XFILL_2_OAI21X1_1503 gnd vdd FILL
XFILL_4_DFFPOSX1_281 gnd vdd FILL
XFILL_0_NAND2X1_17 gnd vdd FILL
XFILL_0_NAND2X1_28 gnd vdd FILL
XFILL_4_DFFPOSX1_270 gnd vdd FILL
XFILL_4_DFFPOSX1_292 gnd vdd FILL
XFILL_0_NAND2X1_39 gnd vdd FILL
XNOR2X1_109 NOR2X1_30/A NOR3X1_9/A gnd NOR2X1_109/Y vdd NOR2X1
XFILL_0_INVX2_6 gnd vdd FILL
XFILL_1_BUFX2_171 gnd vdd FILL
XFILL_1_BUFX2_193 gnd vdd FILL
XFILL_1_OAI21X1_1104 gnd vdd FILL
XFILL_1_BUFX2_182 gnd vdd FILL
XFILL_1_OAI21X1_1126 gnd vdd FILL
XFILL_1_OAI21X1_1115 gnd vdd FILL
XFILL_0_BUFX2_920 gnd vdd FILL
XDFFPOSX1_529 BUFX2_561/A CLKBUF1_79/Y OAI21X1_617/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_942 gnd vdd FILL
XDFFPOSX1_507 BUFX2_537/A CLKBUF1_33/Y OAI21X1_563/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_705 gnd vdd FILL
XFILL_0_BUFX2_931 gnd vdd FILL
XDFFPOSX1_518 BUFX2_549/A CLKBUF1_48/Y OAI21X1_590/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1137 gnd vdd FILL
XFILL_0_BUFX2_975 gnd vdd FILL
XFILL_1_DFFPOSX1_749 gnd vdd FILL
XFILL_1_DFFPOSX1_716 gnd vdd FILL
XFILL_1_DFFPOSX1_727 gnd vdd FILL
XFILL_1_OAI21X1_1148 gnd vdd FILL
XFILL_0_BUFX2_964 gnd vdd FILL
XFILL_0_BUFX2_953 gnd vdd FILL
XFILL_1_OAI21X1_1159 gnd vdd FILL
XFILL_1_DFFPOSX1_738 gnd vdd FILL
XFILL_0_BUFX2_986 gnd vdd FILL
XFILL_0_BUFX2_997 gnd vdd FILL
XFILL_6_DFFPOSX1_375 gnd vdd FILL
XFILL_6_DFFPOSX1_386 gnd vdd FILL
XFILL_6_DFFPOSX1_364 gnd vdd FILL
XNAND2X1_52 BUFX2_880/A BUFX4_191/Y gnd OAI21X1_52/C vdd NAND2X1
XNAND2X1_41 BUFX2_868/A BUFX4_208/Y gnd OAI21X1_41/C vdd NAND2X1
XNAND2X1_30 BUFX2_856/A BUFX4_195/Y gnd OAI21X1_30/C vdd NAND2X1
XFILL_6_DFFPOSX1_397 gnd vdd FILL
XFILL_37_4_1 gnd vdd FILL
XNAND2X1_63 BUFX2_892/A BUFX4_180/Y gnd OAI21X1_63/C vdd NAND2X1
XNAND2X1_74 BUFX2_405/A BUFX4_365/Y gnd NAND2X1_74/Y vdd NAND2X1
XNAND2X1_85 BUFX2_398/A BUFX4_345/Y gnd NAND2X1_85/Y vdd NAND2X1
XFILL_0_XNOR2X1_81 gnd vdd FILL
XNAND2X1_96 BUFX2_410/A OAI21X1_2/A gnd NAND2X1_96/Y vdd NAND2X1
XFILL_0_XNOR2X1_70 gnd vdd FILL
XFILL_1_NAND2X1_105 gnd vdd FILL
XFILL_0_DFFPOSX1_306 gnd vdd FILL
XFILL_0_XNOR2X1_92 gnd vdd FILL
XFILL_1_NAND2X1_138 gnd vdd FILL
XFILL_0_DFFPOSX1_328 gnd vdd FILL
XFILL_0_DFFPOSX1_339 gnd vdd FILL
XFILL_0_DFFPOSX1_317 gnd vdd FILL
XFILL_1_NAND2X1_149 gnd vdd FILL
XFILL_20_3_1 gnd vdd FILL
XFILL_0_NOR3X1_13 gnd vdd FILL
XOAI21X1_1440 INVX2_97/Y INVX4_51/Y OAI21X1_1440/C gnd OAI21X1_1442/A vdd OAI21X1
XFILL_1_OAI21X1_1660 gnd vdd FILL
XOAI21X1_1473 NAND2X1_634/Y BUFX4_292/Y OAI21X1_1473/C gnd OAI21X1_1473/Y vdd OAI21X1
XOAI21X1_1462 XNOR2X1_98/Y BUFX4_292/Y OAI21X1_1462/C gnd OAI21X1_1462/Y vdd OAI21X1
XFILL_0_BUFX4_290 gnd vdd FILL
XOAI21X1_1484 XNOR2X1_100/Y BUFX4_294/Y OAI21X1_1484/C gnd OAI21X1_1484/Y vdd OAI21X1
XOAI21X1_1451 OAI21X1_1451/A INVX8_2/A OAI21X1_1451/C gnd OAI21X1_1451/Y vdd OAI21X1
XFILL_1_OAI21X1_1693 gnd vdd FILL
XFILL_1_OAI21X1_1682 gnd vdd FILL
XFILL_1_OAI21X1_611 gnd vdd FILL
XFILL_1_OAI21X1_1671 gnd vdd FILL
XOAI21X1_1495 BUFX4_157/Y BUFX4_80/Y BUFX2_224/A gnd OAI21X1_1496/C vdd OAI21X1
XFILL_1_OAI21X1_600 gnd vdd FILL
XFILL_0_OAI21X1_440 gnd vdd FILL
XFILL_1_OAI21X1_644 gnd vdd FILL
XFILL_1_NOR2X1_227 gnd vdd FILL
XFILL_2_OAI21X1_804 gnd vdd FILL
XFILL_0_OAI21X1_473 gnd vdd FILL
XFILL_1_OAI21X1_633 gnd vdd FILL
XFILL_0_OAI21X1_462 gnd vdd FILL
XFILL_1_OAI21X1_622 gnd vdd FILL
XFILL_0_OAI21X1_451 gnd vdd FILL
XFILL_1_OAI21X1_655 gnd vdd FILL
XFILL_0_OAI21X1_495 gnd vdd FILL
XFILL_3_NOR3X1_6 gnd vdd FILL
XFILL_1_OAI21X1_666 gnd vdd FILL
XFILL_0_OAI21X1_484 gnd vdd FILL
XFILL_2_OAI21X1_848 gnd vdd FILL
XFILL_1_OAI21X1_688 gnd vdd FILL
XFILL_1_OAI21X1_677 gnd vdd FILL
XFILL_1_INVX1_127 gnd vdd FILL
XFILL_1_OAI21X1_699 gnd vdd FILL
XFILL_28_4_1 gnd vdd FILL
XBUFX2_509 BUFX2_509/A gnd majID2_o[7] vdd BUFX2
XFILL_4_DFFPOSX1_18 gnd vdd FILL
XFILL_4_DFFPOSX1_29 gnd vdd FILL
XFILL_3_4_1 gnd vdd FILL
XFILL_0_OAI21X1_1250 gnd vdd FILL
XFILL_1_NAND2X1_683 gnd vdd FILL
XFILL_0_NAND2X1_490 gnd vdd FILL
XFILL_0_DFFPOSX1_840 gnd vdd FILL
XFILL_0_OAI21X1_1261 gnd vdd FILL
XFILL_0_DFFPOSX1_851 gnd vdd FILL
XFILL_1_NAND2X1_661 gnd vdd FILL
XFILL_0_OAI21X1_1283 gnd vdd FILL
XFILL_0_OAI21X1_1272 gnd vdd FILL
XFILL_0_DFFPOSX1_884 gnd vdd FILL
XFILL_0_OAI21X1_1294 gnd vdd FILL
XFILL_26_18_1 gnd vdd FILL
XFILL_0_DFFPOSX1_873 gnd vdd FILL
XFILL_0_DFFPOSX1_895 gnd vdd FILL
XFILL_0_DFFPOSX1_862 gnd vdd FILL
XDFFPOSX1_1014 BUFX2_651/A CLKBUF1_8/Y OAI21X1_1591/Y gnd vdd DFFPOSX1
XDFFPOSX1_1025 BUFX2_663/A CLKBUF1_64/Y OAI21X1_1602/Y gnd vdd DFFPOSX1
XDFFPOSX1_1003 BUFX2_392/A CLKBUF1_77/Y OAI21X1_1580/Y gnd vdd DFFPOSX1
XFILL_11_3_1 gnd vdd FILL
XFILL_0_BUFX2_205 gnd vdd FILL
XFILL_0_BUFX2_238 gnd vdd FILL
XFILL_0_BUFX2_216 gnd vdd FILL
XFILL_0_BUFX2_227 gnd vdd FILL
XFILL_0_BUFX2_249 gnd vdd FILL
XFILL_20_14_0 gnd vdd FILL
XOAI22X1_1 INVX1_26/Y OAI22X1_1/B OAI22X1_1/C bundleStartMajId_i[50] gnd OAI22X1_1/Y
+ vdd OAI22X1
XFILL_2_DFFPOSX1_901 gnd vdd FILL
XFILL_19_4_1 gnd vdd FILL
XFILL_2_OAI21X1_1344 gnd vdd FILL
XFILL_2_DFFPOSX1_923 gnd vdd FILL
XFILL_2_DFFPOSX1_912 gnd vdd FILL
XFILL_2_OAI21X1_1399 gnd vdd FILL
XFILL_2_DFFPOSX1_967 gnd vdd FILL
XFILL_2_DFFPOSX1_945 gnd vdd FILL
XFILL_2_DFFPOSX1_934 gnd vdd FILL
XFILL_2_DFFPOSX1_956 gnd vdd FILL
XFILL_2_DFFPOSX1_978 gnd vdd FILL
XFILL_2_DFFPOSX1_989 gnd vdd FILL
XFILL_6_DFFPOSX1_1030 gnd vdd FILL
XFILL_25_13_0 gnd vdd FILL
XFILL_3_XNOR2X1_14 gnd vdd FILL
XDFFPOSX1_304 BUFX2_973/A CLKBUF1_25/Y OAI21X1_225/Y gnd vdd DFFPOSX1
XFILL_3_XNOR2X1_36 gnd vdd FILL
XFILL_3_XNOR2X1_25 gnd vdd FILL
XFILL_3_XNOR2X1_47 gnd vdd FILL
XDFFPOSX1_337 BUFX2_1009/A CLKBUF1_102/Y OAI21X1_291/Y gnd vdd DFFPOSX1
XDFFPOSX1_326 BUFX2_997/A CLKBUF1_25/Y OAI21X1_269/Y gnd vdd DFFPOSX1
XDFFPOSX1_315 BUFX2_985/A CLKBUF1_86/Y OAI21X1_247/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_750 gnd vdd FILL
XFILL_1_DFFPOSX1_513 gnd vdd FILL
XFILL_1_DFFPOSX1_502 gnd vdd FILL
XFILL_1_DFFPOSX1_524 gnd vdd FILL
XFILL_0_BUFX2_783 gnd vdd FILL
XFILL_0_BUFX2_761 gnd vdd FILL
XFILL_0_BUFX2_794 gnd vdd FILL
XDFFPOSX1_348 BUFX2_1021/A CLKBUF1_43/Y OAI21X1_313/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_546 gnd vdd FILL
XFILL_1_DFFPOSX1_535 gnd vdd FILL
XFILL_0_NOR2X1_90 gnd vdd FILL
XDFFPOSX1_359 BUFX2_416/A CLKBUF1_4/Y OAI21X1_331/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_772 gnd vdd FILL
XFILL_1_DFFPOSX1_557 gnd vdd FILL
XNAND2X1_407 BUFX2_46/A BUFX4_347/Y gnd NAND2X1_407/Y vdd NAND2X1
XNAND2X1_418 BUFX2_9/A BUFX4_356/Y gnd NAND2X1_418/Y vdd NAND2X1
XFILL_1_DFFPOSX1_568 gnd vdd FILL
XFILL_1_DFFPOSX1_579 gnd vdd FILL
XFILL_6_DFFPOSX1_150 gnd vdd FILL
XNAND2X1_429 BUFX2_21/A BUFX4_317/Y gnd NAND2X1_429/Y vdd NAND2X1
XFILL_6_DFFPOSX1_161 gnd vdd FILL
XFILL_3_DFFPOSX1_1 gnd vdd FILL
XFILL_6_DFFPOSX1_172 gnd vdd FILL
XFILL_6_18_1 gnd vdd FILL
XBUFX4_380 BUFX4_380/A gnd BUFX4_380/Y vdd BUFX4
XFILL_0_DFFPOSX1_114 gnd vdd FILL
XFILL_0_DFFPOSX1_103 gnd vdd FILL
XFILL_0_14_0 gnd vdd FILL
XFILL_0_DFFPOSX1_125 gnd vdd FILL
XFILL_0_DFFPOSX1_147 gnd vdd FILL
XFILL_0_DFFPOSX1_136 gnd vdd FILL
XFILL_1_BUFX2_929 gnd vdd FILL
XFILL_1_BUFX2_918 gnd vdd FILL
XFILL_1_BUFX2_907 gnd vdd FILL
XFILL_0_DFFPOSX1_158 gnd vdd FILL
XFILL_0_DFFPOSX1_169 gnd vdd FILL
XFILL_0_NAND2X1_1 gnd vdd FILL
XOAI21X1_924 BUFX4_2/A BUFX4_352/Y BUFX2_355/A gnd OAI21X1_925/C vdd OAI21X1
XOAI21X1_902 INVX1_103/Y BUFX4_232/Y OAI21X1_902/C gnd OAI21X1_902/Y vdd OAI21X1
XOAI21X1_913 BUFX4_153/Y INVX1_111/Y OAI21X1_913/C gnd OAI21X1_913/Y vdd OAI21X1
XOAI21X1_957 BUFX4_143/Y INVX1_133/Y OAI21X1_957/C gnd OAI21X1_957/Y vdd OAI21X1
XFILL_3_DFFPOSX1_607 gnd vdd FILL
XOAI21X1_935 BUFX4_153/Y INVX1_122/Y OAI21X1_935/C gnd OAI21X1_935/Y vdd OAI21X1
XFILL_3_DFFPOSX1_629 gnd vdd FILL
XFILL_3_DFFPOSX1_618 gnd vdd FILL
XOAI21X1_946 BUFX4_96/Y OAI21X1_7/A BUFX2_336/A gnd OAI21X1_947/C vdd OAI21X1
XOAI21X1_979 BUFX4_291/Y INVX1_144/Y OAI21X1_979/C gnd OAI21X1_979/Y vdd OAI21X1
XOAI21X1_968 BUFX4_111/Y BUFX4_332/Y BUFX2_349/A gnd OAI21X1_969/C vdd OAI21X1
XOAI21X1_1292 AOI21X1_48/Y OR2X2_20/Y OAI21X1_1292/C gnd OAI21X1_1292/Y vdd OAI21X1
XOAI21X1_1281 BUFX4_95/A BUFX4_311/Y BUFX2_148/A gnd OAI21X1_1282/C vdd OAI21X1
XOAI21X1_1270 BUFX4_6/A BUFX4_324/Y BUFX2_143/A gnd OAI21X1_1271/C vdd OAI21X1
XDFFPOSX1_860 BUFX2_113/A CLKBUF1_76/Y OAI21X1_1185/Y gnd vdd DFFPOSX1
XDFFPOSX1_882 BUFX2_131/A CLKBUF1_72/Y OAI21X1_1235/Y gnd vdd DFFPOSX1
XDFFPOSX1_871 BUFX2_125/A CLKBUF1_97/Y OAI21X1_1207/Y gnd vdd DFFPOSX1
XDFFPOSX1_893 BUFX2_143/A CLKBUF1_77/Y OAI21X1_1271/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1490 gnd vdd FILL
XINVX2_10 bundleStartMajId_i[60] gnd INVX2_10/Y vdd INVX2
XINVX2_21 bundleStartMajId_i[41] gnd INVX2_21/Y vdd INVX2
XINVX2_54 bundleAddress_i[63] gnd INVX2_54/Y vdd INVX2
XFILL_0_OAI21X1_270 gnd vdd FILL
XFILL_1_OAI21X1_463 gnd vdd FILL
XINVX2_32 bundleStartMajId_i[16] gnd INVX2_32/Y vdd INVX2
XFILL_2_OAI21X1_623 gnd vdd FILL
XINVX2_43 INVX2_43/A gnd INVX2_43/Y vdd INVX2
XFILL_0_OAI21X1_281 gnd vdd FILL
XFILL_1_OAI21X1_452 gnd vdd FILL
XFILL_1_OAI21X1_430 gnd vdd FILL
XFILL_1_OAI21X1_441 gnd vdd FILL
XINVX2_65 bundleAddress_i[50] gnd INVX2_65/Y vdd INVX2
XFILL_1_OAI21X1_496 gnd vdd FILL
XFILL_1_OAI21X1_474 gnd vdd FILL
XFILL_0_OAI21X1_292 gnd vdd FILL
XINVX2_87 bundleAddress_i[9] gnd INVX2_87/Y vdd INVX2
XFILL_1_OAI21X1_485 gnd vdd FILL
XINVX2_76 bundleAddress_i[28] gnd INVX2_76/Y vdd INVX2
XINVX2_98 INVX2_98/A gnd INVX2_98/Y vdd INVX2
XFILL_5_13_0 gnd vdd FILL
XFILL_2_DFFPOSX1_208 gnd vdd FILL
XBUFX2_306 BUFX2_306/A gnd instr2_o[11] vdd BUFX2
XFILL_0_AOI21X1_6 gnd vdd FILL
XFILL_2_DFFPOSX1_219 gnd vdd FILL
XBUFX2_317 BUFX2_317/A gnd instr2_o[1] vdd BUFX2
XFILL_5_DFFPOSX1_19 gnd vdd FILL
XBUFX2_339 BUFX2_339/A gnd instr3_o[10] vdd BUFX2
XBUFX2_328 BUFX2_328/A gnd instr3_o[20] vdd BUFX2
XFILL_1_INVX4_21 gnd vdd FILL
XFILL_1_INVX4_10 gnd vdd FILL
XFILL_1_INVX4_43 gnd vdd FILL
XFILL_1_BUFX4_211 gnd vdd FILL
XFILL_1_BUFX4_200 gnd vdd FILL
XOAI21X1_17 INVX2_155/Y BUFX4_224/Y OAI21X1_17/C gnd OAI21X1_17/Y vdd OAI21X1
XFILL_1_BUFX4_222 gnd vdd FILL
XFILL_1_NAND2X1_491 gnd vdd FILL
XFILL_0_DFFPOSX1_670 gnd vdd FILL
XFILL_1_NAND2X1_480 gnd vdd FILL
XFILL_0_OAI21X1_1080 gnd vdd FILL
XOAI21X1_39 INVX2_177/Y BUFX4_230/Y OAI21X1_39/C gnd OAI21X1_39/Y vdd OAI21X1
XFILL_1_BUFX4_255 gnd vdd FILL
XFILL_1_BUFX4_244 gnd vdd FILL
XFILL_0_OAI21X1_1091 gnd vdd FILL
XOAI21X1_28 INVX2_166/Y BUFX4_233/Y OAI21X1_28/C gnd OAI21X1_28/Y vdd OAI21X1
XFILL_1_BUFX4_233 gnd vdd FILL
XFILL_0_DFFPOSX1_692 gnd vdd FILL
XFILL_0_DFFPOSX1_681 gnd vdd FILL
XFILL_1_BUFX4_266 gnd vdd FILL
XFILL_1_BUFX4_288 gnd vdd FILL
XFILL_1_BUFX4_277 gnd vdd FILL
XFILL_1_BUFX4_299 gnd vdd FILL
XFILL_0_DFFPOSX1_26 gnd vdd FILL
XFILL_0_DFFPOSX1_15 gnd vdd FILL
XFILL_0_DFFPOSX1_59 gnd vdd FILL
XFILL_0_DFFPOSX1_37 gnd vdd FILL
XFILL_0_DFFPOSX1_48 gnd vdd FILL
XFILL_2_XNOR2X1_4 gnd vdd FILL
XFILL_14_10_1 gnd vdd FILL
XBUFX2_840 BUFX2_840/A gnd tid1_o[54] vdd BUFX2
XFILL_2_DFFPOSX1_720 gnd vdd FILL
XFILL_2_DFFPOSX1_731 gnd vdd FILL
XFILL_2_OAI21X1_1163 gnd vdd FILL
XFILL_2_DFFPOSX1_742 gnd vdd FILL
XFILL_34_2_1 gnd vdd FILL
XBUFX2_873 BUFX2_873/A gnd tid2_o[25] vdd BUFX2
XFILL_2_DFFPOSX1_753 gnd vdd FILL
XFILL_2_DFFPOSX1_775 gnd vdd FILL
XBUFX2_851 BUFX2_851/A gnd tid2_o[45] vdd BUFX2
XBUFX2_862 BUFX2_862/A gnd tid2_o[35] vdd BUFX2
XFILL_2_DFFPOSX1_764 gnd vdd FILL
XBUFX2_884 BUFX2_884/A gnd tid2_o[15] vdd BUFX2
XFILL_0_NOR2X1_213 gnd vdd FILL
XFILL_2_DFFPOSX1_786 gnd vdd FILL
XFILL_0_NOR2X1_202 gnd vdd FILL
XFILL_2_DFFPOSX1_797 gnd vdd FILL
XBUFX2_895 BUFX2_895/A gnd tid2_o[5] vdd BUFX2
XFILL_0_NOR2X1_224 gnd vdd FILL
XOAI21X1_209 INVX2_150/Y BUFX4_291/Y OAI21X1_209/C gnd OAI21X1_209/Y vdd OAI21X1
XFILL_12_1 gnd vdd FILL
XFILL_3_CLKBUF1_4 gnd vdd FILL
XDFFPOSX1_112 BUFX2_781/A CLKBUF1_17/Y OAI21X1_1786/Y gnd vdd DFFPOSX1
XDFFPOSX1_101 BUFX2_778/A CLKBUF1_71/Y OAI21X1_1775/Y gnd vdd DFFPOSX1
XDFFPOSX1_134 BUFX2_805/A CLKBUF1_11/Y OAI21X1_1808/Y gnd vdd DFFPOSX1
XDFFPOSX1_145 BUFX2_817/A CLKBUF1_11/Y OAI21X1_1819/Y gnd vdd DFFPOSX1
XDFFPOSX1_123 BUFX2_793/A CLKBUF1_67/Y OAI21X1_1797/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_321 gnd vdd FILL
XFILL_1_DFFPOSX1_310 gnd vdd FILL
XFILL_1_DFFPOSX1_332 gnd vdd FILL
XDFFPOSX1_178 BUFX2_847/A CLKBUF1_57/Y OAI21X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_156 BUFX2_829/A CLKBUF1_93/Y OAI21X1_1830/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_580 gnd vdd FILL
XDFFPOSX1_189 BUFX2_859/A CLKBUF1_3/Y OAI21X1_33/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_343 gnd vdd FILL
XFILL_1_DFFPOSX1_354 gnd vdd FILL
XFILL_0_BUFX2_591 gnd vdd FILL
XFILL_1_DFFPOSX1_365 gnd vdd FILL
XDFFPOSX1_167 BUFX2_864/A CLKBUF1_41/Y OAI21X1_11/Y gnd vdd DFFPOSX1
XNAND2X1_215 bundleStartMajId_i[25] NOR2X1_33/Y gnd XNOR2X1_18/A vdd NAND2X1
XFILL_1_DFFPOSX1_398 gnd vdd FILL
XFILL_1_DFFPOSX1_376 gnd vdd FILL
XNAND2X1_204 BUFX2_483/A BUFX4_194/Y gnd OAI21X1_449/C vdd NAND2X1
XNAND2X1_226 BUFX2_496/A BUFX4_182/Y gnd OAI21X1_466/C vdd NAND2X1
XFILL_1_DFFPOSX1_387 gnd vdd FILL
XNAND2X1_237 BUFX2_501/A BUFX4_200/Y gnd OAI21X1_475/C vdd NAND2X1
XFILL_4_DFFPOSX1_803 gnd vdd FILL
XNAND2X1_259 BUFX2_514/A BUFX4_221/Y gnd OAI21X1_494/C vdd NAND2X1
XNAND2X1_248 BUFX2_508/A BUFX4_182/Y gnd OAI21X1_485/C vdd NAND2X1
XFILL_4_DFFPOSX1_814 gnd vdd FILL
XFILL_4_DFFPOSX1_825 gnd vdd FILL
XFILL_4_DFFPOSX1_836 gnd vdd FILL
XFILL_16_18_0 gnd vdd FILL
XFILL_4_DFFPOSX1_847 gnd vdd FILL
XFILL_32_11_1 gnd vdd FILL
XFILL_4_DFFPOSX1_869 gnd vdd FILL
XFILL_4_DFFPOSX1_858 gnd vdd FILL
XFILL_4_CLKBUF1_70 gnd vdd FILL
XFILL_25_2_1 gnd vdd FILL
XFILL_0_OAI21X1_9 gnd vdd FILL
XFILL_0_BUFX2_30 gnd vdd FILL
XFILL_0_2_1 gnd vdd FILL
XFILL_4_CLKBUF1_81 gnd vdd FILL
XFILL_4_CLKBUF1_92 gnd vdd FILL
XFILL_0_BUFX2_63 gnd vdd FILL
XFILL_0_BUFX2_41 gnd vdd FILL
XFILL_0_BUFX2_52 gnd vdd FILL
XFILL_1_BUFX2_704 gnd vdd FILL
XFILL_0_BUFX2_85 gnd vdd FILL
XFILL_1_BUFX2_726 gnd vdd FILL
XFILL_1_BUFX2_715 gnd vdd FILL
XFILL_0_BUFX2_74 gnd vdd FILL
XFILL_1_NOR2X1_55 gnd vdd FILL
XFILL_1_NOR2X1_22 gnd vdd FILL
XFILL_0_BUFX2_96 gnd vdd FILL
XFILL_1_BUFX2_759 gnd vdd FILL
XOAI21X1_710 BUFX4_175/Y BUFX4_54/Y BUFX2_595/A gnd OAI21X1_711/C vdd OAI21X1
XOAI21X1_732 BUFX4_133/Y BUFX4_79/A BUFX2_603/A gnd OAI21X1_733/C vdd OAI21X1
XOAI21X1_721 INVX1_37/A INVX4_8/Y INVX2_21/Y gnd OAI21X1_722/C vdd OAI21X1
XFILL_1_NOR2X1_88 gnd vdd FILL
XFILL_3_DFFPOSX1_404 gnd vdd FILL
XFILL_1_NOR2X1_66 gnd vdd FILL
XFILL_3_DFFPOSX1_415 gnd vdd FILL
XOAI21X1_765 XNOR2X1_50/Y BUFX4_291/Y OAI21X1_765/C gnd OAI21X1_765/Y vdd OAI21X1
XOAI21X1_776 NOR3X1_3/A NOR2X1_114/B OAI21X1_776/C gnd OAI21X1_778/A vdd OAI21X1
XOAI21X1_743 XNOR2X1_47/Y BUFX4_295/Y OAI21X1_743/C gnd OAI21X1_743/Y vdd OAI21X1
XOAI21X1_754 OAI21X1_754/A BUFX4_300/Y OAI21X1_754/C gnd OAI21X1_754/Y vdd OAI21X1
XFILL_3_DFFPOSX1_426 gnd vdd FILL
XFILL_3_DFFPOSX1_437 gnd vdd FILL
XOAI21X1_798 BUFX4_161/Y BUFX4_62/Y BUFX2_628/A gnd OAI21X1_799/C vdd OAI21X1
XFILL_3_DFFPOSX1_459 gnd vdd FILL
XOAI21X1_787 INVX4_31/Y INVX2_49/Y INVX2_30/Y gnd OAI21X1_787/Y vdd OAI21X1
XFILL_3_DFFPOSX1_448 gnd vdd FILL
XFILL_6_DFFPOSX1_919 gnd vdd FILL
XFILL_6_DFFPOSX1_908 gnd vdd FILL
XFILL_37_10_1 gnd vdd FILL
XDFFPOSX1_690 BUFX2_327/A CLKBUF1_39/Y OAI21X1_929/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_260 gnd vdd FILL
XFILL_1_OAI21X1_271 gnd vdd FILL
XFILL_2_OAI21X1_420 gnd vdd FILL
XFILL_8_3_1 gnd vdd FILL
XNAND2X1_760 BUFX2_817/A BUFX4_316/Y gnd NAND2X1_760/Y vdd NAND2X1
XNAND2X1_771 BUFX2_829/A BUFX4_361/Y gnd NAND2X1_771/Y vdd NAND2X1
XFILL_1_OAI21X1_282 gnd vdd FILL
XFILL_1_OAI21X1_293 gnd vdd FILL
XFILL_2_XNOR2X1_22 gnd vdd FILL
XFILL_2_XNOR2X1_11 gnd vdd FILL
XBUFX2_103 BUFX2_103/A gnd addr2_o[20] vdd BUFX2
XFILL_2_XNOR2X1_55 gnd vdd FILL
XBUFX2_125 BUFX2_125/A gnd addr2_o[0] vdd BUFX2
XFILL_2_XNOR2X1_33 gnd vdd FILL
XFILL_2_XNOR2X1_44 gnd vdd FILL
XBUFX2_114 BUFX2_114/A gnd addr2_o[10] vdd BUFX2
XBUFX2_136 BUFX2_136/A gnd addr3_o[48] vdd BUFX2
XFILL_2_XNOR2X1_77 gnd vdd FILL
XFILL_2_XNOR2X1_99 gnd vdd FILL
XFILL_2_XNOR2X1_66 gnd vdd FILL
XFILL_2_XNOR2X1_88 gnd vdd FILL
XFILL_16_2_1 gnd vdd FILL
XBUFX2_169 BUFX2_169/A gnd addr3_o[18] vdd BUFX2
XBUFX2_158 BUFX2_158/A gnd addr3_o[28] vdd BUFX2
XBUFX2_147 BUFX2_147/A gnd addr3_o[38] vdd BUFX2
XFILL_0_CLKBUF1_101 gnd vdd FILL
XFILL_5_DFFPOSX1_509 gnd vdd FILL
XBUFX2_1017 BUFX2_1017/A gnd tid4_o[11] vdd BUFX2
XBUFX2_1006 BUFX2_1006/A gnd tid4_o[21] vdd BUFX2
XBUFX2_1028 BUFX2_1028/A gnd tid4_o[1] vdd BUFX2
XFILL_3_DFFPOSX1_982 gnd vdd FILL
XFILL_3_DFFPOSX1_960 gnd vdd FILL
XFILL_3_DFFPOSX1_993 gnd vdd FILL
XFILL_3_DFFPOSX1_971 gnd vdd FILL
XCLKBUF1_29 BUFX4_84/Y gnd CLKBUF1_29/Y vdd CLKBUF1
XCLKBUF1_18 BUFX4_91/Y gnd CLKBUF1_18/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_27 gnd vdd FILL
XFILL_1_DFFPOSX1_38 gnd vdd FILL
XFILL_1_DFFPOSX1_16 gnd vdd FILL
XBUFX4_50 BUFX4_55/A gnd BUFX4_50/Y vdd BUFX4
XBUFX4_61 BUFX4_82/A gnd BUFX4_61/Y vdd BUFX4
XFILL_1_DFFPOSX1_49 gnd vdd FILL
XBUFX4_94 BUFX4_94/A gnd BUFX4_94/Y vdd BUFX4
XBUFX4_83 clock_i gnd BUFX4_83/Y vdd BUFX4
XFILL_2_BUFX4_209 gnd vdd FILL
XBUFX4_72 BUFX4_72/A gnd BUFX4_72/Y vdd BUFX4
XFILL_0_OAI21X1_1805 gnd vdd FILL
XFILL_2_DFFPOSX1_550 gnd vdd FILL
XFILL_0_OAI21X1_1816 gnd vdd FILL
XBUFX2_670 BUFX2_670/A gnd pid1_o[3] vdd BUFX2
XFILL_0_OAI21X1_1827 gnd vdd FILL
XBUFX2_681 BUFX2_681/A gnd pid2_o[31] vdd BUFX2
XFILL_2_DFFPOSX1_583 gnd vdd FILL
XFILL_2_DFFPOSX1_572 gnd vdd FILL
XFILL_2_DFFPOSX1_561 gnd vdd FILL
XFILL_2_DFFPOSX1_594 gnd vdd FILL
XBUFX2_692 BUFX2_692/A gnd pid2_o[12] vdd BUFX2
XOR2X2_20 OR2X2_20/A OR2X2_20/B gnd OR2X2_20/Y vdd OR2X2
XOR2X2_2 OR2X2_5/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XFILL_1_DFFPOSX1_140 gnd vdd FILL
XFILL_1_DFFPOSX1_173 gnd vdd FILL
XFILL_1_DFFPOSX1_151 gnd vdd FILL
XFILL_1_DFFPOSX1_162 gnd vdd FILL
XXNOR2X1_4 NOR2X1_9/B NOR2X1_9/A gnd XNOR2X1_4/Y vdd XNOR2X1
XFILL_1_DFFPOSX1_195 gnd vdd FILL
XFILL_1_DFFPOSX1_184 gnd vdd FILL
XFILL_4_DFFPOSX1_600 gnd vdd FILL
XFILL_4_DFFPOSX1_611 gnd vdd FILL
XFILL_4_DFFPOSX1_622 gnd vdd FILL
XFILL_4_DFFPOSX1_655 gnd vdd FILL
XFILL_4_DFFPOSX1_633 gnd vdd FILL
XFILL_4_DFFPOSX1_644 gnd vdd FILL
XFILL_4_DFFPOSX1_688 gnd vdd FILL
XFILL_4_DFFPOSX1_677 gnd vdd FILL
XFILL_4_DFFPOSX1_666 gnd vdd FILL
XFILL_4_DFFPOSX1_699 gnd vdd FILL
XFILL_1_BUFX2_512 gnd vdd FILL
XINVX1_4 bundleStartMajId_i[4] gnd INVX1_4/Y vdd INVX1
XFILL_1_BUFX2_523 gnd vdd FILL
XFILL_1_BUFX2_578 gnd vdd FILL
XFILL_3_DFFPOSX1_212 gnd vdd FILL
XFILL_1_BUFX2_567 gnd vdd FILL
XFILL_3_DFFPOSX1_201 gnd vdd FILL
XFILL_0_BUFX4_108 gnd vdd FILL
XFILL_23_16_1 gnd vdd FILL
XFILL_0_BUFX4_119 gnd vdd FILL
XOAI21X1_540 BUFX4_98/Y BUFX4_365/Y BUFX2_527/A gnd OAI21X1_541/C vdd OAI21X1
XFILL_1_INVX1_77 gnd vdd FILL
XFILL_10_9_0 gnd vdd FILL
XFILL_1_BUFX2_556 gnd vdd FILL
XFILL_3_DFFPOSX1_245 gnd vdd FILL
XFILL_3_DFFPOSX1_234 gnd vdd FILL
XOAI21X1_584 OAI21X1_584/A BUFX4_149/Y OAI21X1_584/C gnd OAI21X1_584/Y vdd OAI21X1
XOAI21X1_551 BUFX4_4/Y BUFX4_314/Y BUFX2_531/A gnd OAI21X1_552/C vdd OAI21X1
XOAI21X1_573 NOR2X1_70/B OAI21X1_575/B INVX8_6/A gnd OAI21X1_574/B vdd OAI21X1
XFILL_3_DFFPOSX1_223 gnd vdd FILL
XOAI21X1_562 BUFX4_10/A BUFX4_383/Y BUFX2_537/A gnd OAI21X1_563/C vdd OAI21X1
XFILL_3_DFFPOSX1_278 gnd vdd FILL
XFILL_3_DFFPOSX1_267 gnd vdd FILL
XOAI21X1_595 BUFX4_3/Y BUFX4_346/Y BUFX2_551/A gnd OAI21X1_596/C vdd OAI21X1
XFILL_1_BUFX2_19 gnd vdd FILL
XFILL_3_DFFPOSX1_256 gnd vdd FILL
XFILL_3_DFFPOSX1_289 gnd vdd FILL
XFILL_6_DFFPOSX1_705 gnd vdd FILL
XFILL_5_DFFPOSX1_8 gnd vdd FILL
XFILL_2_OAI21X1_272 gnd vdd FILL
XNAND2X1_590 INVX2_56/Y INVX2_57/Y gnd NAND2X1_591/B vdd NAND2X1
XFILL_0_NAND2X1_308 gnd vdd FILL
XFILL_0_NAND2X1_319 gnd vdd FILL
XFILL_1_CLKBUF1_102 gnd vdd FILL
XFILL_1_DFFPOSX1_1003 gnd vdd FILL
XFILL_5_DFFPOSX1_306 gnd vdd FILL
XFILL_1_DFFPOSX1_1014 gnd vdd FILL
XFILL_31_0_1 gnd vdd FILL
XFILL_1_DFFPOSX1_1025 gnd vdd FILL
XFILL_28_15_1 gnd vdd FILL
XFILL_5_DFFPOSX1_317 gnd vdd FILL
XFILL_5_DFFPOSX1_328 gnd vdd FILL
XFILL_5_DFFPOSX1_339 gnd vdd FILL
XFILL_22_11_0 gnd vdd FILL
XOAI21X1_1803 BUFX4_384/Y INVX2_175/Y NAND2X1_744/Y gnd OAI21X1_1803/Y vdd OAI21X1
XOAI21X1_1814 BUFX4_314/Y INVX2_186/Y NAND2X1_755/Y gnd OAI21X1_1814/Y vdd OAI21X1
XOAI21X1_1825 BUFX4_348/Y INVX2_197/Y NAND2X1_766/Y gnd OAI21X1_1825/Y vdd OAI21X1
XFILL_3_DFFPOSX1_790 gnd vdd FILL
XFILL_0_OAI21X1_803 gnd vdd FILL
XFILL_0_OAI21X1_814 gnd vdd FILL
XFILL_0_OAI21X1_836 gnd vdd FILL
XFILL_0_OAI21X1_825 gnd vdd FILL
XFILL_0_OAI21X1_847 gnd vdd FILL
XFILL_0_OAI21X1_858 gnd vdd FILL
XFILL_0_OAI21X1_869 gnd vdd FILL
XFILL_2_DFFPOSX1_17 gnd vdd FILL
XFILL_2_DFFPOSX1_28 gnd vdd FILL
XFILL_2_DFFPOSX1_39 gnd vdd FILL
XFILL_3_16_1 gnd vdd FILL
XFILL_0_OAI21X1_1613 gnd vdd FILL
XFILL_0_OAI21X1_1602 gnd vdd FILL
XFILL_0_OAI21X1_1624 gnd vdd FILL
XFILL_0_OAI21X1_1646 gnd vdd FILL
XFILL_0_OAI21X1_1668 gnd vdd FILL
XFILL_0_OAI21X1_1635 gnd vdd FILL
XFILL_2_DFFPOSX1_391 gnd vdd FILL
XFILL_2_DFFPOSX1_380 gnd vdd FILL
XFILL_0_OAI21X1_1657 gnd vdd FILL
XFILL_0_OAI21X1_1679 gnd vdd FILL
XFILL_22_0_1 gnd vdd FILL
XFILL_5_DFFPOSX1_840 gnd vdd FILL
XFILL_27_10_0 gnd vdd FILL
XFILL_5_DFFPOSX1_851 gnd vdd FILL
XFILL_5_DFFPOSX1_873 gnd vdd FILL
XFILL_5_DFFPOSX1_862 gnd vdd FILL
XFILL_5_DFFPOSX1_884 gnd vdd FILL
XFILL_5_DFFPOSX1_895 gnd vdd FILL
XFILL_1_XNOR2X1_30 gnd vdd FILL
XFILL_1_XNOR2X1_63 gnd vdd FILL
XFILL_1_XNOR2X1_52 gnd vdd FILL
XFILL_1_XNOR2X1_41 gnd vdd FILL
XFILL_1_XNOR2X1_74 gnd vdd FILL
XFILL_4_DFFPOSX1_1018 gnd vdd FILL
XFILL_4_DFFPOSX1_1007 gnd vdd FILL
XFILL_1_XNOR2X1_85 gnd vdd FILL
XFILL_1_XNOR2X1_96 gnd vdd FILL
XFILL_4_DFFPOSX1_1029 gnd vdd FILL
XFILL_8_15_1 gnd vdd FILL
XBUFX4_209 BUFX4_22/Y gnd BUFX4_209/Y vdd BUFX4
XFILL_4_DFFPOSX1_430 gnd vdd FILL
XFILL_2_OAI21X1_1729 gnd vdd FILL
XFILL_0_INVX2_108 gnd vdd FILL
XFILL_4_DFFPOSX1_463 gnd vdd FILL
XFILL_5_1_1 gnd vdd FILL
XFILL_4_DFFPOSX1_452 gnd vdd FILL
XFILL_4_DFFPOSX1_441 gnd vdd FILL
XFILL_0_INVX2_119 gnd vdd FILL
XFILL_4_DFFPOSX1_485 gnd vdd FILL
XFILL_2_11_0 gnd vdd FILL
XFILL_4_DFFPOSX1_496 gnd vdd FILL
XFILL_4_DFFPOSX1_474 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XFILL_1_BUFX2_320 gnd vdd FILL
XFILL_1_BUFX2_331 gnd vdd FILL
XFILL_1_BUFX2_353 gnd vdd FILL
XFILL_1_BUFX2_375 gnd vdd FILL
XFILL_1_BUFX2_364 gnd vdd FILL
XOAI21X1_370 BUFX4_325/Y INVX2_28/Y OAI21X1_370/C gnd OAI21X1_370/Y vdd OAI21X1
XOAI21X1_381 BUFX4_325/Y INVX4_24/Y OAI21X1_381/C gnd OAI21X1_381/Y vdd OAI21X1
XAND2X2_4 bundleStartMajId_i[43] bundleStartMajId_i[40] gnd AND2X2_4/Y vdd AND2X2
XOAI21X1_392 bundleStartMajId_i[63] BUFX4_237/Y OAI21X1_392/C gnd OAI21X1_392/Y vdd
+ OAI21X1
XFILL_1_OAI21X1_1319 gnd vdd FILL
XFILL_1_OAI21X1_1308 gnd vdd FILL
XFILL_1_DFFPOSX1_909 gnd vdd FILL
XFILL_6_DFFPOSX1_546 gnd vdd FILL
XFILL_6_DFFPOSX1_568 gnd vdd FILL
XFILL_6_DFFPOSX1_557 gnd vdd FILL
XFILL_6_DFFPOSX1_579 gnd vdd FILL
XFILL_7_10_0 gnd vdd FILL
XFILL_0_NAND2X1_116 gnd vdd FILL
XFILL_0_NAND2X1_105 gnd vdd FILL
XFILL_0_INVX1_130 gnd vdd FILL
XFILL_0_NAND2X1_138 gnd vdd FILL
XFILL_0_NAND2X1_127 gnd vdd FILL
XFILL_0_NAND2X1_149 gnd vdd FILL
XFILL_1_AOI21X1_41 gnd vdd FILL
XFILL_0_INVX1_152 gnd vdd FILL
XFILL_0_INVX1_141 gnd vdd FILL
XFILL_0_INVX1_163 gnd vdd FILL
XFILL_1_AOI21X1_30 gnd vdd FILL
XFILL_33_8_0 gnd vdd FILL
XFILL_0_INVX1_185 gnd vdd FILL
XFILL_1_AOI21X1_52 gnd vdd FILL
XFILL_0_INVX1_196 gnd vdd FILL
XFILL_1_AOI21X1_63 gnd vdd FILL
XFILL_0_INVX1_174 gnd vdd FILL
XFILL_5_DFFPOSX1_114 gnd vdd FILL
XFILL_5_DFFPOSX1_125 gnd vdd FILL
XFILL_5_DFFPOSX1_103 gnd vdd FILL
XFILL_5_DFFPOSX1_147 gnd vdd FILL
XFILL_5_DFFPOSX1_136 gnd vdd FILL
XFILL_5_DFFPOSX1_158 gnd vdd FILL
XFILL_5_DFFPOSX1_169 gnd vdd FILL
XOAI21X1_1622 INVX2_125/Y BUFX4_193/Y NAND2X1_690/Y gnd DFFPOSX1_12/D vdd OAI21X1
XOAI21X1_1600 BUFX4_321/Y INVX2_136/Y NAND2X1_669/Y gnd OAI21X1_1600/Y vdd OAI21X1
XOAI21X1_1633 INVX2_136/Y BUFX4_233/Y NAND2X1_701/Y gnd DFFPOSX1_23/D vdd OAI21X1
XOAI21X1_1611 BUFX4_373/Y INVX2_115/Y NAND2X1_680/Y gnd DFFPOSX1_2/D vdd OAI21X1
XOAI21X1_1666 BUFX4_105/Y BUFX4_339/Y BUFX2_715/A gnd OAI21X1_1667/C vdd OAI21X1
XOAI21X1_1655 BUFX4_125/Y INVX2_121/Y OAI21X1_1655/C gnd DFFPOSX1_40/D vdd OAI21X1
XFILL_1_OAI21X1_1820 gnd vdd FILL
XOAI21X1_1644 INVX2_115/Y BUFX4_225/Y NAND2X1_712/Y gnd DFFPOSX1_34/D vdd OAI21X1
XOAI21X1_1688 BUFX4_2/A BUFX4_352/Y BUFX2_727/A gnd OAI21X1_1689/C vdd OAI21X1
XOAI21X1_1677 BUFX4_170/Y INVX2_132/Y OAI21X1_1677/C gnd DFFPOSX1_51/D vdd OAI21X1
XOAI21X1_1699 BUFX4_140/Y INVX2_143/Y OAI21X1_1699/C gnd DFFPOSX1_62/D vdd OAI21X1
XFILL_0_OAI21X1_611 gnd vdd FILL
XFILL_0_OAI21X1_600 gnd vdd FILL
XFILL_0_OAI21X1_622 gnd vdd FILL
XFILL_0_OAI21X1_655 gnd vdd FILL
XFILL_0_OAI21X1_644 gnd vdd FILL
XFILL_1_OAI21X1_837 gnd vdd FILL
XFILL_1_OAI21X1_826 gnd vdd FILL
XFILL_1_OAI21X1_804 gnd vdd FILL
XFILL_0_OAI21X1_633 gnd vdd FILL
XFILL_2_OAI22X1_2 gnd vdd FILL
XFILL_1_OAI21X1_815 gnd vdd FILL
XFILL_0_OAI21X1_666 gnd vdd FILL
XFILL_1_OAI21X1_848 gnd vdd FILL
XFILL_1_OAI21X1_859 gnd vdd FILL
XFILL_0_OAI21X1_699 gnd vdd FILL
XFILL_0_OAI21X1_688 gnd vdd FILL
XFILL_0_OAI21X1_677 gnd vdd FILL
XFILL_1_AND2X2_23 gnd vdd FILL
XFILL_1_AND2X2_12 gnd vdd FILL
XFILL_3_DFFPOSX1_18 gnd vdd FILL
XFILL_3_DFFPOSX1_29 gnd vdd FILL
XFILL_13_16_0 gnd vdd FILL
XFILL_0_NAND2X1_650 gnd vdd FILL
XFILL_0_NAND2X1_672 gnd vdd FILL
XFILL_0_OAI21X1_1432 gnd vdd FILL
XFILL_0_OAI21X1_1421 gnd vdd FILL
XFILL_0_OAI21X1_1410 gnd vdd FILL
XFILL_0_NAND2X1_661 gnd vdd FILL
XFILL_0_NAND2X1_683 gnd vdd FILL
XFILL_0_OAI21X1_1465 gnd vdd FILL
XFILL_0_OAI21X1_1476 gnd vdd FILL
XFILL_24_8_0 gnd vdd FILL
XFILL_0_NAND2X1_694 gnd vdd FILL
XFILL_0_OAI21X1_1454 gnd vdd FILL
XFILL_0_OAI21X1_1443 gnd vdd FILL
XFILL_0_OAI21X1_1487 gnd vdd FILL
XFILL_0_OAI21X1_1498 gnd vdd FILL
XFILL_4_DFFPOSX1_5 gnd vdd FILL
XFILL_5_DFFPOSX1_670 gnd vdd FILL
XFILL_0_BUFX2_7 gnd vdd FILL
XFILL_5_DFFPOSX1_681 gnd vdd FILL
XFILL_5_DFFPOSX1_692 gnd vdd FILL
XFILL_0_BUFX2_409 gnd vdd FILL
XFILL_18_15_0 gnd vdd FILL
XFILL_7_9_0 gnd vdd FILL
XFILL_4_DFFPOSX1_271 gnd vdd FILL
XFILL_31_17_0 gnd vdd FILL
XFILL_0_NAND2X1_29 gnd vdd FILL
XFILL_2_OAI21X1_1537 gnd vdd FILL
XFILL_0_NAND2X1_18 gnd vdd FILL
XFILL_4_DFFPOSX1_260 gnd vdd FILL
XFILL_4_DFFPOSX1_282 gnd vdd FILL
XFILL_4_DFFPOSX1_293 gnd vdd FILL
XFILL_0_INVX2_7 gnd vdd FILL
XFILL_15_8_0 gnd vdd FILL
XFILL_1_BUFX2_161 gnd vdd FILL
XFILL_1_OAI21X1_1105 gnd vdd FILL
XFILL_1_BUFX2_172 gnd vdd FILL
XFILL_0_BUFX2_943 gnd vdd FILL
XFILL_0_BUFX2_932 gnd vdd FILL
XFILL_0_BUFX2_921 gnd vdd FILL
XFILL_1_OAI21X1_1116 gnd vdd FILL
XFILL_1_OAI21X1_1127 gnd vdd FILL
XDFFPOSX1_519 BUFX2_550/A CLKBUF1_90/Y OAI21X1_594/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_706 gnd vdd FILL
XFILL_0_BUFX2_910 gnd vdd FILL
XDFFPOSX1_508 BUFX2_538/A CLKBUF1_33/Y OAI21X1_565/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_1138 gnd vdd FILL
XFILL_0_BUFX2_976 gnd vdd FILL
XFILL_0_BUFX2_954 gnd vdd FILL
XINVX1_220 INVX1_220/A gnd INVX1_220/Y vdd INVX1
XFILL_1_OAI21X1_1149 gnd vdd FILL
XFILL_0_BUFX2_965 gnd vdd FILL
XFILL_1_DFFPOSX1_728 gnd vdd FILL
XFILL_1_DFFPOSX1_717 gnd vdd FILL
XFILL_1_DFFPOSX1_739 gnd vdd FILL
XFILL_0_BUFX2_987 gnd vdd FILL
XFILL_0_BUFX2_998 gnd vdd FILL
XFILL_6_DFFPOSX1_310 gnd vdd FILL
XFILL_6_DFFPOSX1_321 gnd vdd FILL
XFILL_6_DFFPOSX1_343 gnd vdd FILL
XFILL_6_DFFPOSX1_332 gnd vdd FILL
XFILL_36_16_0 gnd vdd FILL
XFILL_6_DFFPOSX1_354 gnd vdd FILL
XNAND2X1_42 BUFX2_869/A BUFX4_234/Y gnd OAI21X1_42/C vdd NAND2X1
XNAND2X1_20 BUFX2_845/A BUFX4_227/Y gnd OAI21X1_20/C vdd NAND2X1
XNAND2X1_31 BUFX2_857/A BUFX4_195/Y gnd OAI21X1_31/C vdd NAND2X1
XNAND2X1_64 BUFX2_893/A BUFX4_207/Y gnd OAI21X1_64/C vdd NAND2X1
XNAND2X1_53 BUFX2_881/A BUFX4_198/Y gnd OAI21X1_53/C vdd NAND2X1
XNAND2X1_75 BUFX2_416/A BUFX4_321/Y gnd NAND2X1_75/Y vdd NAND2X1
XNAND2X1_86 BUFX2_399/A BUFX4_335/Y gnd NAND2X1_86/Y vdd NAND2X1
XNAND2X1_97 BUFX2_411/A BUFX4_378/Y gnd NAND2X1_97/Y vdd NAND2X1
XFILL_0_XNOR2X1_71 gnd vdd FILL
XFILL_0_XNOR2X1_60 gnd vdd FILL
XFILL_0_XNOR2X1_93 gnd vdd FILL
XFILL_1_NAND2X1_128 gnd vdd FILL
XFILL_1_NAND2X1_117 gnd vdd FILL
XFILL_0_XNOR2X1_82 gnd vdd FILL
XFILL_1_NAND2X1_106 gnd vdd FILL
XFILL_0_DFFPOSX1_318 gnd vdd FILL
XFILL_0_DFFPOSX1_307 gnd vdd FILL
XFILL_0_DFFPOSX1_329 gnd vdd FILL
XFILL_1_NAND2X1_139 gnd vdd FILL
XFILL_0_NOR3X1_14 gnd vdd FILL
XOAI21X1_1430 INVX1_221/Y INVX2_67/Y INVX4_34/Y gnd OAI21X1_1431/C vdd OAI21X1
XOAI21X1_1441 BUFX4_174/Y BUFX4_31/Y BUFX2_204/A gnd OAI21X1_1442/C vdd OAI21X1
XFILL_1_OAI21X1_1650 gnd vdd FILL
XOAI21X1_1474 BUFX4_128/Y BUFX4_45/Y BUFX2_218/A gnd OAI21X1_1475/C vdd OAI21X1
XOAI21X1_1463 XNOR2X1_98/A INVX2_72/Y INVX1_176/Y gnd OAI21X1_1464/C vdd OAI21X1
XFILL_0_BUFX4_291 gnd vdd FILL
XFILL_0_BUFX4_280 gnd vdd FILL
XOAI21X1_1452 BUFX4_169/Y BUFX4_78/Y BUFX2_209/A gnd OAI21X1_1453/C vdd OAI21X1
XFILL_1_OAI21X1_1661 gnd vdd FILL
XFILL_1_OAI21X1_1694 gnd vdd FILL
XFILL_1_OAI21X1_1683 gnd vdd FILL
XFILL_1_OAI21X1_612 gnd vdd FILL
XFILL_1_OAI21X1_1672 gnd vdd FILL
XOAI21X1_1496 OAI21X1_1496/A BUFX4_294/Y OAI21X1_1496/C gnd OAI21X1_1496/Y vdd OAI21X1
XOAI21X1_1485 INVX1_223/A INVX4_40/Y INVX2_76/Y gnd OAI21X1_1486/C vdd OAI21X1
XFILL_1_OAI21X1_601 gnd vdd FILL
XFILL_0_OAI21X1_430 gnd vdd FILL
XFILL_1_OAI21X1_645 gnd vdd FILL
XFILL_1_NOR2X1_217 gnd vdd FILL
XFILL_1_OAI21X1_634 gnd vdd FILL
XFILL_0_OAI21X1_474 gnd vdd FILL
XFILL_1_NOR2X1_206 gnd vdd FILL
XFILL_0_OAI21X1_463 gnd vdd FILL
XFILL_1_OAI21X1_623 gnd vdd FILL
XFILL_1_NOR2X1_228 gnd vdd FILL
XFILL_0_OAI21X1_452 gnd vdd FILL
XFILL_0_OAI21X1_441 gnd vdd FILL
XFILL_1_OAI21X1_656 gnd vdd FILL
XFILL_0_OAI21X1_496 gnd vdd FILL
XFILL_3_NOR3X1_7 gnd vdd FILL
XFILL_1_OAI21X1_667 gnd vdd FILL
XFILL_0_OAI21X1_485 gnd vdd FILL
XFILL_1_OAI21X1_678 gnd vdd FILL
XFILL_1_OAI21X1_689 gnd vdd FILL
XFILL_4_DFFPOSX1_19 gnd vdd FILL
XFILL_0_OAI21X1_1251 gnd vdd FILL
XFILL_0_OAI21X1_1240 gnd vdd FILL
XFILL_0_NAND2X1_480 gnd vdd FILL
XFILL_1_NAND2X1_673 gnd vdd FILL
XFILL_0_NAND2X1_491 gnd vdd FILL
XFILL_1_NAND2X1_684 gnd vdd FILL
XFILL_0_DFFPOSX1_841 gnd vdd FILL
XFILL_0_DFFPOSX1_852 gnd vdd FILL
XFILL_0_OAI21X1_1284 gnd vdd FILL
XFILL_1_NAND2X1_662 gnd vdd FILL
XFILL_0_OAI21X1_1262 gnd vdd FILL
XFILL_0_OAI21X1_1273 gnd vdd FILL
XFILL_0_DFFPOSX1_830 gnd vdd FILL
XFILL_0_DFFPOSX1_874 gnd vdd FILL
XFILL_0_OAI21X1_1295 gnd vdd FILL
XFILL_0_DFFPOSX1_885 gnd vdd FILL
XFILL_0_DFFPOSX1_863 gnd vdd FILL
XDFFPOSX1_1004 BUFX2_649/A CLKBUF1_8/Y OAI21X1_1581/Y gnd vdd DFFPOSX1
XDFFPOSX1_1026 BUFX2_664/A CLKBUF1_43/Y OAI21X1_1603/Y gnd vdd DFFPOSX1
XDFFPOSX1_1015 BUFX2_652/A CLKBUF1_64/Y OAI21X1_1592/Y gnd vdd DFFPOSX1
XFILL_0_DFFPOSX1_896 gnd vdd FILL
XFILL_0_BUFX2_217 gnd vdd FILL
XFILL_0_BUFX2_206 gnd vdd FILL
XFILL_0_BUFX2_228 gnd vdd FILL
XFILL_20_14_1 gnd vdd FILL
XOAI22X1_2 INVX2_48/Y OR2X2_9/A OAI22X1_2/C bundleStartMajId_i[27] gnd OAI22X1_2/Y
+ vdd OAI22X1
XFILL_0_BUFX2_239 gnd vdd FILL
XFILL_0_AOI21X1_60 gnd vdd FILL
XFILL_2_OAI21X1_1301 gnd vdd FILL
XFILL_2_DFFPOSX1_902 gnd vdd FILL
XFILL_2_DFFPOSX1_924 gnd vdd FILL
XFILL_2_DFFPOSX1_913 gnd vdd FILL
XFILL_2_DFFPOSX1_946 gnd vdd FILL
XFILL_2_DFFPOSX1_935 gnd vdd FILL
XFILL_2_DFFPOSX1_957 gnd vdd FILL
XFILL_2_DFFPOSX1_968 gnd vdd FILL
XFILL_2_DFFPOSX1_979 gnd vdd FILL
XFILL_30_6_0 gnd vdd FILL
XFILL_25_13_1 gnd vdd FILL
XFILL_3_XNOR2X1_37 gnd vdd FILL
XFILL_3_XNOR2X1_26 gnd vdd FILL
XDFFPOSX1_316 BUFX2_986/A CLKBUF1_43/Y OAI21X1_249/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_751 gnd vdd FILL
XFILL_3_XNOR2X1_59 gnd vdd FILL
XDFFPOSX1_327 BUFX2_998/A CLKBUF1_22/Y OAI21X1_271/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_503 gnd vdd FILL
XFILL_1_DFFPOSX1_514 gnd vdd FILL
XDFFPOSX1_338 BUFX2_1010/A CLKBUF1_4/Y OAI21X1_293/Y gnd vdd DFFPOSX1
XDFFPOSX1_305 BUFX2_974/A CLKBUF1_66/Y OAI21X1_227/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_740 gnd vdd FILL
XFILL_0_BUFX2_784 gnd vdd FILL
XFILL_0_BUFX2_762 gnd vdd FILL
XFILL_1_DFFPOSX1_547 gnd vdd FILL
XDFFPOSX1_349 BUFX2_1022/A CLKBUF1_47/Y OAI21X1_315/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_525 gnd vdd FILL
XFILL_1_DFFPOSX1_536 gnd vdd FILL
XFILL_0_NOR2X1_80 gnd vdd FILL
XFILL_0_NOR2X1_91 gnd vdd FILL
XFILL_0_BUFX2_773 gnd vdd FILL
XFILL_0_BUFX2_795 gnd vdd FILL
XNAND2X1_408 BUFX2_57/A BUFX4_347/Y gnd NAND2X1_408/Y vdd NAND2X1
XFILL_1_DFFPOSX1_569 gnd vdd FILL
XFILL_1_DFFPOSX1_558 gnd vdd FILL
XNAND2X1_419 BUFX2_10/A BUFX4_359/Y gnd NAND2X1_419/Y vdd NAND2X1
XFILL_3_DFFPOSX1_2 gnd vdd FILL
XFILL_6_DFFPOSX1_195 gnd vdd FILL
XFILL_38_7_0 gnd vdd FILL
XBUFX4_381 BUFX4_381/A gnd BUFX4_381/Y vdd BUFX4
XBUFX4_370 BUFX4_384/A gnd BUFX4_370/Y vdd BUFX4
XFILL_0_DFFPOSX1_104 gnd vdd FILL
XFILL_0_14_1 gnd vdd FILL
XFILL_0_DFFPOSX1_126 gnd vdd FILL
XFILL_0_DFFPOSX1_115 gnd vdd FILL
XFILL_0_DFFPOSX1_137 gnd vdd FILL
XFILL_0_DFFPOSX1_148 gnd vdd FILL
XFILL_1_BUFX2_908 gnd vdd FILL
XFILL_0_DFFPOSX1_159 gnd vdd FILL
XOAI21X1_914 BUFX4_100/Y BUFX4_329/Y BUFX2_348/A gnd OAI21X1_915/C vdd OAI21X1
XOAI21X1_925 BUFX4_143/Y INVX1_117/Y OAI21X1_925/C gnd OAI21X1_925/Y vdd OAI21X1
XFILL_21_6_0 gnd vdd FILL
XFILL_0_NAND2X1_2 gnd vdd FILL
XOAI21X1_903 INVX1_104/Y BUFX4_181/Y OAI21X1_903/C gnd OAI21X1_903/Y vdd OAI21X1
XOAI21X1_936 BUFX4_247/Y BUFX4_329/Y BUFX2_331/A gnd OAI21X1_937/C vdd OAI21X1
XFILL_3_DFFPOSX1_608 gnd vdd FILL
XFILL_3_DFFPOSX1_619 gnd vdd FILL
XOAI21X1_958 BUFX4_1/A OAI21X1_7/A BUFX2_343/A gnd OAI21X1_959/C vdd OAI21X1
XOAI21X1_947 BUFX4_154/Y INVX1_128/Y OAI21X1_947/C gnd OAI21X1_947/Y vdd OAI21X1
XOAI21X1_969 BUFX4_123/Y INVX1_139/Y OAI21X1_969/C gnd OAI21X1_969/Y vdd OAI21X1
XOAI21X1_1260 NOR2X1_184/B NOR2X1_185/B BUFX4_305/Y gnd OAI21X1_1261/B vdd OAI21X1
XOAI21X1_1282 XNOR2X1_79/Y BUFX4_159/Y OAI21X1_1282/C gnd OAI21X1_1282/Y vdd OAI21X1
XDFFPOSX1_850 BUFX2_102/A CLKBUF1_85/Y OAI21X1_1169/Y gnd vdd DFFPOSX1
XOAI21X1_1271 OAI21X1_1271/A BUFX4_129/Y OAI21X1_1271/C gnd OAI21X1_1271/Y vdd OAI21X1
XDFFPOSX1_883 BUFX2_132/A CLKBUF1_11/Y OAI21X1_1237/Y gnd vdd DFFPOSX1
XDFFPOSX1_872 BUFX2_129/A CLKBUF1_7/Y OAI21X1_1209/Y gnd vdd DFFPOSX1
XOAI21X1_1293 BUFX4_103/Y BUFX4_339/Y BUFX2_154/A gnd OAI21X1_1294/C vdd OAI21X1
XFILL_1_OAI21X1_1480 gnd vdd FILL
XFILL_1_OAI21X1_1491 gnd vdd FILL
XFILL_1_OAI21X1_420 gnd vdd FILL
XINVX2_11 bundleStartMajId_i[59] gnd INVX2_11/Y vdd INVX2
XDFFPOSX1_861 BUFX2_114/A CLKBUF1_76/Y OAI21X1_1187/Y gnd vdd DFFPOSX1
XFILL_0_OAI21X1_260 gnd vdd FILL
XFILL_0_OAI21X1_282 gnd vdd FILL
XINVX2_33 bundleStartMajId_i[13] gnd INVX2_33/Y vdd INVX2
XFILL_0_OAI21X1_271 gnd vdd FILL
XINVX2_44 INVX2_44/A gnd NOR3X1_2/B vdd INVX2
XDFFPOSX1_894 BUFX2_144/A CLKBUF1_83/Y OAI21X1_1274/Y gnd vdd DFFPOSX1
XINVX2_22 bundleStartMajId_i[37] gnd INVX2_22/Y vdd INVX2
XFILL_1_OAI21X1_453 gnd vdd FILL
XFILL_1_OAI21X1_431 gnd vdd FILL
XFILL_1_OAI21X1_442 gnd vdd FILL
XFILL_2_OAI21X1_657 gnd vdd FILL
XFILL_2_OAI21X1_646 gnd vdd FILL
XINVX2_66 bundleAddress_i[49] gnd INVX2_66/Y vdd INVX2
XINVX2_55 bundleAddress_i[62] gnd INVX2_55/Y vdd INVX2
XFILL_1_OAI21X1_486 gnd vdd FILL
XFILL_1_OAI21X1_475 gnd vdd FILL
XFILL_1_OAI21X1_464 gnd vdd FILL
XFILL_0_OAI21X1_293 gnd vdd FILL
XINVX2_88 bundleAddress_i[7] gnd INVX2_88/Y vdd INVX2
XINVX2_77 bundleAddress_i[27] gnd INVX2_77/Y vdd INVX2
XINVX2_99 INVX2_99/A gnd INVX2_99/Y vdd INVX2
XFILL_1_OAI21X1_497 gnd vdd FILL
XFILL_5_13_1 gnd vdd FILL
XFILL_2_DFFPOSX1_209 gnd vdd FILL
XBUFX2_318 BUFX2_318/A gnd instr2_o[0] vdd BUFX2
XFILL_29_7_0 gnd vdd FILL
XFILL_0_AOI21X1_7 gnd vdd FILL
XBUFX2_307 BUFX2_307/A gnd instr2_o[10] vdd BUFX2
XFILL_4_7_0 gnd vdd FILL
XBUFX2_329 BUFX2_329/A gnd instr3_o[19] vdd BUFX2
XFILL_1_INVX4_33 gnd vdd FILL
XFILL_1_INVX4_22 gnd vdd FILL
XFILL_1_BUFX4_212 gnd vdd FILL
XFILL_1_BUFX4_201 gnd vdd FILL
XFILL_1_BUFX4_234 gnd vdd FILL
XFILL_0_DFFPOSX1_660 gnd vdd FILL
XFILL_1_NAND2X1_492 gnd vdd FILL
XFILL_1_NAND2X1_470 gnd vdd FILL
XFILL_1_BUFX4_223 gnd vdd FILL
XOAI21X1_29 INVX2_167/Y BUFX4_200/Y OAI21X1_29/C gnd OAI21X1_29/Y vdd OAI21X1
XFILL_0_OAI21X1_1081 gnd vdd FILL
XFILL_0_OAI21X1_1070 gnd vdd FILL
XFILL_1_BUFX4_245 gnd vdd FILL
XOAI21X1_18 INVX2_156/Y OAI21X1_9/B OAI21X1_18/C gnd OAI21X1_18/Y vdd OAI21X1
XFILL_0_OAI21X1_1092 gnd vdd FILL
XFILL_1_BUFX4_289 gnd vdd FILL
XFILL_1_BUFX4_278 gnd vdd FILL
XFILL_1_BUFX4_256 gnd vdd FILL
XFILL_1_BUFX4_267 gnd vdd FILL
XFILL_12_6_0 gnd vdd FILL
XFILL_0_DFFPOSX1_693 gnd vdd FILL
XFILL_0_DFFPOSX1_671 gnd vdd FILL
XFILL_0_DFFPOSX1_682 gnd vdd FILL
XFILL_0_DFFPOSX1_16 gnd vdd FILL
XFILL_0_DFFPOSX1_27 gnd vdd FILL
XFILL_0_DFFPOSX1_38 gnd vdd FILL
XFILL_2_BUFX4_72 gnd vdd FILL
XFILL_0_DFFPOSX1_49 gnd vdd FILL
XFILL_2_XNOR2X1_5 gnd vdd FILL
XBUFX2_830 NAND2X1_1/A gnd tid1_o[6] vdd BUFX2
XFILL_2_DFFPOSX1_710 gnd vdd FILL
XFILL_2_DFFPOSX1_721 gnd vdd FILL
XFILL_2_DFFPOSX1_732 gnd vdd FILL
XFILL_2_OAI21X1_1142 gnd vdd FILL
XBUFX2_841 NAND2X1_8/A gnd tid2_o[63] vdd BUFX2
XBUFX2_852 BUFX2_852/A gnd tid2_o[44] vdd BUFX2
XFILL_2_DFFPOSX1_754 gnd vdd FILL
XFILL_2_DFFPOSX1_743 gnd vdd FILL
XBUFX2_863 BUFX2_863/A gnd tid2_o[34] vdd BUFX2
XFILL_2_DFFPOSX1_765 gnd vdd FILL
XBUFX2_885 BUFX2_885/A gnd tid2_o[14] vdd BUFX2
XFILL_2_DFFPOSX1_776 gnd vdd FILL
XFILL_2_DFFPOSX1_787 gnd vdd FILL
XFILL_0_NOR2X1_203 gnd vdd FILL
XBUFX2_874 BUFX2_874/A gnd tid2_o[24] vdd BUFX2
XBUFX2_896 BUFX2_896/A gnd tid2_o[4] vdd BUFX2
XFILL_2_DFFPOSX1_798 gnd vdd FILL
XFILL_0_NOR2X1_225 gnd vdd FILL
XFILL_0_NOR2X1_214 gnd vdd FILL
XFILL_12_2 gnd vdd FILL
XFILL_3_CLKBUF1_5 gnd vdd FILL
XDFFPOSX1_102 BUFX2_789/A CLKBUF1_92/Y OAI21X1_1776/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_322 gnd vdd FILL
XDFFPOSX1_124 BUFX2_794/A CLKBUF1_93/Y OAI21X1_1798/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_311 gnd vdd FILL
XDFFPOSX1_135 BUFX2_806/A CLKBUF1_73/Y OAI21X1_1809/Y gnd vdd DFFPOSX1
XFILL_1_DFFPOSX1_300 gnd vdd FILL
XDFFPOSX1_146 BUFX2_818/A CLKBUF1_41/Y OAI21X1_1820/Y gnd vdd DFFPOSX1
XDFFPOSX1_113 BUFX2_782/A CLKBUF1_56/Y OAI21X1_1787/Y gnd vdd DFFPOSX1
XDFFPOSX1_157 NAND2X1_1/A CLKBUF1_43/Y OAI21X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_179 BUFX2_848/A CLKBUF1_12/Y OAI21X1_23/Y gnd vdd DFFPOSX1
XDFFPOSX1_168 BUFX2_875/A CLKBUF1_101/Y OAI21X1_12/Y gnd vdd DFFPOSX1
XFILL_0_BUFX2_581 gnd vdd FILL
XFILL_0_BUFX2_570 gnd vdd FILL
XFILL_1_DFFPOSX1_333 gnd vdd FILL
XFILL_0_BUFX2_592 gnd vdd FILL
XFILL_1_DFFPOSX1_366 gnd vdd FILL
XFILL_1_DFFPOSX1_355 gnd vdd FILL
XFILL_1_DFFPOSX1_344 gnd vdd FILL
XFILL_1_DFFPOSX1_399 gnd vdd FILL
XNAND2X1_216 bundleStartMajId_i[25] bundleStartMajId_i[24] gnd NOR2X1_34/B vdd NAND2X1
XFILL_1_DFFPOSX1_388 gnd vdd FILL
XFILL_1_DFFPOSX1_377 gnd vdd FILL
XNAND2X1_205 BUFX2_484/A BUFX4_182/Y gnd OAI21X1_450/C vdd NAND2X1
XNAND2X1_238 bundleStartMajId_i[15] bundleStartMajId_i[14] gnd NOR2X1_44/A vdd NAND2X1
XNAND2X1_249 bundleStartMajId_i[8] INVX2_46/A gnd INVX1_21/A vdd NAND2X1
XFILL_4_DFFPOSX1_804 gnd vdd FILL
XNAND2X1_227 BUFX2_497/A BUFX4_225/Y gnd OAI21X1_467/C vdd NAND2X1
XFILL_4_DFFPOSX1_815 gnd vdd FILL
XFILL_4_DFFPOSX1_837 gnd vdd FILL
XFILL_16_18_1 gnd vdd FILL
XFILL_4_DFFPOSX1_826 gnd vdd FILL
XFILL_4_DFFPOSX1_848 gnd vdd FILL
XFILL_4_DFFPOSX1_859 gnd vdd FILL
XFILL_4_CLKBUF1_60 gnd vdd FILL
XFILL_10_14_0 gnd vdd FILL
XFILL_4_CLKBUF1_93 gnd vdd FILL
XFILL_0_BUFX2_20 gnd vdd FILL
XFILL_4_CLKBUF1_71 gnd vdd FILL
XFILL_0_BUFX2_42 gnd vdd FILL
XFILL_1_NOR2X1_12 gnd vdd FILL
XFILL_0_BUFX2_53 gnd vdd FILL
XFILL_0_BUFX2_31 gnd vdd FILL
XFILL_0_BUFX2_64 gnd vdd FILL
XFILL_1_NOR2X1_45 gnd vdd FILL
XFILL_0_BUFX2_97 gnd vdd FILL
XFILL_1_BUFX2_705 gnd vdd FILL
XFILL_0_BUFX2_86 gnd vdd FILL
XFILL_0_BUFX2_75 gnd vdd FILL
XFILL_1_NOR2X1_56 gnd vdd FILL
XOAI21X1_711 AOI21X1_31/Y OAI21X1_711/B OAI21X1_711/C gnd OAI21X1_711/Y vdd OAI21X1
XFILL_1_BUFX2_749 gnd vdd FILL
XOAI21X1_733 OAI21X1_733/A BUFX4_295/Y OAI21X1_733/C gnd OAI21X1_733/Y vdd OAI21X1
XOAI21X1_722 NOR2X1_69/A INVX1_37/A OAI21X1_722/C gnd OAI21X1_724/A vdd OAI21X1
XFILL_1_BUFX2_738 gnd vdd FILL
XOAI21X1_700 OAI21X1_700/A BUFX4_299/Y OAI21X1_700/C gnd OAI21X1_700/Y vdd OAI21X1
XFILL_3_DFFPOSX1_416 gnd vdd FILL
XOAI21X1_744 BUFX4_127/Y BUFX4_64/Y BUFX2_609/A gnd OAI21X1_745/C vdd OAI21X1
XFILL_3_DFFPOSX1_405 gnd vdd FILL
XOAI21X1_766 AND2X2_21/Y NOR2X1_113/Y BUFX4_287/Y gnd OAI21X1_767/C vdd OAI21X1
XOAI21X1_755 NOR2X1_110/Y bundleStartMajId_i[29] BUFX4_285/Y gnd OAI21X1_757/B vdd
+ OAI21X1
XFILL_3_DFFPOSX1_427 gnd vdd FILL
XOAI21X1_799 OAI21X1_799/A BUFX4_290/Y OAI21X1_799/C gnd OAI21X1_799/Y vdd OAI21X1
XOAI21X1_777 BUFX4_135/Y BUFX4_72/A BUFX2_622/A gnd OAI21X1_778/C vdd OAI21X1
XOAI21X1_788 BUFX4_142/Y BUFX4_74/Y BUFX2_625/A gnd OAI21X1_789/C vdd OAI21X1
XFILL_3_DFFPOSX1_449 gnd vdd FILL
XFILL_3_DFFPOSX1_438 gnd vdd FILL
XOAI21X1_1090 BUFX4_374/Y INVX2_87/Y NAND2X1_456/Y gnd OAI21X1_1090/Y vdd OAI21X1
XDFFPOSX1_691 BUFX2_328/A CLKBUF1_32/Y OAI21X1_931/Y gnd vdd DFFPOSX1
XDFFPOSX1_680 BUFX2_325/A CLKBUF1_101/Y OAI21X1_909/Y gnd vdd DFFPOSX1
XFILL_1_OAI21X1_261 gnd vdd FILL
XFILL_1_OAI21X1_250 gnd vdd FILL
XFILL_1_OAI21X1_294 gnd vdd FILL
XFILL_1_OAI21X1_272 gnd vdd FILL
XFILL_1_OAI21X1_283 gnd vdd FILL
XNAND2X1_750 BUFX2_806/A BUFX4_376/Y gnd NAND2X1_750/Y vdd NAND2X1
XNAND2X1_761 BUFX2_818/A OAI21X1_6/A gnd NAND2X1_761/Y vdd NAND2X1
XFILL_2_XNOR2X1_23 gnd vdd FILL
XFILL_2_OAI21X1_487 gnd vdd FILL
XFILL_2_XNOR2X1_12 gnd vdd FILL
XFILL_15_13_0 gnd vdd FILL
XBUFX2_126 BUFX2_126/A gnd addr2_o[56] vdd BUFX2
XFILL_2_XNOR2X1_56 gnd vdd FILL
XBUFX2_104 BUFX2_104/A gnd addr2_o[19] vdd BUFX2
XFILL_2_XNOR2X1_45 gnd vdd FILL
XBUFX2_115 BUFX2_115/A gnd addr2_o[9] vdd BUFX2
XFILL_2_XNOR2X1_34 gnd vdd FILL
XBUFX2_137 BUFX2_137/A gnd addr3_o[47] vdd BUFX2
XBUFX2_148 BUFX2_148/A gnd addr3_o[37] vdd BUFX2
XFILL_2_XNOR2X1_89 gnd vdd FILL
XFILL_2_XNOR2X1_78 gnd vdd FILL
XBUFX2_159 BUFX2_159/A gnd addr3_o[27] vdd BUFX2
XFILL_2_XNOR2X1_67 gnd vdd FILL
XFILL_0_CLKBUF1_102 gnd vdd FILL
XFILL_0_DFFPOSX1_490 gnd vdd FILL
XBUFX2_1018 BUFX2_1018/A gnd tid4_o[10] vdd BUFX2
XBUFX2_1007 BUFX2_1007/A gnd tid4_o[20] vdd BUFX2
XFILL_3_DFFPOSX1_950 gnd vdd FILL
XFILL_3_DFFPOSX1_961 gnd vdd FILL
XFILL_3_DFFPOSX1_983 gnd vdd FILL
XFILL_3_DFFPOSX1_972 gnd vdd FILL
XBUFX2_1029 BUFX2_1029/A gnd tid4_o[0] vdd BUFX2
XFILL_3_DFFPOSX1_994 gnd vdd FILL
XCLKBUF1_19 BUFX4_91/Y gnd CLKBUF1_19/Y vdd CLKBUF1
XFILL_1_DFFPOSX1_39 gnd vdd FILL
XFILL_1_DFFPOSX1_17 gnd vdd FILL
XFILL_1_DFFPOSX1_28 gnd vdd FILL
XFILL_33_14_0 gnd vdd FILL
XBUFX4_40 BUFX4_67/A gnd BUFX4_40/Y vdd BUFX4
XBUFX4_62 BUFX4_82/A gnd BUFX4_62/Y vdd BUFX4
XBUFX4_51 BUFX4_51/A gnd BUFX4_51/Y vdd BUFX4
XBUFX4_95 BUFX4_95/A gnd BUFX4_95/Y vdd BUFX4
XBUFX4_84 clock_i gnd BUFX4_84/Y vdd BUFX4
XBUFX4_73 BUFX4_73/A gnd BUFX4_73/Y vdd BUFX4
XFILL_35_5_0 gnd vdd FILL
XFILL_0_OAI21X1_1817 gnd vdd FILL
XFILL_2_DFFPOSX1_540 gnd vdd FILL
XFILL_0_OAI21X1_1806 gnd vdd FILL
XBUFX2_682 BUFX2_682/A gnd pid2_o[30] vdd BUFX2
XFILL_0_OAI21X1_1828 gnd vdd FILL
XFILL_2_DFFPOSX1_551 gnd vdd FILL
XBUFX2_671 BUFX2_671/A gnd pid1_o[2] vdd BUFX2
XBUFX2_660 BUFX2_660/A gnd pid1_o[12] vdd BUFX2
XFILL_2_DFFPOSX1_573 gnd vdd FILL
XFILL_2_DFFPOSX1_562 gnd vdd FILL
XFILL_2_DFFPOSX1_595 gnd vdd FILL
XFILL_2_DFFPOSX1_584 gnd vdd FILL
XBUFX2_693 BUFX2_693/A gnd pid2_o[29] vdd BUFX2
XOR2X2_21 OR2X2_21/A OR2X2_21/B gnd OR2X2_21/Y vdd OR2X2
XOR2X2_10 OR2X2_10/A OR2X2_10/B gnd OR2X2_10/Y vdd OR2X2
XFILL_1_DFFPOSX1_130 gnd vdd FILL
XFILL_2_AOI21X1_34 gnd vdd FILL
XOR2X2_3 OR2X2_5/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XFILL_38_13_0 gnd vdd FILL
XFILL_1_DFFPOSX1_163 gnd vdd FILL
XFILL_1_DFFPOSX1_152 gnd vdd FILL
XFILL_1_DFFPOSX1_174 gnd vdd FILL
XXNOR2X1_5 NOR2X1_9/Y bundleStartMajId_i[48] gnd XNOR2X1_5/Y vdd XNOR2X1
XFILL_1_DFFPOSX1_141 gnd vdd FILL
XFILL_1_DFFPOSX1_185 gnd vdd FILL
XFILL_1_DFFPOSX1_196 gnd vdd FILL
XFILL_4_DFFPOSX1_601 gnd vdd FILL
XFILL_4_DFFPOSX1_612 gnd vdd FILL
XFILL_4_DFFPOSX1_645 gnd vdd FILL
XFILL_4_DFFPOSX1_634 gnd vdd FILL
XFILL_4_DFFPOSX1_623 gnd vdd FILL
XFILL_4_DFFPOSX1_656 gnd vdd FILL
XFILL_4_DFFPOSX1_678 gnd vdd FILL
XFILL_4_DFFPOSX1_667 gnd vdd FILL
XFILL_4_DFFPOSX1_689 gnd vdd FILL
XFILL_26_5_0 gnd vdd FILL
XFILL_1_5_0 gnd vdd FILL
XFILL_1_BUFX2_502 gnd vdd FILL
XFILL_1_BUFX2_546 gnd vdd FILL
XINVX1_5 bundleStartMajId_i[1] gnd INVX1_5/Y vdd INVX1
XFILL_1_BUFX2_535 gnd vdd FILL
XFILL_1_BUFX2_513 gnd vdd FILL
XFILL_3_DFFPOSX1_202 gnd vdd FILL
XFILL_1_BUFX2_557 gnd vdd FILL
XFILL_0_BUFX4_109 gnd vdd FILL
XOAI21X1_541 OAI21X1_541/A BUFX4_135/Y OAI21X1_541/C gnd OAI21X1_541/Y vdd OAI21X1
XFILL_10_9_1 gnd vdd FILL
XOAI21X1_530 OAI21X1_530/A BUFX4_163/Y OAI21X1_530/C gnd OAI21X1_530/Y vdd OAI21X1
XFILL_3_DFFPOSX1_246 gnd vdd FILL
XFILL_3_DFFPOSX1_213 gnd vdd FILL
XFILL_3_DFFPOSX1_235 gnd vdd FILL
XOAI21X1_552 OAI21X1_552/A BUFX4_130/Y OAI21X1_552/C gnd OAI21X1_552/Y vdd OAI21X1
XOAI21X1_563 XNOR2X1_30/Y BUFX4_130/Y OAI21X1_563/C gnd OAI21X1_563/Y vdd OAI21X1
XFILL_3_DFFPOSX1_224 gnd vdd FILL
XOAI21X1_574 NOR2X1_71/Y OAI21X1_574/B OAI21X1_574/C gnd OAI21X1_574/Y vdd OAI21X1
XOAI21X1_596 OAI22X1_2/Y BUFX4_155/Y OAI21X1_596/C gnd OAI21X1_596/Y vdd OAI21X1
XFILL_3_DFFPOSX1_279 gnd vdd FILL
XFILL_3_DFFPOSX1_268 gnd vdd FILL
XFILL_3_DFFPOSX1_257 gnd vdd FILL
XOAI21X1_585 BUFX4_93/Y BUFX4_335/Y BUFX2_548/A gnd OAI21X1_586/C vdd OAI21X1
.ends

