module BundleParser (clock_i, enable_i, bundle_i, bundleAddress_i, bundleLen_i, is64Bit_i, bundlePid_i, bundleTid_i, bundleStartMajId_i, enable1_i, enable2_i, enable3_i, enable4_i, enable1_o, enable2_o, enable3_o, enable4_o, instr1_o, instr2_o, instr3_o, instr4_o, addr1_o, addr2_o, addr3_o, addr4_o, is64b1_o, is64b2_o, is64b3_o, is64b4_o, pid1_o, pid2_o, pid3_o, pid4_o, tid1_o, tid2_o, tid3_o, tid4_o, majID1_o, majID2_o, majID3_o, majID4_o);

input clock_i;
input enable_i;
input is64Bit_i;
input enable1_i;
input enable2_i;
input enable3_i;
input enable4_i;
output enable1_o;
output enable2_o;
output enable3_o;
output enable4_o;
output is64b1_o;
output is64b2_o;
output is64b3_o;
output is64b4_o;
input [127:0] bundle_i;
input [63:0] bundleAddress_i;
input [1:0] bundleLen_i;
input [31:0] bundlePid_i;
input [63:0] bundleTid_i;
input [63:0] bundleStartMajId_i;
output [31:0] instr1_o;
output [31:0] instr2_o;
output [31:0] instr3_o;
output [31:0] instr4_o;
output [63:0] addr1_o;
output [63:0] addr2_o;
output [63:0] addr3_o;
output [63:0] addr4_o;
output [31:0] pid1_o;
output [31:0] pid2_o;
output [31:0] pid3_o;
output [31:0] pid4_o;
output [63:0] tid1_o;
output [63:0] tid2_o;
output [63:0] tid3_o;
output [63:0] tid4_o;
output [63:0] majID1_o;
output [63:0] majID2_o;
output [63:0] majID3_o;
output [63:0] majID4_o;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX4 BUFX4_1 ( .A(_1100__bF_buf2), .Y(_1100__bF_buf7_bF_buf3) );
BUFX4 BUFX4_2 ( .A(_1100__bF_buf4), .Y(_1100__bF_buf7_bF_buf2) );
BUFX4 BUFX4_3 ( .A(_1100__bF_buf14), .Y(_1100__bF_buf7_bF_buf1) );
BUFX4 BUFX4_4 ( .A(_1100__bF_buf5), .Y(_1100__bF_buf7_bF_buf0) );
BUFX4 BUFX4_5 ( .A(_1100__bF_buf1), .Y(_1100__bF_buf8_bF_buf3) );
BUFX4 BUFX4_6 ( .A(_1100__bF_buf1), .Y(_1100__bF_buf8_bF_buf2) );
BUFX4 BUFX4_7 ( .A(_1100__bF_buf6), .Y(_1100__bF_buf8_bF_buf1) );
BUFX4 BUFX4_8 ( .A(_1100__bF_buf11), .Y(_1100__bF_buf8_bF_buf0) );
BUFX4 BUFX4_9 ( .A(_1100__bF_buf8), .Y(_1100__bF_buf9_bF_buf3) );
BUFX4 BUFX4_10 ( .A(_1100__bF_buf0), .Y(_1100__bF_buf9_bF_buf2) );
BUFX4 BUFX4_11 ( .A(_1100__bF_buf3), .Y(_1100__bF_buf9_bF_buf1) );
BUFX4 BUFX4_12 ( .A(_1100__bF_buf2), .Y(_1100__bF_buf9_bF_buf0) );
BUFX4 BUFX4_13 ( .A(_1101_), .Y(_1101__hier0_bF_buf6) );
BUFX4 BUFX4_14 ( .A(_1101_), .Y(_1101__hier0_bF_buf5) );
BUFX4 BUFX4_15 ( .A(_1101_), .Y(_1101__hier0_bF_buf4) );
BUFX4 BUFX4_16 ( .A(_1101_), .Y(_1101__hier0_bF_buf3) );
BUFX4 BUFX4_17 ( .A(_1101_), .Y(_1101__hier0_bF_buf2) );
BUFX4 BUFX4_18 ( .A(_1101_), .Y(_1101__hier0_bF_buf1) );
BUFX4 BUFX4_19 ( .A(_1101_), .Y(_1101__hier0_bF_buf0) );
BUFX4 BUFX4_20 ( .A(_1039_), .Y(_1039__hier0_bF_buf6) );
BUFX4 BUFX4_21 ( .A(_1039_), .Y(_1039__hier0_bF_buf5) );
BUFX4 BUFX4_22 ( .A(_1039_), .Y(_1039__hier0_bF_buf4) );
BUFX4 BUFX4_23 ( .A(_1039_), .Y(_1039__hier0_bF_buf3) );
BUFX4 BUFX4_24 ( .A(_1039_), .Y(_1039__hier0_bF_buf2) );
BUFX4 BUFX4_25 ( .A(_1039_), .Y(_1039__hier0_bF_buf1) );
BUFX4 BUFX4_26 ( .A(_1039_), .Y(_1039__hier0_bF_buf0) );
BUFX4 BUFX4_27 ( .A(_1135__bF_buf8), .Y(_1135__bF_buf1_bF_buf3) );
BUFX4 BUFX4_28 ( .A(_1135__bF_buf6), .Y(_1135__bF_buf1_bF_buf2) );
BUFX4 BUFX4_29 ( .A(_1135__bF_buf0), .Y(_1135__bF_buf1_bF_buf1) );
BUFX4 BUFX4_30 ( .A(_1135__bF_buf0), .Y(_1135__bF_buf1_bF_buf0) );
BUFX4 BUFX4_31 ( .A(_1135__bF_buf8), .Y(_1135__bF_buf2_bF_buf3) );
BUFX4 BUFX4_32 ( .A(_1135__bF_buf5), .Y(_1135__bF_buf2_bF_buf2) );
BUFX4 BUFX4_33 ( .A(_1135__bF_buf0), .Y(_1135__bF_buf2_bF_buf1) );
BUFX4 BUFX4_34 ( .A(_1135__bF_buf11), .Y(_1135__bF_buf2_bF_buf0) );
BUFX4 BUFX4_35 ( .A(_1135__bF_buf10), .Y(_1135__bF_buf3_bF_buf3) );
BUFX4 BUFX4_36 ( .A(_1135__bF_buf4), .Y(_1135__bF_buf3_bF_buf2) );
BUFX4 BUFX4_37 ( .A(_1135__bF_buf0), .Y(_1135__bF_buf3_bF_buf1) );
BUFX4 BUFX4_38 ( .A(_1135__bF_buf13), .Y(_1135__bF_buf3_bF_buf0) );
BUFX4 BUFX4_39 ( .A(_1135__bF_buf7), .Y(_1135__bF_buf4_bF_buf3) );
BUFX4 BUFX4_40 ( .A(_1135__bF_buf4), .Y(_1135__bF_buf4_bF_buf2) );
BUFX4 BUFX4_41 ( .A(_1135__bF_buf12), .Y(_1135__bF_buf4_bF_buf1) );
BUFX4 BUFX4_42 ( .A(_1135__bF_buf14), .Y(_1135__bF_buf4_bF_buf0) );
BUFX4 BUFX4_43 ( .A(_1135__bF_buf2), .Y(_1135__bF_buf5_bF_buf3) );
BUFX4 BUFX4_44 ( .A(_1135__bF_buf0), .Y(_1135__bF_buf5_bF_buf2) );
BUFX4 BUFX4_45 ( .A(_1135__bF_buf13), .Y(_1135__bF_buf5_bF_buf1) );
BUFX4 BUFX4_46 ( .A(_1135__bF_buf1), .Y(_1135__bF_buf5_bF_buf0) );
BUFX4 BUFX4_47 ( .A(_1135__bF_buf13), .Y(_1135__bF_buf6_bF_buf3) );
BUFX4 BUFX4_48 ( .A(_1135__bF_buf2), .Y(_1135__bF_buf6_bF_buf2) );
BUFX4 BUFX4_49 ( .A(_1135__bF_buf1), .Y(_1135__bF_buf6_bF_buf1) );
BUFX4 BUFX4_50 ( .A(_1135__bF_buf10), .Y(_1135__bF_buf6_bF_buf0) );
BUFX4 BUFX4_51 ( .A(_1135__bF_buf13), .Y(_1135__bF_buf7_bF_buf3) );
BUFX4 BUFX4_52 ( .A(_1135__bF_buf9), .Y(_1135__bF_buf7_bF_buf2) );
BUFX4 BUFX4_53 ( .A(_1135__bF_buf5), .Y(_1135__bF_buf7_bF_buf1) );
BUFX4 BUFX4_54 ( .A(_1135__bF_buf12), .Y(_1135__bF_buf7_bF_buf0) );
BUFX4 BUFX4_55 ( .A(_1135__bF_buf10), .Y(_1135__bF_buf8_bF_buf3) );
BUFX4 BUFX4_56 ( .A(_1135__bF_buf12), .Y(_1135__bF_buf8_bF_buf2) );
BUFX4 BUFX4_57 ( .A(_1135__bF_buf0), .Y(_1135__bF_buf8_bF_buf1) );
BUFX4 BUFX4_58 ( .A(_1135__bF_buf6), .Y(_1135__bF_buf8_bF_buf0) );
BUFX4 BUFX4_59 ( .A(_1135__bF_buf5), .Y(_1135__bF_buf9_bF_buf3) );
BUFX4 BUFX4_60 ( .A(_1135__bF_buf11), .Y(_1135__bF_buf9_bF_buf2) );
BUFX4 BUFX4_61 ( .A(_1135__bF_buf0), .Y(_1135__bF_buf9_bF_buf1) );
BUFX4 BUFX4_62 ( .A(_1135__bF_buf0), .Y(_1135__bF_buf9_bF_buf0) );
BUFX4 BUFX4_63 ( .A(_1135__bF_buf0), .Y(_1135__bF_buf10_bF_buf3) );
BUFX4 BUFX4_64 ( .A(_1135__bF_buf2), .Y(_1135__bF_buf10_bF_buf2) );
BUFX4 BUFX4_65 ( .A(_1135__bF_buf0), .Y(_1135__bF_buf10_bF_buf1) );
BUFX4 BUFX4_66 ( .A(_1135__bF_buf7), .Y(_1135__bF_buf10_bF_buf0) );
BUFX4 BUFX4_67 ( .A(_1135__bF_buf4), .Y(_1135__bF_buf11_bF_buf3) );
BUFX4 BUFX4_68 ( .A(_1135__bF_buf6), .Y(_1135__bF_buf11_bF_buf2) );
BUFX4 BUFX4_69 ( .A(_1135__bF_buf9), .Y(_1135__bF_buf11_bF_buf1) );
BUFX4 BUFX4_70 ( .A(_1135__bF_buf14), .Y(_1135__bF_buf11_bF_buf0) );
BUFX4 BUFX4_71 ( .A(_1135__bF_buf12), .Y(_1135__bF_buf12_bF_buf3) );
BUFX4 BUFX4_72 ( .A(_1135__bF_buf9), .Y(_1135__bF_buf12_bF_buf2) );
BUFX4 BUFX4_73 ( .A(_1135__bF_buf6), .Y(_1135__bF_buf12_bF_buf1) );
BUFX4 BUFX4_74 ( .A(_1135__bF_buf0), .Y(_1135__bF_buf12_bF_buf0) );
BUFX4 BUFX4_75 ( .A(_1135__bF_buf14), .Y(_1135__bF_buf13_bF_buf3) );
BUFX4 BUFX4_76 ( .A(_1135__bF_buf0), .Y(_1135__bF_buf13_bF_buf2) );
BUFX4 BUFX4_77 ( .A(_1135__bF_buf0), .Y(_1135__bF_buf13_bF_buf1) );
BUFX4 BUFX4_78 ( .A(_1135__bF_buf3), .Y(_1135__bF_buf13_bF_buf0) );
BUFX4 BUFX4_79 ( .A(_1135__bF_buf8), .Y(_1135__bF_buf14_bF_buf3) );
BUFX4 BUFX4_80 ( .A(_1135__bF_buf3), .Y(_1135__bF_buf14_bF_buf2) );
BUFX4 BUFX4_81 ( .A(_1135__bF_buf1), .Y(_1135__bF_buf14_bF_buf1) );
BUFX4 BUFX4_82 ( .A(_1135__bF_buf0), .Y(_1135__bF_buf14_bF_buf0) );
BUFX4 BUFX4_83 ( .A(clock_i), .Y(clock_i_hier0_bF_buf9) );
BUFX4 BUFX4_84 ( .A(clock_i), .Y(clock_i_hier0_bF_buf8) );
BUFX4 BUFX4_85 ( .A(clock_i), .Y(clock_i_hier0_bF_buf7) );
BUFX4 BUFX4_86 ( .A(clock_i), .Y(clock_i_hier0_bF_buf6) );
BUFX4 BUFX4_87 ( .A(clock_i), .Y(clock_i_hier0_bF_buf5) );
BUFX4 BUFX4_88 ( .A(clock_i), .Y(clock_i_hier0_bF_buf4) );
BUFX4 BUFX4_89 ( .A(clock_i), .Y(clock_i_hier0_bF_buf3) );
BUFX4 BUFX4_90 ( .A(clock_i), .Y(clock_i_hier0_bF_buf2) );
BUFX4 BUFX4_91 ( .A(clock_i), .Y(clock_i_hier0_bF_buf1) );
BUFX4 BUFX4_92 ( .A(clock_i), .Y(clock_i_hier0_bF_buf0) );
BUFX4 BUFX4_93 ( .A(_1100__bF_buf8), .Y(_1100__bF_buf10_bF_buf3) );
BUFX4 BUFX4_94 ( .A(_1100__bF_buf10), .Y(_1100__bF_buf10_bF_buf2) );
BUFX4 BUFX4_95 ( .A(_1100__bF_buf7), .Y(_1100__bF_buf10_bF_buf1) );
BUFX4 BUFX4_96 ( .A(_1100__bF_buf2), .Y(_1100__bF_buf10_bF_buf0) );
BUFX4 BUFX4_97 ( .A(_1100__bF_buf5), .Y(_1100__bF_buf11_bF_buf3) );
BUFX4 BUFX4_98 ( .A(_1100__bF_buf4), .Y(_1100__bF_buf11_bF_buf2) );
BUFX4 BUFX4_99 ( .A(_1100__bF_buf1), .Y(_1100__bF_buf11_bF_buf1) );
BUFX4 BUFX4_100 ( .A(_1100__bF_buf4), .Y(_1100__bF_buf11_bF_buf0) );
BUFX4 BUFX4_101 ( .A(_1100__bF_buf10), .Y(_1100__bF_buf12_bF_buf3) );
BUFX4 BUFX4_102 ( .A(_1100__bF_buf6), .Y(_1100__bF_buf12_bF_buf2) );
BUFX4 BUFX4_103 ( .A(_1100__bF_buf3), .Y(_1100__bF_buf12_bF_buf1) );
BUFX4 BUFX4_104 ( .A(_1100__bF_buf7), .Y(_1100__bF_buf12_bF_buf0) );
BUFX4 BUFX4_105 ( .A(_1100__bF_buf2), .Y(_1100__bF_buf13_bF_buf3) );
BUFX4 BUFX4_106 ( .A(_1100__bF_buf5), .Y(_1100__bF_buf13_bF_buf2) );
BUFX4 BUFX4_107 ( .A(_1100__bF_buf4), .Y(_1100__bF_buf13_bF_buf1) );
BUFX4 BUFX4_108 ( .A(_1100__bF_buf0), .Y(_1100__bF_buf13_bF_buf0) );
BUFX4 BUFX4_109 ( .A(_1100__bF_buf7), .Y(_1100__bF_buf14_bF_buf3) );
BUFX4 BUFX4_110 ( .A(_1100__bF_buf0), .Y(_1100__bF_buf14_bF_buf2) );
BUFX4 BUFX4_111 ( .A(_1100__bF_buf2), .Y(_1100__bF_buf14_bF_buf1) );
BUFX4 BUFX4_112 ( .A(_1100__bF_buf8), .Y(_1100__bF_buf14_bF_buf0) );
BUFX4 BUFX4_113 ( .A(_1031_), .Y(_1031__hier0_bF_buf7) );
BUFX4 BUFX4_114 ( .A(_1031_), .Y(_1031__hier0_bF_buf6) );
BUFX4 BUFX4_115 ( .A(_1031_), .Y(_1031__hier0_bF_buf5) );
BUFX4 BUFX4_116 ( .A(_1031_), .Y(_1031__hier0_bF_buf4) );
BUFX4 BUFX4_117 ( .A(_1031_), .Y(_1031__hier0_bF_buf3) );
BUFX4 BUFX4_118 ( .A(_1031_), .Y(_1031__hier0_bF_buf2) );
BUFX4 BUFX4_119 ( .A(_1031_), .Y(_1031__hier0_bF_buf1) );
BUFX4 BUFX4_120 ( .A(_1031_), .Y(_1031__hier0_bF_buf0) );
BUFX4 BUFX4_121 ( .A(_1101__hier0_bF_buf5), .Y(_1101__bF_buf58) );
BUFX4 BUFX4_122 ( .A(_1101__hier0_bF_buf6), .Y(_1101__bF_buf57) );
BUFX4 BUFX4_123 ( .A(_1101__hier0_bF_buf5), .Y(_1101__bF_buf56) );
BUFX4 BUFX4_124 ( .A(_1101__hier0_bF_buf3), .Y(_1101__bF_buf55) );
BUFX4 BUFX4_125 ( .A(_1101__hier0_bF_buf1), .Y(_1101__bF_buf54) );
BUFX4 BUFX4_126 ( .A(_1101__hier0_bF_buf1), .Y(_1101__bF_buf53) );
BUFX4 BUFX4_127 ( .A(_1101__hier0_bF_buf0), .Y(_1101__bF_buf52) );
BUFX4 BUFX4_128 ( .A(_1101__hier0_bF_buf5), .Y(_1101__bF_buf51) );
BUFX4 BUFX4_129 ( .A(_1101__hier0_bF_buf4), .Y(_1101__bF_buf50) );
BUFX4 BUFX4_130 ( .A(_1101__hier0_bF_buf0), .Y(_1101__bF_buf49) );
BUFX4 BUFX4_131 ( .A(_1101__hier0_bF_buf6), .Y(_1101__bF_buf48) );
BUFX4 BUFX4_132 ( .A(_1101__hier0_bF_buf1), .Y(_1101__bF_buf47) );
BUFX4 BUFX4_133 ( .A(_1101__hier0_bF_buf0), .Y(_1101__bF_buf46) );
BUFX4 BUFX4_134 ( .A(_1101__hier0_bF_buf6), .Y(_1101__bF_buf45) );
BUFX4 BUFX4_135 ( .A(_1101__hier0_bF_buf6), .Y(_1101__bF_buf44) );
BUFX4 BUFX4_136 ( .A(_1101__hier0_bF_buf1), .Y(_1101__bF_buf43) );
BUFX4 BUFX4_137 ( .A(_1101__hier0_bF_buf5), .Y(_1101__bF_buf42) );
BUFX4 BUFX4_138 ( .A(_1101__hier0_bF_buf4), .Y(_1101__bF_buf41) );
BUFX4 BUFX4_139 ( .A(_1101__hier0_bF_buf3), .Y(_1101__bF_buf40) );
BUFX4 BUFX4_140 ( .A(_1101__hier0_bF_buf5), .Y(_1101__bF_buf39) );
BUFX4 BUFX4_141 ( .A(_1101__hier0_bF_buf3), .Y(_1101__bF_buf38) );
BUFX4 BUFX4_142 ( .A(_1101__hier0_bF_buf2), .Y(_1101__bF_buf37) );
BUFX4 BUFX4_143 ( .A(_1101__hier0_bF_buf1), .Y(_1101__bF_buf36) );
BUFX4 BUFX4_144 ( .A(_1101__hier0_bF_buf3), .Y(_1101__bF_buf35) );
BUFX4 BUFX4_145 ( .A(_1101__hier0_bF_buf1), .Y(_1101__bF_buf34) );
BUFX4 BUFX4_146 ( .A(_1101__hier0_bF_buf2), .Y(_1101__bF_buf33) );
BUFX4 BUFX4_147 ( .A(_1101__hier0_bF_buf0), .Y(_1101__bF_buf32) );
BUFX4 BUFX4_148 ( .A(_1101__hier0_bF_buf4), .Y(_1101__bF_buf31) );
BUFX4 BUFX4_149 ( .A(_1101__hier0_bF_buf0), .Y(_1101__bF_buf30) );
BUFX4 BUFX4_150 ( .A(_1101__hier0_bF_buf2), .Y(_1101__bF_buf29) );
BUFX4 BUFX4_151 ( .A(_1101__hier0_bF_buf1), .Y(_1101__bF_buf28) );
BUFX4 BUFX4_152 ( .A(_1101__hier0_bF_buf3), .Y(_1101__bF_buf27) );
BUFX4 BUFX4_153 ( .A(_1101__hier0_bF_buf6), .Y(_1101__bF_buf26) );
BUFX4 BUFX4_154 ( .A(_1101__hier0_bF_buf3), .Y(_1101__bF_buf25) );
BUFX4 BUFX4_155 ( .A(_1101__hier0_bF_buf2), .Y(_1101__bF_buf24) );
BUFX4 BUFX4_156 ( .A(_1101__hier0_bF_buf2), .Y(_1101__bF_buf23) );
BUFX4 BUFX4_157 ( .A(_1101__hier0_bF_buf4), .Y(_1101__bF_buf22) );
BUFX4 BUFX4_158 ( .A(_1101__hier0_bF_buf3), .Y(_1101__bF_buf21) );
BUFX4 BUFX4_159 ( .A(_1101__hier0_bF_buf4), .Y(_1101__bF_buf20) );
BUFX4 BUFX4_160 ( .A(_1101__hier0_bF_buf4), .Y(_1101__bF_buf19) );
BUFX4 BUFX4_161 ( .A(_1101__hier0_bF_buf2), .Y(_1101__bF_buf18) );
BUFX4 BUFX4_162 ( .A(_1101__hier0_bF_buf5), .Y(_1101__bF_buf17) );
BUFX4 BUFX4_163 ( .A(_1101__hier0_bF_buf6), .Y(_1101__bF_buf16) );
BUFX4 BUFX4_164 ( .A(_1101__hier0_bF_buf0), .Y(_1101__bF_buf15) );
BUFX4 BUFX4_165 ( .A(_1101__hier0_bF_buf5), .Y(_1101__bF_buf14) );
BUFX4 BUFX4_166 ( .A(_1101__hier0_bF_buf4), .Y(_1101__bF_buf13) );
BUFX4 BUFX4_167 ( .A(_1101__hier0_bF_buf6), .Y(_1101__bF_buf12) );
BUFX4 BUFX4_168 ( .A(_1101__hier0_bF_buf0), .Y(_1101__bF_buf11) );
BUFX4 BUFX4_169 ( .A(_1101__hier0_bF_buf3), .Y(_1101__bF_buf10) );
BUFX4 BUFX4_170 ( .A(_1101__hier0_bF_buf5), .Y(_1101__bF_buf9) );
BUFX4 BUFX4_171 ( .A(_1101__hier0_bF_buf2), .Y(_1101__bF_buf8) );
BUFX4 BUFX4_172 ( .A(_1101__hier0_bF_buf5), .Y(_1101__bF_buf7) );
BUFX4 BUFX4_173 ( .A(_1101__hier0_bF_buf6), .Y(_1101__bF_buf6) );
BUFX4 BUFX4_174 ( .A(_1101__hier0_bF_buf4), .Y(_1101__bF_buf5) );
BUFX4 BUFX4_175 ( .A(_1101__hier0_bF_buf0), .Y(_1101__bF_buf4) );
BUFX4 BUFX4_176 ( .A(_1101__hier0_bF_buf6), .Y(_1101__bF_buf3) );
BUFX4 BUFX4_177 ( .A(_1101__hier0_bF_buf2), .Y(_1101__bF_buf2) );
BUFX4 BUFX4_178 ( .A(_1101__hier0_bF_buf4), .Y(_1101__bF_buf1) );
BUFX4 BUFX4_179 ( .A(_1101__hier0_bF_buf1), .Y(_1101__bF_buf0) );
BUFX4 BUFX4_180 ( .A(_1039__hier0_bF_buf2), .Y(_1039__bF_buf57) );
BUFX4 BUFX4_181 ( .A(_1039__hier0_bF_buf6), .Y(_1039__bF_buf56) );
BUFX4 BUFX4_182 ( .A(_1039__hier0_bF_buf6), .Y(_1039__bF_buf55) );
BUFX4 BUFX4_183 ( .A(_1039__hier0_bF_buf2), .Y(_1039__bF_buf54) );
BUFX4 BUFX4_184 ( .A(_1039__hier0_bF_buf2), .Y(_1039__bF_buf53) );
BUFX4 BUFX4_185 ( .A(_1039__hier0_bF_buf5), .Y(_1039__bF_buf52) );
BUFX4 BUFX4_186 ( .A(_1039__hier0_bF_buf0), .Y(_1039__bF_buf51) );
BUFX4 BUFX4_187 ( .A(_1039__hier0_bF_buf5), .Y(_1039__bF_buf50) );
BUFX4 BUFX4_188 ( .A(_1039__hier0_bF_buf5), .Y(_1039__bF_buf49) );
BUFX4 BUFX4_189 ( .A(_1039__hier0_bF_buf5), .Y(_1039__bF_buf48) );
BUFX4 BUFX4_190 ( .A(_1039__hier0_bF_buf4), .Y(_1039__bF_buf47) );
BUFX4 BUFX4_191 ( .A(_1039__hier0_bF_buf0), .Y(_1039__bF_buf46) );
BUFX4 BUFX4_192 ( .A(_1039__hier0_bF_buf0), .Y(_1039__bF_buf45) );
BUFX4 BUFX4_193 ( .A(_1039__hier0_bF_buf3), .Y(_1039__bF_buf44) );
BUFX4 BUFX4_194 ( .A(_1039__hier0_bF_buf4), .Y(_1039__bF_buf43) );
BUFX4 BUFX4_195 ( .A(_1039__hier0_bF_buf3), .Y(_1039__bF_buf42) );
BUFX4 BUFX4_196 ( .A(_1039__hier0_bF_buf5), .Y(_1039__bF_buf41) );
BUFX4 BUFX4_197 ( .A(_1039__hier0_bF_buf2), .Y(_1039__bF_buf40) );
BUFX4 BUFX4_198 ( .A(_1039__hier0_bF_buf1), .Y(_1039__bF_buf39) );
BUFX4 BUFX4_199 ( .A(_1039__hier0_bF_buf6), .Y(_1039__bF_buf38) );
BUFX4 BUFX4_200 ( .A(_1039__hier0_bF_buf1), .Y(_1039__bF_buf37) );
BUFX4 BUFX4_201 ( .A(_1039__hier0_bF_buf5), .Y(_1039__bF_buf36) );
BUFX4 BUFX4_202 ( .A(_1039__hier0_bF_buf0), .Y(_1039__bF_buf35) );
BUFX4 BUFX4_203 ( .A(_1039__hier0_bF_buf3), .Y(_1039__bF_buf34) );
BUFX4 BUFX4_204 ( .A(_1039__hier0_bF_buf1), .Y(_1039__bF_buf33) );
BUFX4 BUFX4_205 ( .A(_1039__hier0_bF_buf3), .Y(_1039__bF_buf32) );
BUFX4 BUFX4_206 ( .A(_1039__hier0_bF_buf5), .Y(_1039__bF_buf31) );
BUFX4 BUFX4_207 ( .A(_1039__hier0_bF_buf0), .Y(_1039__bF_buf30) );
BUFX4 BUFX4_208 ( .A(_1039__hier0_bF_buf2), .Y(_1039__bF_buf29) );
BUFX4 BUFX4_209 ( .A(_1039__hier0_bF_buf4), .Y(_1039__bF_buf28) );
BUFX4 BUFX4_210 ( .A(_1039__hier0_bF_buf1), .Y(_1039__bF_buf27) );
BUFX4 BUFX4_211 ( .A(_1039__hier0_bF_buf2), .Y(_1039__bF_buf26) );
BUFX4 BUFX4_212 ( .A(_1039__hier0_bF_buf5), .Y(_1039__bF_buf25) );
BUFX4 BUFX4_213 ( .A(_1039__hier0_bF_buf1), .Y(_1039__bF_buf24) );
BUFX4 BUFX4_214 ( .A(_1039__hier0_bF_buf4), .Y(_1039__bF_buf23) );
BUFX4 BUFX4_215 ( .A(_1039__hier0_bF_buf6), .Y(_1039__bF_buf22) );
BUFX4 BUFX4_216 ( .A(_1039__hier0_bF_buf2), .Y(_1039__bF_buf21) );
BUFX4 BUFX4_217 ( .A(_1039__hier0_bF_buf6), .Y(_1039__bF_buf20) );
BUFX4 BUFX4_218 ( .A(_1039__hier0_bF_buf3), .Y(_1039__bF_buf19) );
BUFX4 BUFX4_219 ( .A(_1039__hier0_bF_buf3), .Y(_1039__bF_buf18) );
BUFX4 BUFX4_220 ( .A(_1039__hier0_bF_buf0), .Y(_1039__bF_buf17) );
BUFX4 BUFX4_221 ( .A(_1039__hier0_bF_buf1), .Y(_1039__bF_buf16) );
BUFX4 BUFX4_222 ( .A(_1039__hier0_bF_buf6), .Y(_1039__bF_buf15) );
BUFX4 BUFX4_223 ( .A(_1039__hier0_bF_buf4), .Y(_1039__bF_buf14) );
BUFX4 BUFX4_224 ( .A(_1039__hier0_bF_buf4), .Y(_1039__bF_buf13) );
BUFX4 BUFX4_225 ( .A(_1039__hier0_bF_buf6), .Y(_1039__bF_buf12) );
BUFX4 BUFX4_226 ( .A(_1039__hier0_bF_buf5), .Y(_1039__bF_buf11) );
BUFX4 BUFX4_227 ( .A(_1039__hier0_bF_buf3), .Y(_1039__bF_buf10) );
BUFX4 BUFX4_228 ( .A(_1039__hier0_bF_buf0), .Y(_1039__bF_buf9) );
BUFX4 BUFX4_229 ( .A(_1039__hier0_bF_buf0), .Y(_1039__bF_buf8) );
BUFX4 BUFX4_230 ( .A(_1039__hier0_bF_buf2), .Y(_1039__bF_buf7) );
BUFX4 BUFX4_231 ( .A(_1039__hier0_bF_buf1), .Y(_1039__bF_buf6) );
BUFX4 BUFX4_232 ( .A(_1039__hier0_bF_buf6), .Y(_1039__bF_buf5) );
BUFX4 BUFX4_233 ( .A(_1039__hier0_bF_buf4), .Y(_1039__bF_buf4) );
BUFX4 BUFX4_234 ( .A(_1039__hier0_bF_buf3), .Y(_1039__bF_buf3) );
BUFX4 BUFX4_235 ( .A(_1039__hier0_bF_buf1), .Y(_1039__bF_buf2) );
BUFX4 BUFX4_236 ( .A(_1039__hier0_bF_buf4), .Y(_1039__bF_buf1) );
BUFX4 BUFX4_237 ( .A(_1039__hier0_bF_buf6), .Y(_1039__bF_buf0) );
BUFX4 BUFX4_238 ( .A(_611_), .Y(_611__bF_buf7) );
BUFX4 BUFX4_239 ( .A(_611_), .Y(_611__bF_buf6) );
BUFX4 BUFX4_240 ( .A(_611_), .Y(_611__bF_buf5) );
BUFX4 BUFX4_241 ( .A(_611_), .Y(_611__bF_buf4) );
BUFX4 BUFX4_242 ( .A(_611_), .Y(_611__bF_buf3) );
BUFX4 BUFX4_243 ( .A(_611_), .Y(_611__bF_buf2) );
BUFX4 BUFX4_244 ( .A(_611_), .Y(_611__bF_buf1) );
BUFX4 BUFX4_245 ( .A(_611_), .Y(_611__bF_buf0) );
BUFX4 BUFX4_246 ( .A(_1100_), .Y(_1100__bF_buf14) );
BUFX4 BUFX4_247 ( .A(_1100_), .Y(_1100__bF_buf13) );
BUFX4 BUFX4_248 ( .A(_1100_), .Y(_1100__bF_buf12) );
BUFX4 BUFX4_249 ( .A(_1100_), .Y(_1100__bF_buf11) );
BUFX4 BUFX4_250 ( .A(_1100_), .Y(_1100__bF_buf10) );
BUFX4 BUFX4_251 ( .A(_1100_), .Y(_1100__bF_buf9) );
BUFX4 BUFX4_252 ( .A(_1100_), .Y(_1100__bF_buf8) );
BUFX4 BUFX4_253 ( .A(_1100_), .Y(_1100__bF_buf7) );
BUFX4 BUFX4_254 ( .A(_1100_), .Y(_1100__bF_buf6) );
BUFX4 BUFX4_255 ( .A(_1100_), .Y(_1100__bF_buf5) );
BUFX4 BUFX4_256 ( .A(_1100_), .Y(_1100__bF_buf4) );
BUFX4 BUFX4_257 ( .A(_1100_), .Y(_1100__bF_buf3) );
BUFX4 BUFX4_258 ( .A(_1100_), .Y(_1100__bF_buf2) );
BUFX4 BUFX4_259 ( .A(_1100_), .Y(_1100__bF_buf1) );
BUFX4 BUFX4_260 ( .A(_1100_), .Y(_1100__bF_buf0) );
BUFX4 BUFX4_261 ( .A(enable_i), .Y(enable_i_bF_buf7) );
BUFX4 BUFX4_262 ( .A(enable_i), .Y(enable_i_bF_buf6) );
BUFX4 BUFX4_263 ( .A(enable_i), .Y(enable_i_bF_buf5) );
BUFX4 BUFX4_264 ( .A(enable_i), .Y(enable_i_bF_buf4) );
BUFX4 BUFX4_265 ( .A(enable_i), .Y(enable_i_bF_buf3) );
BUFX4 BUFX4_266 ( .A(enable_i), .Y(enable_i_bF_buf2) );
BUFX4 BUFX4_267 ( .A(enable_i), .Y(enable_i_bF_buf1) );
BUFX4 BUFX4_268 ( .A(enable_i), .Y(enable_i_bF_buf0) );
BUFX4 BUFX4_269 ( .A(_1135_), .Y(_1135__bF_buf14) );
BUFX4 BUFX4_270 ( .A(_1135_), .Y(_1135__bF_buf13) );
BUFX4 BUFX4_271 ( .A(_1135_), .Y(_1135__bF_buf12) );
BUFX4 BUFX4_272 ( .A(_1135_), .Y(_1135__bF_buf11) );
BUFX4 BUFX4_273 ( .A(_1135_), .Y(_1135__bF_buf10) );
BUFX4 BUFX4_274 ( .A(_1135_), .Y(_1135__bF_buf9) );
BUFX4 BUFX4_275 ( .A(_1135_), .Y(_1135__bF_buf8) );
BUFX4 BUFX4_276 ( .A(_1135_), .Y(_1135__bF_buf7) );
BUFX4 BUFX4_277 ( .A(_1135_), .Y(_1135__bF_buf6) );
BUFX4 BUFX4_278 ( .A(_1135_), .Y(_1135__bF_buf5) );
BUFX4 BUFX4_279 ( .A(_1135_), .Y(_1135__bF_buf4) );
BUFX4 BUFX4_280 ( .A(_1135_), .Y(_1135__bF_buf3) );
BUFX4 BUFX4_281 ( .A(_1135_), .Y(_1135__bF_buf2) );
BUFX4 BUFX4_282 ( .A(_1135_), .Y(_1135__bF_buf1) );
BUFX4 BUFX4_283 ( .A(_1135_), .Y(_1135__bF_buf0) );
CLKBUF1 CLKBUF1_1 ( .A(clock_i_hier0_bF_buf1), .Y(clock_i_bF_buf101) );
CLKBUF1 CLKBUF1_2 ( .A(clock_i_hier0_bF_buf4), .Y(clock_i_bF_buf100) );
CLKBUF1 CLKBUF1_3 ( .A(clock_i_hier0_bF_buf6), .Y(clock_i_bF_buf99) );
CLKBUF1 CLKBUF1_4 ( .A(clock_i_hier0_bF_buf9), .Y(clock_i_bF_buf98) );
CLKBUF1 CLKBUF1_5 ( .A(clock_i_hier0_bF_buf7), .Y(clock_i_bF_buf97) );
CLKBUF1 CLKBUF1_6 ( .A(clock_i_hier0_bF_buf8), .Y(clock_i_bF_buf96) );
CLKBUF1 CLKBUF1_7 ( .A(clock_i_hier0_bF_buf6), .Y(clock_i_bF_buf95) );
CLKBUF1 CLKBUF1_8 ( .A(clock_i_hier0_bF_buf5), .Y(clock_i_bF_buf94) );
CLKBUF1 CLKBUF1_9 ( .A(clock_i_hier0_bF_buf8), .Y(clock_i_bF_buf93) );
CLKBUF1 CLKBUF1_10 ( .A(clock_i_hier0_bF_buf2), .Y(clock_i_bF_buf92) );
CLKBUF1 CLKBUF1_11 ( .A(clock_i_hier0_bF_buf8), .Y(clock_i_bF_buf91) );
CLKBUF1 CLKBUF1_12 ( .A(clock_i_hier0_bF_buf7), .Y(clock_i_bF_buf90) );
CLKBUF1 CLKBUF1_13 ( .A(clock_i_hier0_bF_buf2), .Y(clock_i_bF_buf89) );
CLKBUF1 CLKBUF1_14 ( .A(clock_i_hier0_bF_buf0), .Y(clock_i_bF_buf88) );
CLKBUF1 CLKBUF1_15 ( .A(clock_i_hier0_bF_buf4), .Y(clock_i_bF_buf87) );
CLKBUF1 CLKBUF1_16 ( .A(clock_i_hier0_bF_buf6), .Y(clock_i_bF_buf86) );
CLKBUF1 CLKBUF1_17 ( .A(clock_i_hier0_bF_buf5), .Y(clock_i_bF_buf85) );
CLKBUF1 CLKBUF1_18 ( .A(clock_i_hier0_bF_buf1), .Y(clock_i_bF_buf84) );
CLKBUF1 CLKBUF1_19 ( .A(clock_i_hier0_bF_buf1), .Y(clock_i_bF_buf83) );
CLKBUF1 CLKBUF1_20 ( .A(clock_i_hier0_bF_buf3), .Y(clock_i_bF_buf82) );
CLKBUF1 CLKBUF1_21 ( .A(clock_i_hier0_bF_buf0), .Y(clock_i_bF_buf81) );
CLKBUF1 CLKBUF1_22 ( .A(clock_i_hier0_bF_buf9), .Y(clock_i_bF_buf80) );
CLKBUF1 CLKBUF1_23 ( .A(clock_i_hier0_bF_buf1), .Y(clock_i_bF_buf79) );
CLKBUF1 CLKBUF1_24 ( .A(clock_i_hier0_bF_buf8), .Y(clock_i_bF_buf78) );
CLKBUF1 CLKBUF1_25 ( .A(clock_i_hier0_bF_buf5), .Y(clock_i_bF_buf77) );
CLKBUF1 CLKBUF1_26 ( .A(clock_i_hier0_bF_buf5), .Y(clock_i_bF_buf76) );
CLKBUF1 CLKBUF1_27 ( .A(clock_i_hier0_bF_buf0), .Y(clock_i_bF_buf75) );
CLKBUF1 CLKBUF1_28 ( .A(clock_i_hier0_bF_buf4), .Y(clock_i_bF_buf74) );
CLKBUF1 CLKBUF1_29 ( .A(clock_i_hier0_bF_buf8), .Y(clock_i_bF_buf73) );
CLKBUF1 CLKBUF1_30 ( .A(clock_i_hier0_bF_buf5), .Y(clock_i_bF_buf72) );
CLKBUF1 CLKBUF1_31 ( .A(clock_i_hier0_bF_buf7), .Y(clock_i_bF_buf71) );
CLKBUF1 CLKBUF1_32 ( .A(clock_i_hier0_bF_buf5), .Y(clock_i_bF_buf70) );
CLKBUF1 CLKBUF1_33 ( .A(clock_i_hier0_bF_buf1), .Y(clock_i_bF_buf69) );
CLKBUF1 CLKBUF1_34 ( .A(clock_i_hier0_bF_buf4), .Y(clock_i_bF_buf68) );
CLKBUF1 CLKBUF1_35 ( .A(clock_i_hier0_bF_buf6), .Y(clock_i_bF_buf67) );
CLKBUF1 CLKBUF1_36 ( .A(clock_i_hier0_bF_buf0), .Y(clock_i_bF_buf66) );
CLKBUF1 CLKBUF1_37 ( .A(clock_i_hier0_bF_buf3), .Y(clock_i_bF_buf65) );
CLKBUF1 CLKBUF1_38 ( .A(clock_i_hier0_bF_buf3), .Y(clock_i_bF_buf64) );
CLKBUF1 CLKBUF1_39 ( .A(clock_i_hier0_bF_buf7), .Y(clock_i_bF_buf63) );
CLKBUF1 CLKBUF1_40 ( .A(clock_i_hier0_bF_buf3), .Y(clock_i_bF_buf62) );
CLKBUF1 CLKBUF1_41 ( .A(clock_i_hier0_bF_buf2), .Y(clock_i_bF_buf61) );
CLKBUF1 CLKBUF1_42 ( .A(clock_i_hier0_bF_buf5), .Y(clock_i_bF_buf60) );
CLKBUF1 CLKBUF1_43 ( .A(clock_i_hier0_bF_buf6), .Y(clock_i_bF_buf59) );
CLKBUF1 CLKBUF1_44 ( .A(clock_i_hier0_bF_buf8), .Y(clock_i_bF_buf58) );
CLKBUF1 CLKBUF1_45 ( .A(clock_i_hier0_bF_buf9), .Y(clock_i_bF_buf57) );
CLKBUF1 CLKBUF1_46 ( .A(clock_i_hier0_bF_buf2), .Y(clock_i_bF_buf56) );
CLKBUF1 CLKBUF1_47 ( .A(clock_i_hier0_bF_buf6), .Y(clock_i_bF_buf55) );
CLKBUF1 CLKBUF1_48 ( .A(clock_i_hier0_bF_buf8), .Y(clock_i_bF_buf54) );
CLKBUF1 CLKBUF1_49 ( .A(clock_i_hier0_bF_buf0), .Y(clock_i_bF_buf53) );
CLKBUF1 CLKBUF1_50 ( .A(clock_i_hier0_bF_buf1), .Y(clock_i_bF_buf52) );
CLKBUF1 CLKBUF1_51 ( .A(clock_i_hier0_bF_buf4), .Y(clock_i_bF_buf51) );
CLKBUF1 CLKBUF1_52 ( .A(clock_i_hier0_bF_buf4), .Y(clock_i_bF_buf50) );
CLKBUF1 CLKBUF1_53 ( .A(clock_i_hier0_bF_buf4), .Y(clock_i_bF_buf49) );
CLKBUF1 CLKBUF1_54 ( .A(clock_i_hier0_bF_buf2), .Y(clock_i_bF_buf48) );
CLKBUF1 CLKBUF1_55 ( .A(clock_i_hier0_bF_buf6), .Y(clock_i_bF_buf47) );
CLKBUF1 CLKBUF1_56 ( .A(clock_i_hier0_bF_buf2), .Y(clock_i_bF_buf46) );
CLKBUF1 CLKBUF1_57 ( .A(clock_i_hier0_bF_buf0), .Y(clock_i_bF_buf45) );
CLKBUF1 CLKBUF1_58 ( .A(clock_i_hier0_bF_buf3), .Y(clock_i_bF_buf44) );
CLKBUF1 CLKBUF1_59 ( .A(clock_i_hier0_bF_buf1), .Y(clock_i_bF_buf43) );
CLKBUF1 CLKBUF1_60 ( .A(clock_i_hier0_bF_buf6), .Y(clock_i_bF_buf42) );
CLKBUF1 CLKBUF1_61 ( .A(clock_i_hier0_bF_buf9), .Y(clock_i_bF_buf41) );
CLKBUF1 CLKBUF1_62 ( .A(clock_i_hier0_bF_buf4), .Y(clock_i_bF_buf40) );
CLKBUF1 CLKBUF1_63 ( .A(clock_i_hier0_bF_buf1), .Y(clock_i_bF_buf39) );
CLKBUF1 CLKBUF1_64 ( .A(clock_i_hier0_bF_buf9), .Y(clock_i_bF_buf38) );
CLKBUF1 CLKBUF1_65 ( .A(clock_i_hier0_bF_buf8), .Y(clock_i_bF_buf37) );
CLKBUF1 CLKBUF1_66 ( .A(clock_i_hier0_bF_buf2), .Y(clock_i_bF_buf36) );
CLKBUF1 CLKBUF1_67 ( .A(clock_i_hier0_bF_buf5), .Y(clock_i_bF_buf35) );
CLKBUF1 CLKBUF1_68 ( .A(clock_i_hier0_bF_buf0), .Y(clock_i_bF_buf34) );
CLKBUF1 CLKBUF1_69 ( .A(clock_i_hier0_bF_buf3), .Y(clock_i_bF_buf33) );
CLKBUF1 CLKBUF1_70 ( .A(clock_i_hier0_bF_buf8), .Y(clock_i_bF_buf32) );
CLKBUF1 CLKBUF1_71 ( .A(clock_i_hier0_bF_buf3), .Y(clock_i_bF_buf31) );
CLKBUF1 CLKBUF1_72 ( .A(clock_i_hier0_bF_buf7), .Y(clock_i_bF_buf30) );
CLKBUF1 CLKBUF1_73 ( .A(clock_i_hier0_bF_buf9), .Y(clock_i_bF_buf29) );
CLKBUF1 CLKBUF1_74 ( .A(clock_i_hier0_bF_buf7), .Y(clock_i_bF_buf28) );
CLKBUF1 CLKBUF1_75 ( .A(clock_i_hier0_bF_buf2), .Y(clock_i_bF_buf27) );
CLKBUF1 CLKBUF1_76 ( .A(clock_i_hier0_bF_buf3), .Y(clock_i_bF_buf26) );
CLKBUF1 CLKBUF1_77 ( .A(clock_i_hier0_bF_buf4), .Y(clock_i_bF_buf25) );
CLKBUF1 CLKBUF1_78 ( .A(clock_i_hier0_bF_buf9), .Y(clock_i_bF_buf24) );
CLKBUF1 CLKBUF1_79 ( .A(clock_i_hier0_bF_buf8), .Y(clock_i_bF_buf23) );
CLKBUF1 CLKBUF1_80 ( .A(clock_i_hier0_bF_buf9), .Y(clock_i_bF_buf22) );
CLKBUF1 CLKBUF1_81 ( .A(clock_i_hier0_bF_buf3), .Y(clock_i_bF_buf21) );
CLKBUF1 CLKBUF1_82 ( .A(clock_i_hier0_bF_buf3), .Y(clock_i_bF_buf20) );
CLKBUF1 CLKBUF1_83 ( .A(clock_i_hier0_bF_buf6), .Y(clock_i_bF_buf19) );
CLKBUF1 CLKBUF1_84 ( .A(clock_i_hier0_bF_buf9), .Y(clock_i_bF_buf18) );
CLKBUF1 CLKBUF1_85 ( .A(clock_i_hier0_bF_buf4), .Y(clock_i_bF_buf17) );
CLKBUF1 CLKBUF1_86 ( .A(clock_i_hier0_bF_buf0), .Y(clock_i_bF_buf16) );
CLKBUF1 CLKBUF1_87 ( .A(clock_i_hier0_bF_buf9), .Y(clock_i_bF_buf15) );
CLKBUF1 CLKBUF1_88 ( .A(clock_i_hier0_bF_buf1), .Y(clock_i_bF_buf14) );
CLKBUF1 CLKBUF1_89 ( .A(clock_i_hier0_bF_buf0), .Y(clock_i_bF_buf13) );
CLKBUF1 CLKBUF1_90 ( .A(clock_i_hier0_bF_buf2), .Y(clock_i_bF_buf12) );
CLKBUF1 CLKBUF1_91 ( .A(clock_i_hier0_bF_buf9), .Y(clock_i_bF_buf11) );
CLKBUF1 CLKBUF1_92 ( .A(clock_i_hier0_bF_buf8), .Y(clock_i_bF_buf10) );
CLKBUF1 CLKBUF1_93 ( .A(clock_i_hier0_bF_buf6), .Y(clock_i_bF_buf9) );
CLKBUF1 CLKBUF1_94 ( .A(clock_i_hier0_bF_buf2), .Y(clock_i_bF_buf8) );
CLKBUF1 CLKBUF1_95 ( .A(clock_i_hier0_bF_buf0), .Y(clock_i_bF_buf7) );
CLKBUF1 CLKBUF1_96 ( .A(clock_i_hier0_bF_buf7), .Y(clock_i_bF_buf6) );
CLKBUF1 CLKBUF1_97 ( .A(clock_i_hier0_bF_buf5), .Y(clock_i_bF_buf5) );
CLKBUF1 CLKBUF1_98 ( .A(clock_i_hier0_bF_buf7), .Y(clock_i_bF_buf4) );
CLKBUF1 CLKBUF1_99 ( .A(clock_i_hier0_bF_buf5), .Y(clock_i_bF_buf3) );
CLKBUF1 CLKBUF1_100 ( .A(clock_i_hier0_bF_buf7), .Y(clock_i_bF_buf2) );
CLKBUF1 CLKBUF1_101 ( .A(clock_i_hier0_bF_buf7), .Y(clock_i_bF_buf1) );
CLKBUF1 CLKBUF1_102 ( .A(clock_i_hier0_bF_buf1), .Y(clock_i_bF_buf0) );
BUFX4 BUFX4_284 ( .A(_613_), .Y(_613__bF_buf4) );
BUFX4 BUFX4_285 ( .A(_613_), .Y(_613__bF_buf3) );
BUFX4 BUFX4_286 ( .A(_613_), .Y(_613__bF_buf2) );
BUFX4 BUFX4_287 ( .A(_613_), .Y(_613__bF_buf1) );
BUFX4 BUFX4_288 ( .A(_613_), .Y(_613__bF_buf0) );
BUFX4 BUFX4_289 ( .A(_1134_), .Y(_1134__bF_buf14) );
BUFX4 BUFX4_290 ( .A(_1134_), .Y(_1134__bF_buf13) );
BUFX4 BUFX4_291 ( .A(_1134_), .Y(_1134__bF_buf12) );
BUFX4 BUFX4_292 ( .A(_1134_), .Y(_1134__bF_buf11) );
BUFX4 BUFX4_293 ( .A(_1134_), .Y(_1134__bF_buf10) );
BUFX4 BUFX4_294 ( .A(_1134_), .Y(_1134__bF_buf9) );
BUFX4 BUFX4_295 ( .A(_1134_), .Y(_1134__bF_buf8) );
BUFX4 BUFX4_296 ( .A(_1134_), .Y(_1134__bF_buf7) );
BUFX4 BUFX4_297 ( .A(_1134_), .Y(_1134__bF_buf6) );
BUFX4 BUFX4_298 ( .A(_1134_), .Y(_1134__bF_buf5) );
BUFX4 BUFX4_299 ( .A(_1134_), .Y(_1134__bF_buf4) );
BUFX4 BUFX4_300 ( .A(_1134_), .Y(_1134__bF_buf3) );
BUFX4 BUFX4_301 ( .A(_1134_), .Y(_1134__bF_buf2) );
BUFX4 BUFX4_302 ( .A(_1134_), .Y(_1134__bF_buf1) );
BUFX4 BUFX4_303 ( .A(_1134_), .Y(_1134__bF_buf0) );
BUFX4 BUFX4_304 ( .A(_612_), .Y(_612__bF_buf6) );
BUFX4 BUFX4_305 ( .A(_612_), .Y(_612__bF_buf5) );
BUFX4 BUFX4_306 ( .A(_612_), .Y(_612__bF_buf4) );
BUFX4 BUFX4_307 ( .A(_612_), .Y(_612__bF_buf3) );
BUFX4 BUFX4_308 ( .A(_612_), .Y(_612__bF_buf2) );
BUFX4 BUFX4_309 ( .A(_612_), .Y(_612__bF_buf1) );
BUFX4 BUFX4_310 ( .A(_612_), .Y(_612__bF_buf0) );
BUFX4 BUFX4_311 ( .A(_1031__hier0_bF_buf7), .Y(_1031__bF_buf77) );
BUFX4 BUFX4_312 ( .A(_1031__hier0_bF_buf4), .Y(_1031__bF_buf76) );
BUFX4 BUFX4_313 ( .A(_1031__hier0_bF_buf2), .Y(_1031__bF_buf75) );
BUFX4 BUFX4_314 ( .A(_1031__hier0_bF_buf7), .Y(_1031__bF_buf74) );
BUFX4 BUFX4_315 ( .A(_1031__hier0_bF_buf6), .Y(_1031__bF_buf73) );
BUFX4 BUFX4_316 ( .A(_1031__hier0_bF_buf4), .Y(_1031__bF_buf72) );
BUFX4 BUFX4_317 ( .A(_1031__hier0_bF_buf7), .Y(_1031__bF_buf71) );
BUFX4 BUFX4_318 ( .A(_1031__hier0_bF_buf3), .Y(_1031__bF_buf70) );
BUFX4 BUFX4_319 ( .A(_1031__hier0_bF_buf1), .Y(_1031__bF_buf69) );
BUFX4 BUFX4_320 ( .A(_1031__hier0_bF_buf6), .Y(_1031__bF_buf68) );
BUFX4 BUFX4_321 ( .A(_1031__hier0_bF_buf5), .Y(_1031__bF_buf67) );
BUFX4 BUFX4_322 ( .A(_1031__hier0_bF_buf2), .Y(_1031__bF_buf66) );
BUFX4 BUFX4_323 ( .A(_1031__hier0_bF_buf5), .Y(_1031__bF_buf65) );
BUFX4 BUFX4_324 ( .A(_1031__hier0_bF_buf7), .Y(_1031__bF_buf64) );
BUFX4 BUFX4_325 ( .A(_1031__hier0_bF_buf4), .Y(_1031__bF_buf63) );
BUFX4 BUFX4_326 ( .A(_1031__hier0_bF_buf7), .Y(_1031__bF_buf62) );
BUFX4 BUFX4_327 ( .A(_1031__hier0_bF_buf6), .Y(_1031__bF_buf61) );
BUFX4 BUFX4_328 ( .A(_1031__hier0_bF_buf4), .Y(_1031__bF_buf60) );
BUFX4 BUFX4_329 ( .A(_1031__hier0_bF_buf5), .Y(_1031__bF_buf59) );
BUFX4 BUFX4_330 ( .A(_1031__hier0_bF_buf3), .Y(_1031__bF_buf58) );
BUFX4 BUFX4_331 ( .A(_1031__hier0_bF_buf0), .Y(_1031__bF_buf57) );
BUFX4 BUFX4_332 ( .A(_1031__hier0_bF_buf2), .Y(_1031__bF_buf56) );
BUFX4 BUFX4_333 ( .A(_1031__hier0_bF_buf7), .Y(_1031__bF_buf55) );
BUFX4 BUFX4_334 ( .A(_1031__hier0_bF_buf7), .Y(_1031__bF_buf54) );
BUFX4 BUFX4_335 ( .A(_1031__hier0_bF_buf4), .Y(_1031__bF_buf53) );
BUFX4 BUFX4_336 ( .A(_1031__hier0_bF_buf2), .Y(_1031__bF_buf52) );
BUFX4 BUFX4_337 ( .A(_1031__hier0_bF_buf1), .Y(_1031__bF_buf51) );
BUFX4 BUFX4_338 ( .A(_1031__hier0_bF_buf0), .Y(_1031__bF_buf50) );
BUFX4 BUFX4_339 ( .A(_1031__hier0_bF_buf3), .Y(_1031__bF_buf49) );
BUFX4 BUFX4_340 ( .A(_1031__hier0_bF_buf1), .Y(_1031__bF_buf48) );
BUFX4 BUFX4_341 ( .A(_1031__hier0_bF_buf2), .Y(_1031__bF_buf47) );
BUFX4 BUFX4_342 ( .A(_1031__hier0_bF_buf3), .Y(_1031__bF_buf46) );
BUFX4 BUFX4_343 ( .A(_1031__hier0_bF_buf0), .Y(_1031__bF_buf45) );
BUFX4 BUFX4_344 ( .A(_1031__hier0_bF_buf3), .Y(_1031__bF_buf44) );
BUFX4 BUFX4_345 ( .A(_1031__hier0_bF_buf6), .Y(_1031__bF_buf43) );
BUFX4 BUFX4_346 ( .A(_1031__hier0_bF_buf4), .Y(_1031__bF_buf42) );
BUFX4 BUFX4_347 ( .A(_1031__hier0_bF_buf5), .Y(_1031__bF_buf41) );
BUFX4 BUFX4_348 ( .A(_1031__hier0_bF_buf3), .Y(_1031__bF_buf40) );
BUFX4 BUFX4_349 ( .A(_1031__hier0_bF_buf2), .Y(_1031__bF_buf39) );
BUFX4 BUFX4_350 ( .A(_1031__hier0_bF_buf0), .Y(_1031__bF_buf38) );
BUFX4 BUFX4_351 ( .A(_1031__hier0_bF_buf1), .Y(_1031__bF_buf37) );
BUFX4 BUFX4_352 ( .A(_1031__hier0_bF_buf5), .Y(_1031__bF_buf36) );
BUFX4 BUFX4_353 ( .A(_1031__hier0_bF_buf4), .Y(_1031__bF_buf35) );
BUFX4 BUFX4_354 ( .A(_1031__hier0_bF_buf7), .Y(_1031__bF_buf34) );
BUFX4 BUFX4_355 ( .A(_1031__hier0_bF_buf6), .Y(_1031__bF_buf33) );
BUFX4 BUFX4_356 ( .A(_1031__hier0_bF_buf1), .Y(_1031__bF_buf32) );
BUFX4 BUFX4_357 ( .A(_1031__hier0_bF_buf3), .Y(_1031__bF_buf31) );
BUFX4 BUFX4_358 ( .A(_1031__hier0_bF_buf6), .Y(_1031__bF_buf30) );
BUFX4 BUFX4_359 ( .A(_1031__hier0_bF_buf1), .Y(_1031__bF_buf29) );
BUFX4 BUFX4_360 ( .A(_1031__hier0_bF_buf3), .Y(_1031__bF_buf28) );
BUFX4 BUFX4_361 ( .A(_1031__hier0_bF_buf2), .Y(_1031__bF_buf27) );
BUFX4 BUFX4_362 ( .A(_1031__hier0_bF_buf5), .Y(_1031__bF_buf26) );
BUFX4 BUFX4_363 ( .A(_1031__hier0_bF_buf2), .Y(_1031__bF_buf25) );
BUFX4 BUFX4_364 ( .A(_1031__hier0_bF_buf0), .Y(_1031__bF_buf24) );
BUFX4 BUFX4_365 ( .A(_1031__hier0_bF_buf6), .Y(_1031__bF_buf23) );
BUFX4 BUFX4_366 ( .A(_1031__hier0_bF_buf5), .Y(_1031__bF_buf22) );
BUFX4 BUFX4_367 ( .A(_1031__hier0_bF_buf5), .Y(_1031__bF_buf21) );
BUFX4 BUFX4_368 ( .A(_1031__hier0_bF_buf5), .Y(_1031__bF_buf20) );
BUFX4 BUFX4_369 ( .A(_1031__hier0_bF_buf0), .Y(_1031__bF_buf19) );
BUFX4 BUFX4_370 ( .A(_1031__hier0_bF_buf0), .Y(_1031__bF_buf18) );
BUFX4 BUFX4_371 ( .A(_1031__hier0_bF_buf7), .Y(_1031__bF_buf17) );
BUFX4 BUFX4_372 ( .A(_1031__hier0_bF_buf6), .Y(_1031__bF_buf16) );
BUFX4 BUFX4_373 ( .A(_1031__hier0_bF_buf4), .Y(_1031__bF_buf15) );
BUFX4 BUFX4_374 ( .A(_1031__hier0_bF_buf0), .Y(_1031__bF_buf14) );
BUFX4 BUFX4_375 ( .A(_1031__hier0_bF_buf3), .Y(_1031__bF_buf13) );
BUFX4 BUFX4_376 ( .A(_1031__hier0_bF_buf5), .Y(_1031__bF_buf12) );
BUFX4 BUFX4_377 ( .A(_1031__hier0_bF_buf2), .Y(_1031__bF_buf11) );
BUFX4 BUFX4_378 ( .A(_1031__hier0_bF_buf7), .Y(_1031__bF_buf10) );
BUFX4 BUFX4_379 ( .A(_1031__hier0_bF_buf1), .Y(_1031__bF_buf9) );
BUFX4 BUFX4_380 ( .A(_1031__hier0_bF_buf2), .Y(_1031__bF_buf8) );
BUFX4 BUFX4_381 ( .A(_1031__hier0_bF_buf3), .Y(_1031__bF_buf7) );
BUFX4 BUFX4_382 ( .A(_1031__hier0_bF_buf4), .Y(_1031__bF_buf6) );
BUFX4 BUFX4_383 ( .A(_1031__hier0_bF_buf1), .Y(_1031__bF_buf5) );
BUFX4 BUFX4_384 ( .A(_1031__hier0_bF_buf0), .Y(_1031__bF_buf4) );
BUFX4 BUFX4_385 ( .A(_1031__hier0_bF_buf1), .Y(_1031__bF_buf3) );
BUFX4 BUFX4_386 ( .A(_1031__hier0_bF_buf4), .Y(_1031__bF_buf2) );
BUFX4 BUFX4_387 ( .A(_1031__hier0_bF_buf6), .Y(_1031__bF_buf1) );
BUFX4 BUFX4_388 ( .A(_1031__hier0_bF_buf6), .Y(_1031__bF_buf0) );
INVX2 INVX2_1 ( .A(bundleTid_i[6]), .Y(_1282_) );
NAND2X1 NAND2X1_1 ( .A(_3660__6_), .B(_1031__bF_buf9), .Y(_1283_) );
OAI21X1 OAI21X1_1 ( .A(_1031__bF_buf9), .B(_1282_), .C(_1283_), .Y(_156_) );
INVX2 INVX2_2 ( .A(bundleTid_i[5]), .Y(_1284_) );
NAND2X1 NAND2X1_2 ( .A(_3660__5_), .B(_1031__bF_buf55), .Y(_1285_) );
OAI21X1 OAI21X1_2 ( .A(_1031__bF_buf55), .B(_1284_), .C(_1285_), .Y(_157_) );
INVX2 INVX2_3 ( .A(bundleTid_i[4]), .Y(_1286_) );
NAND2X1 NAND2X1_3 ( .A(_3660__4_), .B(_1031__bF_buf19), .Y(_1287_) );
OAI21X1 OAI21X1_3 ( .A(_1031__bF_buf19), .B(_1286_), .C(_1287_), .Y(_158_) );
INVX2 INVX2_4 ( .A(bundleTid_i[3]), .Y(_1288_) );
NAND2X1 NAND2X1_4 ( .A(_3660__3_), .B(_1031__bF_buf19), .Y(_1289_) );
OAI21X1 OAI21X1_4 ( .A(_1031__bF_buf19), .B(_1288_), .C(_1289_), .Y(_159_) );
INVX2 INVX2_5 ( .A(bundleTid_i[2]), .Y(_1290_) );
NAND2X1 NAND2X1_5 ( .A(_3660__2_), .B(_1031__bF_buf17), .Y(_1291_) );
OAI21X1 OAI21X1_5 ( .A(_1031__bF_buf17), .B(_1290_), .C(_1291_), .Y(_160_) );
INVX2 INVX2_6 ( .A(bundleTid_i[1]), .Y(_1292_) );
NAND2X1 NAND2X1_6 ( .A(_3660__1_), .B(_1031__bF_buf61), .Y(_1293_) );
OAI21X1 OAI21X1_6 ( .A(_1031__bF_buf61), .B(_1292_), .C(_1293_), .Y(_161_) );
INVX2 INVX2_7 ( .A(bundleTid_i[0]), .Y(_1294_) );
NAND2X1 NAND2X1_7 ( .A(_3660__0_), .B(_1031__bF_buf57), .Y(_1295_) );
OAI21X1 OAI21X1_7 ( .A(_1031__bF_buf50), .B(_1294_), .C(_1295_), .Y(_162_) );
NAND2X1 NAND2X1_8 ( .A(_3661__63_), .B(_1039__bF_buf27), .Y(_1296_) );
OAI21X1 OAI21X1_8 ( .A(_1168_), .B(_1039__bF_buf27), .C(_1296_), .Y(_163_) );
NAND2X1 NAND2X1_9 ( .A(_3661__62_), .B(_1039__bF_buf52), .Y(_1297_) );
OAI21X1 OAI21X1_9 ( .A(_1170_), .B(_1039__bF_buf52), .C(_1297_), .Y(_164_) );
NAND2X1 NAND2X1_10 ( .A(_3661__61_), .B(_1039__bF_buf4), .Y(_1298_) );
OAI21X1 OAI21X1_10 ( .A(_1172_), .B(_1039__bF_buf4), .C(_1298_), .Y(_165_) );
NAND2X1 NAND2X1_11 ( .A(_3661__60_), .B(_1039__bF_buf15), .Y(_1299_) );
OAI21X1 OAI21X1_11 ( .A(_1174_), .B(_1039__bF_buf15), .C(_1299_), .Y(_166_) );
NAND2X1 NAND2X1_12 ( .A(_3661__59_), .B(_1039__bF_buf40), .Y(_1300_) );
OAI21X1 OAI21X1_12 ( .A(_1176_), .B(_1039__bF_buf40), .C(_1300_), .Y(_167_) );
NAND2X1 NAND2X1_13 ( .A(_3661__58_), .B(_1039__bF_buf41), .Y(_1301_) );
OAI21X1 OAI21X1_13 ( .A(_1178_), .B(_1039__bF_buf41), .C(_1301_), .Y(_168_) );
NAND2X1 NAND2X1_14 ( .A(_3661__57_), .B(_1039__bF_buf18), .Y(_1302_) );
OAI21X1 OAI21X1_14 ( .A(_1180_), .B(_1039__bF_buf18), .C(_1302_), .Y(_169_) );
NAND2X1 NAND2X1_15 ( .A(_3661__56_), .B(_1039__bF_buf18), .Y(_1303_) );
OAI21X1 OAI21X1_15 ( .A(_1182_), .B(_1039__bF_buf18), .C(_1303_), .Y(_170_) );
NAND2X1 NAND2X1_16 ( .A(_3661__55_), .B(_1039__bF_buf0), .Y(_1304_) );
OAI21X1 OAI21X1_16 ( .A(_1184_), .B(_1039__bF_buf0), .C(_1304_), .Y(_171_) );
NAND2X1 NAND2X1_17 ( .A(_3661__54_), .B(_1039__bF_buf13), .Y(_1305_) );
OAI21X1 OAI21X1_17 ( .A(_1186_), .B(_1039__bF_buf13), .C(_1305_), .Y(_172_) );
NAND2X1 NAND2X1_18 ( .A(_3661__53_), .B(_1039__bF_buf52), .Y(_1306_) );
OAI21X1 OAI21X1_18 ( .A(_1188_), .B(_1039__bF_buf52), .C(_1306_), .Y(_173_) );
NAND2X1 NAND2X1_19 ( .A(_3661__52_), .B(_1039__bF_buf17), .Y(_1307_) );
OAI21X1 OAI21X1_19 ( .A(_1190_), .B(_1039__bF_buf46), .C(_1307_), .Y(_174_) );
NAND2X1 NAND2X1_20 ( .A(_3661__51_), .B(_1039__bF_buf10), .Y(_1308_) );
OAI21X1 OAI21X1_20 ( .A(_1192_), .B(_1039__bF_buf10), .C(_1308_), .Y(_175_) );
NAND2X1 NAND2X1_21 ( .A(_3661__50_), .B(_1039__bF_buf0), .Y(_1309_) );
OAI21X1 OAI21X1_21 ( .A(_1194_), .B(_1039__bF_buf0), .C(_1309_), .Y(_176_) );
NAND2X1 NAND2X1_22 ( .A(_3661__49_), .B(_1039__bF_buf19), .Y(_1310_) );
OAI21X1 OAI21X1_22 ( .A(_1196_), .B(_1039__bF_buf19), .C(_1310_), .Y(_177_) );
NAND2X1 NAND2X1_23 ( .A(_3661__48_), .B(_1039__bF_buf21), .Y(_1311_) );
OAI21X1 OAI21X1_23 ( .A(_1198_), .B(_1039__bF_buf21), .C(_1311_), .Y(_178_) );
NAND2X1 NAND2X1_24 ( .A(_3661__47_), .B(_1039__bF_buf14), .Y(_1312_) );
OAI21X1 OAI21X1_24 ( .A(_1200_), .B(_1039__bF_buf14), .C(_1312_), .Y(_179_) );
NAND2X1 NAND2X1_25 ( .A(_3661__46_), .B(_1039__bF_buf21), .Y(_1313_) );
OAI21X1 OAI21X1_25 ( .A(_1202_), .B(_1039__bF_buf39), .C(_1313_), .Y(_180_) );
NAND2X1 NAND2X1_26 ( .A(_3661__45_), .B(_1039__bF_buf18), .Y(_1314_) );
OAI21X1 OAI21X1_26 ( .A(_1204_), .B(_1039__bF_buf50), .C(_1314_), .Y(_181_) );
NAND2X1 NAND2X1_27 ( .A(_3661__44_), .B(_1039__bF_buf29), .Y(_1315_) );
OAI21X1 OAI21X1_27 ( .A(_1206_), .B(_1039__bF_buf37), .C(_1315_), .Y(_182_) );
NAND2X1 NAND2X1_28 ( .A(_3661__43_), .B(_1039__bF_buf4), .Y(_1316_) );
OAI21X1 OAI21X1_28 ( .A(_1208_), .B(_1039__bF_buf4), .C(_1316_), .Y(_183_) );
NAND2X1 NAND2X1_29 ( .A(_3661__42_), .B(_1039__bF_buf37), .Y(_1317_) );
OAI21X1 OAI21X1_29 ( .A(_1210_), .B(_1039__bF_buf37), .C(_1317_), .Y(_184_) );
NAND2X1 NAND2X1_30 ( .A(_3661__41_), .B(_1039__bF_buf42), .Y(_1318_) );
OAI21X1 OAI21X1_30 ( .A(_1212_), .B(_1039__bF_buf42), .C(_1318_), .Y(_185_) );
NAND2X1 NAND2X1_31 ( .A(_3661__40_), .B(_1039__bF_buf42), .Y(_1319_) );
OAI21X1 OAI21X1_31 ( .A(_1214_), .B(_1039__bF_buf42), .C(_1319_), .Y(_186_) );
NAND2X1 NAND2X1_32 ( .A(_3661__39_), .B(_1039__bF_buf30), .Y(_1320_) );
OAI21X1 OAI21X1_32 ( .A(_1216_), .B(_1039__bF_buf30), .C(_1320_), .Y(_187_) );
NAND2X1 NAND2X1_33 ( .A(_3661__38_), .B(_1039__bF_buf46), .Y(_1321_) );
OAI21X1 OAI21X1_33 ( .A(_1218_), .B(_1039__bF_buf8), .C(_1321_), .Y(_188_) );
NAND2X1 NAND2X1_34 ( .A(_3661__37_), .B(_1039__bF_buf46), .Y(_1322_) );
OAI21X1 OAI21X1_34 ( .A(_1220_), .B(_1039__bF_buf46), .C(_1322_), .Y(_189_) );
NAND2X1 NAND2X1_35 ( .A(_3661__36_), .B(_1039__bF_buf3), .Y(_1323_) );
OAI21X1 OAI21X1_35 ( .A(_1222_), .B(_1039__bF_buf3), .C(_1323_), .Y(_190_) );
NAND2X1 NAND2X1_36 ( .A(_3661__35_), .B(_1039__bF_buf41), .Y(_1324_) );
OAI21X1 OAI21X1_36 ( .A(_1224_), .B(_1039__bF_buf41), .C(_1324_), .Y(_191_) );
NAND2X1 NAND2X1_37 ( .A(_3661__34_), .B(_1039__bF_buf48), .Y(_1325_) );
OAI21X1 OAI21X1_37 ( .A(_1226_), .B(_1039__bF_buf36), .C(_1325_), .Y(_192_) );
NAND2X1 NAND2X1_38 ( .A(_3661__33_), .B(_1039__bF_buf27), .Y(_1326_) );
OAI21X1 OAI21X1_38 ( .A(_1228_), .B(_1039__bF_buf27), .C(_1326_), .Y(_193_) );
NAND2X1 NAND2X1_39 ( .A(_3661__32_), .B(_1039__bF_buf7), .Y(_1327_) );
OAI21X1 OAI21X1_39 ( .A(_1230_), .B(_1039__bF_buf7), .C(_1327_), .Y(_194_) );
NAND2X1 NAND2X1_40 ( .A(_3661__31_), .B(_1039__bF_buf22), .Y(_1328_) );
OAI21X1 OAI21X1_40 ( .A(_1232_), .B(_1039__bF_buf22), .C(_1328_), .Y(_195_) );
NAND2X1 NAND2X1_41 ( .A(_3661__30_), .B(_1039__bF_buf29), .Y(_1329_) );
OAI21X1 OAI21X1_41 ( .A(_1234_), .B(_1039__bF_buf29), .C(_1329_), .Y(_196_) );
NAND2X1 NAND2X1_42 ( .A(_3661__29_), .B(_1039__bF_buf3), .Y(_1330_) );
OAI21X1 OAI21X1_42 ( .A(_1236_), .B(_1039__bF_buf3), .C(_1330_), .Y(_197_) );
NAND2X1 NAND2X1_43 ( .A(_3661__28_), .B(_1039__bF_buf54), .Y(_1331_) );
OAI21X1 OAI21X1_43 ( .A(_1238_), .B(_1039__bF_buf54), .C(_1331_), .Y(_198_) );
NAND2X1 NAND2X1_44 ( .A(_3661__27_), .B(_1039__bF_buf14), .Y(_1332_) );
OAI21X1 OAI21X1_44 ( .A(_1240_), .B(_1039__bF_buf8), .C(_1332_), .Y(_199_) );
NAND2X1 NAND2X1_45 ( .A(_3661__26_), .B(_1039__bF_buf37), .Y(_1333_) );
OAI21X1 OAI21X1_45 ( .A(_1242_), .B(_1039__bF_buf37), .C(_1333_), .Y(_200_) );
NAND2X1 NAND2X1_46 ( .A(_3661__25_), .B(_1039__bF_buf44), .Y(_1334_) );
OAI21X1 OAI21X1_46 ( .A(_1244_), .B(_1039__bF_buf10), .C(_1334_), .Y(_201_) );
NAND2X1 NAND2X1_47 ( .A(_3661__24_), .B(_1039__bF_buf49), .Y(_1335_) );
OAI21X1 OAI21X1_47 ( .A(_1246_), .B(_1039__bF_buf49), .C(_1335_), .Y(_202_) );
NAND2X1 NAND2X1_48 ( .A(_3661__23_), .B(_1039__bF_buf47), .Y(_1336_) );
OAI21X1 OAI21X1_48 ( .A(_1248_), .B(_1039__bF_buf47), .C(_1336_), .Y(_203_) );
NAND2X1 NAND2X1_49 ( .A(_3661__22_), .B(_1039__bF_buf49), .Y(_1337_) );
OAI21X1 OAI21X1_49 ( .A(_1250_), .B(_1039__bF_buf49), .C(_1337_), .Y(_204_) );
NAND2X1 NAND2X1_50 ( .A(_3661__21_), .B(_1039__bF_buf9), .Y(_1338_) );
OAI21X1 OAI21X1_50 ( .A(_1252_), .B(_1039__bF_buf9), .C(_1338_), .Y(_205_) );
NAND2X1 NAND2X1_51 ( .A(_3661__20_), .B(_1039__bF_buf44), .Y(_1339_) );
OAI21X1 OAI21X1_51 ( .A(_1254_), .B(_1039__bF_buf44), .C(_1339_), .Y(_206_) );
NAND2X1 NAND2X1_52 ( .A(_3661__19_), .B(_1039__bF_buf46), .Y(_1340_) );
OAI21X1 OAI21X1_52 ( .A(_1256_), .B(_1039__bF_buf46), .C(_1340_), .Y(_207_) );
NAND2X1 NAND2X1_53 ( .A(_3661__18_), .B(_1039__bF_buf39), .Y(_1341_) );
OAI21X1 OAI21X1_53 ( .A(_1258_), .B(_1039__bF_buf39), .C(_1341_), .Y(_208_) );
NAND2X1 NAND2X1_54 ( .A(_3661__17_), .B(_1039__bF_buf15), .Y(_1342_) );
OAI21X1 OAI21X1_54 ( .A(_1260_), .B(_1039__bF_buf15), .C(_1342_), .Y(_209_) );
NAND2X1 NAND2X1_55 ( .A(_3661__16_), .B(_1039__bF_buf30), .Y(_1343_) );
OAI21X1 OAI21X1_55 ( .A(_1262_), .B(_1039__bF_buf30), .C(_1343_), .Y(_210_) );
NAND2X1 NAND2X1_56 ( .A(_3661__15_), .B(_1039__bF_buf46), .Y(_1344_) );
OAI21X1 OAI21X1_56 ( .A(_1264_), .B(_1039__bF_buf46), .C(_1344_), .Y(_211_) );
NAND2X1 NAND2X1_57 ( .A(_3661__14_), .B(_1039__bF_buf42), .Y(_1345_) );
OAI21X1 OAI21X1_57 ( .A(_1266_), .B(_1039__bF_buf42), .C(_1345_), .Y(_212_) );
NAND2X1 NAND2X1_58 ( .A(_3661__13_), .B(_1039__bF_buf19), .Y(_1346_) );
OAI21X1 OAI21X1_58 ( .A(_1268_), .B(_1039__bF_buf19), .C(_1346_), .Y(_213_) );
NAND2X1 NAND2X1_59 ( .A(_3661__12_), .B(_1039__bF_buf18), .Y(_1347_) );
OAI21X1 OAI21X1_59 ( .A(_1270_), .B(_1039__bF_buf18), .C(_1347_), .Y(_214_) );
NAND2X1 NAND2X1_60 ( .A(_3661__11_), .B(_1039__bF_buf47), .Y(_1348_) );
OAI21X1 OAI21X1_60 ( .A(_1272_), .B(_1039__bF_buf47), .C(_1348_), .Y(_215_) );
NAND2X1 NAND2X1_61 ( .A(_3661__10_), .B(_1039__bF_buf17), .Y(_1349_) );
OAI21X1 OAI21X1_61 ( .A(_1274_), .B(_1039__bF_buf17), .C(_1349_), .Y(_216_) );
NAND2X1 NAND2X1_62 ( .A(_3661__9_), .B(_1039__bF_buf29), .Y(_1350_) );
OAI21X1 OAI21X1_62 ( .A(_1276_), .B(_1039__bF_buf29), .C(_1350_), .Y(_217_) );
NAND2X1 NAND2X1_63 ( .A(_3661__8_), .B(_1039__bF_buf57), .Y(_1351_) );
OAI21X1 OAI21X1_63 ( .A(_1278_), .B(_1039__bF_buf57), .C(_1351_), .Y(_218_) );
NAND2X1 NAND2X1_64 ( .A(_3661__7_), .B(_1039__bF_buf30), .Y(_1352_) );
OAI21X1 OAI21X1_64 ( .A(_1280_), .B(_1039__bF_buf30), .C(_1352_), .Y(_219_) );
NAND2X1 NAND2X1_65 ( .A(_3661__6_), .B(_1039__bF_buf14), .Y(_1353_) );
OAI21X1 OAI21X1_65 ( .A(_1282_), .B(_1039__bF_buf14), .C(_1353_), .Y(_220_) );
NAND2X1 NAND2X1_66 ( .A(_3661__5_), .B(_1039__bF_buf47), .Y(_1354_) );
OAI21X1 OAI21X1_66 ( .A(_1284_), .B(_1039__bF_buf47), .C(_1354_), .Y(_221_) );
NAND2X1 NAND2X1_67 ( .A(_3661__4_), .B(_1039__bF_buf52), .Y(_1355_) );
OAI21X1 OAI21X1_67 ( .A(_1286_), .B(_1039__bF_buf52), .C(_1355_), .Y(_222_) );
NAND2X1 NAND2X1_68 ( .A(_3661__3_), .B(_1039__bF_buf51), .Y(_1356_) );
OAI21X1 OAI21X1_68 ( .A(_1288_), .B(_1039__bF_buf51), .C(_1356_), .Y(_223_) );
NAND2X1 NAND2X1_69 ( .A(_3661__2_), .B(_1039__bF_buf7), .Y(_1357_) );
OAI21X1 OAI21X1_69 ( .A(_1290_), .B(_1039__bF_buf7), .C(_1357_), .Y(_224_) );
NAND2X1 NAND2X1_70 ( .A(_3661__1_), .B(_1039__bF_buf20), .Y(_1358_) );
OAI21X1 OAI21X1_70 ( .A(_1292_), .B(_1039__bF_buf20), .C(_1358_), .Y(_225_) );
NAND2X1 NAND2X1_71 ( .A(_3661__0_), .B(_1039__bF_buf41), .Y(_1359_) );
OAI21X1 OAI21X1_71 ( .A(_1294_), .B(_1039__bF_buf41), .C(_1359_), .Y(_226_) );
OAI21X1 OAI21X1_72 ( .A(_1100__bF_buf14_bF_buf2), .B(_1031__bF_buf29), .C(_3662__63_), .Y(_1360_) );
OAI21X1 OAI21X1_73 ( .A(_1101__bF_buf30), .B(_1168_), .C(_1360_), .Y(_227_) );
OAI21X1 OAI21X1_74 ( .A(_1100__bF_buf13_bF_buf2), .B(_1031__bF_buf70), .C(_3662__62_), .Y(_1361_) );
OAI21X1 OAI21X1_75 ( .A(_1101__bF_buf13), .B(_1170_), .C(_1361_), .Y(_228_) );
OAI21X1 OAI21X1_76 ( .A(_1100__bF_buf12_bF_buf3), .B(_1031__bF_buf15), .C(_3662__61_), .Y(_1362_) );
OAI21X1 OAI21X1_77 ( .A(_1101__bF_buf48), .B(_1172_), .C(_1362_), .Y(_229_) );
OAI21X1 OAI21X1_78 ( .A(_1100__bF_buf11_bF_buf2), .B(_1031__bF_buf67), .C(_3662__60_), .Y(_1363_) );
OAI21X1 OAI21X1_79 ( .A(_1101__bF_buf44), .B(_1174_), .C(_1363_), .Y(_230_) );
OAI21X1 OAI21X1_80 ( .A(_1100__bF_buf10_bF_buf2), .B(_1031__bF_buf76), .C(_3662__59_), .Y(_1364_) );
OAI21X1 OAI21X1_81 ( .A(_1101__bF_buf47), .B(_1176_), .C(_1364_), .Y(_231_) );
OAI21X1 OAI21X1_82 ( .A(_1100__bF_buf9_bF_buf0), .B(_1031__bF_buf14), .C(_3662__58_), .Y(_1365_) );
OAI21X1 OAI21X1_83 ( .A(_1101__bF_buf40), .B(_1178_), .C(_1365_), .Y(_232_) );
OAI21X1 OAI21X1_84 ( .A(_1100__bF_buf8_bF_buf3), .B(_1031__bF_buf47), .C(_3662__57_), .Y(_1366_) );
OAI21X1 OAI21X1_85 ( .A(_1101__bF_buf9), .B(_1180_), .C(_1366_), .Y(_233_) );
OAI21X1 OAI21X1_86 ( .A(_1100__bF_buf7_bF_buf3), .B(_1031__bF_buf40), .C(_3662__56_), .Y(_1367_) );
OAI21X1 OAI21X1_87 ( .A(_1101__bF_buf17), .B(_1182_), .C(_1367_), .Y(_234_) );
OAI21X1 OAI21X1_88 ( .A(_1100__bF_buf6), .B(_1031__bF_buf73), .C(_3662__55_), .Y(_1368_) );
OAI21X1 OAI21X1_89 ( .A(_1101__bF_buf26), .B(_1184_), .C(_1368_), .Y(_235_) );
OAI21X1 OAI21X1_90 ( .A(_1100__bF_buf10), .B(_1031__bF_buf48), .C(_3662__54_), .Y(_1369_) );
OAI21X1 OAI21X1_91 ( .A(_1101__bF_buf29), .B(_1186_), .C(_1369_), .Y(_236_) );
OAI21X1 OAI21X1_92 ( .A(_1100__bF_buf1), .B(_1031__bF_buf64), .C(_3662__53_), .Y(_1370_) );
OAI21X1 OAI21X1_93 ( .A(_1101__bF_buf50), .B(_1188_), .C(_1370_), .Y(_237_) );
OAI21X1 OAI21X1_94 ( .A(_1100__bF_buf3), .B(_1031__bF_buf70), .C(_3662__52_), .Y(_1371_) );
OAI21X1 OAI21X1_95 ( .A(_1101__bF_buf1), .B(_1190_), .C(_1371_), .Y(_238_) );
OAI21X1 OAI21X1_96 ( .A(_1100__bF_buf3), .B(_1031__bF_buf66), .C(_3662__51_), .Y(_1372_) );
OAI21X1 OAI21X1_97 ( .A(_1101__bF_buf14), .B(_1192_), .C(_1372_), .Y(_239_) );
OAI21X1 OAI21X1_98 ( .A(_1100__bF_buf6), .B(_1031__bF_buf73), .C(_3662__50_), .Y(_1373_) );
OAI21X1 OAI21X1_99 ( .A(_1101__bF_buf26), .B(_1194_), .C(_1373_), .Y(_240_) );
OAI21X1 OAI21X1_100 ( .A(_1100__bF_buf3), .B(_1031__bF_buf47), .C(_3662__49_), .Y(_1374_) );
OAI21X1 OAI21X1_101 ( .A(_1101__bF_buf14), .B(_1196_), .C(_1374_), .Y(_241_) );
OAI21X1 OAI21X1_102 ( .A(_1100__bF_buf14_bF_buf0), .B(_1031__bF_buf35), .C(_3662__48_), .Y(_1375_) );
OAI21X1 OAI21X1_103 ( .A(_1101__bF_buf47), .B(_1198_), .C(_1375_), .Y(_242_) );
OAI21X1 OAI21X1_104 ( .A(_1100__bF_buf13_bF_buf0), .B(_1031__bF_buf54), .C(_3662__47_), .Y(_1376_) );
OAI21X1 OAI21X1_105 ( .A(_1101__bF_buf32), .B(_1200_), .C(_1376_), .Y(_243_) );
OAI21X1 OAI21X1_106 ( .A(_1100__bF_buf12_bF_buf3), .B(_1031__bF_buf76), .C(_3662__46_), .Y(_1377_) );
OAI21X1 OAI21X1_107 ( .A(_1101__bF_buf47), .B(_1202_), .C(_1377_), .Y(_244_) );
OAI21X1 OAI21X1_108 ( .A(_1100__bF_buf11_bF_buf3), .B(_1031__bF_buf11), .C(_3662__45_), .Y(_1378_) );
OAI21X1 OAI21X1_109 ( .A(_1101__bF_buf41), .B(_1204_), .C(_1378_), .Y(_245_) );
OAI21X1 OAI21X1_110 ( .A(_1100__bF_buf10_bF_buf1), .B(_1031__bF_buf54), .C(_3662__44_), .Y(_1379_) );
OAI21X1 OAI21X1_111 ( .A(_1101__bF_buf52), .B(_1206_), .C(_1379_), .Y(_246_) );
OAI21X1 OAI21X1_112 ( .A(_1100__bF_buf9_bF_buf2), .B(_1031__bF_buf48), .C(_3662__43_), .Y(_1380_) );
OAI21X1 OAI21X1_113 ( .A(_1101__bF_buf29), .B(_1208_), .C(_1380_), .Y(_247_) );
OAI21X1 OAI21X1_114 ( .A(_1100__bF_buf8_bF_buf0), .B(_1031__bF_buf20), .C(_3662__42_), .Y(_1381_) );
OAI21X1 OAI21X1_115 ( .A(_1101__bF_buf43), .B(_1210_), .C(_1381_), .Y(_248_) );
OAI21X1 OAI21X1_116 ( .A(_1100__bF_buf7_bF_buf3), .B(_1031__bF_buf40), .C(_3662__41_), .Y(_1382_) );
OAI21X1 OAI21X1_117 ( .A(_1101__bF_buf17), .B(_1212_), .C(_1382_), .Y(_249_) );
OAI21X1 OAI21X1_118 ( .A(_1100__bF_buf3), .B(_1031__bF_buf66), .C(_3662__40_), .Y(_1383_) );
OAI21X1 OAI21X1_119 ( .A(_1101__bF_buf7), .B(_1214_), .C(_1383_), .Y(_250_) );
OAI21X1 OAI21X1_120 ( .A(_1100__bF_buf12), .B(_1031__bF_buf27), .C(_3662__39_), .Y(_1384_) );
OAI21X1 OAI21X1_121 ( .A(_1101__bF_buf11), .B(_1216_), .C(_1384_), .Y(_251_) );
OAI21X1 OAI21X1_122 ( .A(_1100__bF_buf5), .B(_1031__bF_buf71), .C(_3662__38_), .Y(_1385_) );
OAI21X1 OAI21X1_123 ( .A(_1101__bF_buf41), .B(_1218_), .C(_1385_), .Y(_252_) );
OAI21X1 OAI21X1_124 ( .A(_1100__bF_buf5), .B(_1031__bF_buf25), .C(_3662__37_), .Y(_1386_) );
OAI21X1 OAI21X1_125 ( .A(_1101__bF_buf31), .B(_1220_), .C(_1386_), .Y(_253_) );
OAI21X1 OAI21X1_126 ( .A(_1100__bF_buf3), .B(_1031__bF_buf56), .C(_3662__36_), .Y(_1387_) );
OAI21X1 OAI21X1_127 ( .A(_1101__bF_buf56), .B(_1222_), .C(_1387_), .Y(_254_) );
OAI21X1 OAI21X1_128 ( .A(_1100__bF_buf2), .B(_1031__bF_buf45), .C(_3662__35_), .Y(_1388_) );
OAI21X1 OAI21X1_129 ( .A(_1101__bF_buf21), .B(_1224_), .C(_1388_), .Y(_255_) );
OAI21X1 OAI21X1_130 ( .A(_1100__bF_buf1), .B(_1031__bF_buf18), .C(_3662__34_), .Y(_1389_) );
OAI21X1 OAI21X1_131 ( .A(_1101__bF_buf27), .B(_1226_), .C(_1389_), .Y(_256_) );
OAI21X1 OAI21X1_132 ( .A(_1100__bF_buf14_bF_buf2), .B(_1031__bF_buf29), .C(_3662__33_), .Y(_1390_) );
OAI21X1 OAI21X1_133 ( .A(_1101__bF_buf30), .B(_1228_), .C(_1390_), .Y(_257_) );
OAI21X1 OAI21X1_134 ( .A(_1100__bF_buf13_bF_buf1), .B(_1031__bF_buf22), .C(_3662__32_), .Y(_1391_) );
OAI21X1 OAI21X1_135 ( .A(_1101__bF_buf54), .B(_1230_), .C(_1391_), .Y(_258_) );
OAI21X1 OAI21X1_136 ( .A(_1100__bF_buf12_bF_buf2), .B(_1031__bF_buf61), .C(_3662__31_), .Y(_1392_) );
OAI21X1 OAI21X1_137 ( .A(_1101__bF_buf6), .B(_1232_), .C(_1392_), .Y(_259_) );
OAI21X1 OAI21X1_138 ( .A(_1100__bF_buf11_bF_buf0), .B(_1031__bF_buf59), .C(_3662__30_), .Y(_1393_) );
OAI21X1 OAI21X1_139 ( .A(_1101__bF_buf36), .B(_1234_), .C(_1393_), .Y(_260_) );
OAI21X1 OAI21X1_140 ( .A(_1100__bF_buf10_bF_buf2), .B(_1031__bF_buf2), .C(_3662__29_), .Y(_1394_) );
OAI21X1 OAI21X1_141 ( .A(_1101__bF_buf33), .B(_1236_), .C(_1394_), .Y(_261_) );
OAI21X1 OAI21X1_142 ( .A(_1100__bF_buf9_bF_buf3), .B(_1031__bF_buf12), .C(_3662__28_), .Y(_1395_) );
OAI21X1 OAI21X1_143 ( .A(_1101__bF_buf54), .B(_1238_), .C(_1395_), .Y(_262_) );
OAI21X1 OAI21X1_144 ( .A(_1100__bF_buf8_bF_buf3), .B(_1031__bF_buf71), .C(_3662__27_), .Y(_1396_) );
OAI21X1 OAI21X1_145 ( .A(_1101__bF_buf22), .B(_1240_), .C(_1396_), .Y(_263_) );
OAI21X1 OAI21X1_146 ( .A(_1100__bF_buf7_bF_buf1), .B(_1031__bF_buf32), .C(_3662__26_), .Y(_1397_) );
OAI21X1 OAI21X1_147 ( .A(_1101__bF_buf29), .B(_1242_), .C(_1397_), .Y(_264_) );
OAI21X1 OAI21X1_148 ( .A(_1100__bF_buf3), .B(_1031__bF_buf66), .C(_3662__25_), .Y(_1398_) );
OAI21X1 OAI21X1_149 ( .A(_1101__bF_buf42), .B(_1244_), .C(_1398_), .Y(_265_) );
OAI21X1 OAI21X1_150 ( .A(_1100__bF_buf2), .B(_1031__bF_buf58), .C(_3662__24_), .Y(_1399_) );
OAI21X1 OAI21X1_151 ( .A(_1101__bF_buf38), .B(_1246_), .C(_1399_), .Y(_266_) );
OAI21X1 OAI21X1_152 ( .A(_1100__bF_buf5), .B(_1031__bF_buf55), .C(_3662__23_), .Y(_1400_) );
OAI21X1 OAI21X1_153 ( .A(_1101__bF_buf46), .B(_1248_), .C(_1400_), .Y(_267_) );
OAI21X1 OAI21X1_154 ( .A(_1100__bF_buf2), .B(_1031__bF_buf14), .C(_3662__22_), .Y(_1401_) );
OAI21X1 OAI21X1_155 ( .A(_1101__bF_buf40), .B(_1250_), .C(_1401_), .Y(_268_) );
OAI21X1 OAI21X1_156 ( .A(_1100__bF_buf5), .B(_1031__bF_buf62), .C(_3662__21_), .Y(_1402_) );
OAI21X1 OAI21X1_157 ( .A(_1101__bF_buf55), .B(_1252_), .C(_1402_), .Y(_269_) );
OAI21X1 OAI21X1_158 ( .A(_1100__bF_buf3), .B(_1031__bF_buf8), .C(_3662__20_), .Y(_1403_) );
OAI21X1 OAI21X1_159 ( .A(_1101__bF_buf7), .B(_1254_), .C(_1403_), .Y(_270_) );
OAI21X1 OAI21X1_160 ( .A(_1100__bF_buf5), .B(_1031__bF_buf52), .C(_3662__19_), .Y(_1404_) );
OAI21X1 OAI21X1_161 ( .A(_1101__bF_buf31), .B(_1256_), .C(_1404_), .Y(_271_) );
OAI21X1 OAI21X1_162 ( .A(_1100__bF_buf14_bF_buf2), .B(_1031__bF_buf9), .C(_3662__18_), .Y(_1405_) );
OAI21X1 OAI21X1_163 ( .A(_1101__bF_buf15), .B(_1258_), .C(_1405_), .Y(_272_) );
OAI21X1 OAI21X1_164 ( .A(_1100__bF_buf13_bF_buf1), .B(_1031__bF_buf21), .C(_3662__17_), .Y(_1406_) );
OAI21X1 OAI21X1_165 ( .A(_1101__bF_buf45), .B(_1260_), .C(_1406_), .Y(_273_) );
OAI21X1 OAI21X1_166 ( .A(_1100__bF_buf12_bF_buf0), .B(_1031__bF_buf27), .C(_3662__16_), .Y(_1407_) );
OAI21X1 OAI21X1_167 ( .A(_1101__bF_buf20), .B(_1262_), .C(_1407_), .Y(_274_) );
OAI21X1 OAI21X1_168 ( .A(_1100__bF_buf11_bF_buf3), .B(_1031__bF_buf11), .C(_3662__15_), .Y(_1408_) );
OAI21X1 OAI21X1_169 ( .A(_1101__bF_buf31), .B(_1264_), .C(_1408_), .Y(_275_) );
OAI21X1 OAI21X1_170 ( .A(_1100__bF_buf10_bF_buf0), .B(_1031__bF_buf58), .C(_3662__14_), .Y(_1409_) );
OAI21X1 OAI21X1_171 ( .A(_1101__bF_buf38), .B(_1266_), .C(_1409_), .Y(_276_) );
OAI21X1 OAI21X1_172 ( .A(_1100__bF_buf9_bF_buf2), .B(_1031__bF_buf3), .C(_3662__13_), .Y(_1410_) );
OAI21X1 OAI21X1_173 ( .A(_1101__bF_buf15), .B(_1268_), .C(_1410_), .Y(_277_) );
OAI21X1 OAI21X1_174 ( .A(_1100__bF_buf8_bF_buf2), .B(_1031__bF_buf57), .C(_3662__12_), .Y(_1411_) );
OAI21X1 OAI21X1_175 ( .A(_1101__bF_buf35), .B(_1270_), .C(_1411_), .Y(_278_) );
OAI21X1 OAI21X1_176 ( .A(_1100__bF_buf7_bF_buf0), .B(_1031__bF_buf74), .C(_3662__11_), .Y(_1412_) );
OAI21X1 OAI21X1_177 ( .A(_1101__bF_buf49), .B(_1272_), .C(_1412_), .Y(_279_) );
OAI21X1 OAI21X1_178 ( .A(_1100__bF_buf3), .B(_1031__bF_buf70), .C(_3662__10_), .Y(_1413_) );
OAI21X1 OAI21X1_179 ( .A(_1101__bF_buf1), .B(_1274_), .C(_1413_), .Y(_280_) );
OAI21X1 OAI21X1_180 ( .A(_1100__bF_buf13), .B(_1031__bF_buf36), .C(_3662__9_), .Y(_1414_) );
OAI21X1 OAI21X1_181 ( .A(_1101__bF_buf36), .B(_1276_), .C(_1414_), .Y(_281_) );
OAI21X1 OAI21X1_182 ( .A(_1100__bF_buf6), .B(_1031__bF_buf21), .C(_3662__8_), .Y(_1415_) );
OAI21X1 OAI21X1_183 ( .A(_1101__bF_buf45), .B(_1278_), .C(_1415_), .Y(_282_) );
OAI21X1 OAI21X1_184 ( .A(_1100__bF_buf0), .B(_1031__bF_buf29), .C(_3662__7_), .Y(_1416_) );
OAI21X1 OAI21X1_185 ( .A(_1101__bF_buf30), .B(_1280_), .C(_1416_), .Y(_283_) );
OAI21X1 OAI21X1_186 ( .A(_1100__bF_buf12), .B(_1031__bF_buf9), .C(_3662__6_), .Y(_1417_) );
OAI21X1 OAI21X1_187 ( .A(_1101__bF_buf11), .B(_1282_), .C(_1417_), .Y(_284_) );
OAI21X1 OAI21X1_188 ( .A(_1100__bF_buf5), .B(_1031__bF_buf34), .C(_3662__5_), .Y(_1418_) );
OAI21X1 OAI21X1_189 ( .A(_1101__bF_buf46), .B(_1284_), .C(_1418_), .Y(_285_) );
OAI21X1 OAI21X1_190 ( .A(_1100__bF_buf1), .B(_1031__bF_buf18), .C(_3662__4_), .Y(_1419_) );
OAI21X1 OAI21X1_191 ( .A(_1101__bF_buf10), .B(_1286_), .C(_1419_), .Y(_286_) );
OAI21X1 OAI21X1_192 ( .A(_1100__bF_buf14_bF_buf3), .B(_1031__bF_buf34), .C(_3662__3_), .Y(_1420_) );
OAI21X1 OAI21X1_193 ( .A(_1101__bF_buf55), .B(_1288_), .C(_1420_), .Y(_287_) );
OAI21X1 OAI21X1_194 ( .A(_1100__bF_buf13_bF_buf2), .B(_1031__bF_buf77), .C(_3662__2_), .Y(_1421_) );
OAI21X1 OAI21X1_195 ( .A(_1101__bF_buf20), .B(_1290_), .C(_1421_), .Y(_288_) );
OAI21X1 OAI21X1_196 ( .A(_1100__bF_buf12_bF_buf2), .B(_1031__bF_buf21), .C(_3662__1_), .Y(_1422_) );
OAI21X1 OAI21X1_197 ( .A(_1101__bF_buf45), .B(_1292_), .C(_1422_), .Y(_289_) );
OAI21X1 OAI21X1_198 ( .A(_1100__bF_buf11_bF_buf1), .B(_1031__bF_buf57), .C(_3662__0_), .Y(_1423_) );
OAI21X1 OAI21X1_199 ( .A(_1101__bF_buf35), .B(_1294_), .C(_1423_), .Y(_290_) );
OAI21X1 OAI21X1_200 ( .A(_1101__bF_buf30), .B(_1135__bF_buf14_bF_buf3), .C(_3663__63_), .Y(_1424_) );
OAI21X1 OAI21X1_201 ( .A(_1168_), .B(_1134__bF_buf12), .C(_1424_), .Y(_291_) );
OAI21X1 OAI21X1_202 ( .A(_1101__bF_buf10), .B(_1135__bF_buf13_bF_buf0), .C(_3663__62_), .Y(_1425_) );
OAI21X1 OAI21X1_203 ( .A(_1170_), .B(_1134__bF_buf9), .C(_1425_), .Y(_292_) );
OAI21X1 OAI21X1_204 ( .A(_1101__bF_buf2), .B(_1135__bF_buf12_bF_buf0), .C(_3663__61_), .Y(_1426_) );
OAI21X1 OAI21X1_205 ( .A(_1172_), .B(_1134__bF_buf3), .C(_1426_), .Y(_293_) );
OAI21X1 OAI21X1_206 ( .A(_1101__bF_buf4), .B(_1135__bF_buf11_bF_buf3), .C(_3663__60_), .Y(_1427_) );
OAI21X1 OAI21X1_207 ( .A(_1174_), .B(_1134__bF_buf3), .C(_1427_), .Y(_294_) );
OAI21X1 OAI21X1_208 ( .A(_1101__bF_buf15), .B(_1135__bF_buf10_bF_buf2), .C(_3663__59_), .Y(_1428_) );
OAI21X1 OAI21X1_209 ( .A(_1176_), .B(_1134__bF_buf12), .C(_1428_), .Y(_295_) );
OAI21X1 OAI21X1_210 ( .A(_1101__bF_buf21), .B(_1135__bF_buf9_bF_buf3), .C(_3663__58_), .Y(_1429_) );
OAI21X1 OAI21X1_211 ( .A(_1178_), .B(_1134__bF_buf0), .C(_1429_), .Y(_296_) );
OAI21X1 OAI21X1_212 ( .A(_1101__bF_buf5), .B(_1135__bF_buf8_bF_buf2), .C(_3663__57_), .Y(_1430_) );
OAI21X1 OAI21X1_213 ( .A(_1180_), .B(_1134__bF_buf5), .C(_1430_), .Y(_297_) );
OAI21X1 OAI21X1_214 ( .A(_1101__bF_buf17), .B(_1135__bF_buf7_bF_buf3), .C(_3663__56_), .Y(_1431_) );
OAI21X1 OAI21X1_215 ( .A(_1182_), .B(_1134__bF_buf6), .C(_1431_), .Y(_298_) );
OAI21X1 OAI21X1_216 ( .A(_1101__bF_buf44), .B(_1135__bF_buf6_bF_buf1), .C(_3663__55_), .Y(_1432_) );
OAI21X1 OAI21X1_217 ( .A(_1184_), .B(_1134__bF_buf1), .C(_1432_), .Y(_299_) );
OAI21X1 OAI21X1_218 ( .A(_1101__bF_buf23), .B(_1135__bF_buf5_bF_buf3), .C(_3663__54_), .Y(_1433_) );
OAI21X1 OAI21X1_219 ( .A(_1186_), .B(_1134__bF_buf14), .C(_1433_), .Y(_300_) );
OAI21X1 OAI21X1_220 ( .A(_1101__bF_buf55), .B(_1135__bF_buf4_bF_buf2), .C(_3663__53_), .Y(_1434_) );
OAI21X1 OAI21X1_221 ( .A(_1188_), .B(_1134__bF_buf5), .C(_1434_), .Y(_301_) );
OAI21X1 OAI21X1_222 ( .A(_1101__bF_buf31), .B(_1135__bF_buf3_bF_buf3), .C(_3663__52_), .Y(_1435_) );
OAI21X1 OAI21X1_223 ( .A(_1190_), .B(_1134__bF_buf11), .C(_1435_), .Y(_302_) );
OAI21X1 OAI21X1_224 ( .A(_1101__bF_buf14), .B(_1135__bF_buf2_bF_buf0), .C(_3663__51_), .Y(_1436_) );
OAI21X1 OAI21X1_225 ( .A(_1192_), .B(_1134__bF_buf10), .C(_1436_), .Y(_303_) );
OAI21X1 OAI21X1_226 ( .A(_1101__bF_buf16), .B(_1135__bF_buf1_bF_buf0), .C(_3663__50_), .Y(_1437_) );
OAI21X1 OAI21X1_227 ( .A(_1194_), .B(_1134__bF_buf1), .C(_1437_), .Y(_304_) );
OAI21X1 OAI21X1_228 ( .A(_1101__bF_buf14), .B(_1135__bF_buf11), .C(_3663__49_), .Y(_1438_) );
OAI21X1 OAI21X1_229 ( .A(_1196_), .B(_1134__bF_buf10), .C(_1438_), .Y(_305_) );
OAI21X1 OAI21X1_230 ( .A(_1101__bF_buf47), .B(_1135__bF_buf14_bF_buf0), .C(_3663__48_), .Y(_1439_) );
OAI21X1 OAI21X1_231 ( .A(_1198_), .B(_1134__bF_buf13), .C(_1439_), .Y(_306_) );
OAI21X1 OAI21X1_232 ( .A(_1101__bF_buf32), .B(_1135__bF_buf13_bF_buf1), .C(_3663__47_), .Y(_1440_) );
OAI21X1 OAI21X1_233 ( .A(_1200_), .B(_1134__bF_buf8), .C(_1440_), .Y(_307_) );
OAI21X1 OAI21X1_234 ( .A(_1101__bF_buf29), .B(_1135__bF_buf12_bF_buf3), .C(_3663__46_), .Y(_1441_) );
OAI21X1 OAI21X1_235 ( .A(_1202_), .B(_1134__bF_buf14), .C(_1441_), .Y(_308_) );
OAI21X1 OAI21X1_236 ( .A(_1101__bF_buf50), .B(_1135__bF_buf11_bF_buf3), .C(_3663__45_), .Y(_1442_) );
OAI21X1 OAI21X1_237 ( .A(_1204_), .B(_1134__bF_buf9), .C(_1442_), .Y(_309_) );
OAI21X1 OAI21X1_238 ( .A(_1101__bF_buf18), .B(_1135__bF_buf10_bF_buf3), .C(_3663__44_), .Y(_1443_) );
OAI21X1 OAI21X1_239 ( .A(_1206_), .B(_1134__bF_buf14), .C(_1443_), .Y(_310_) );
OAI21X1 OAI21X1_240 ( .A(_1101__bF_buf23), .B(_1135__bF_buf9_bF_buf0), .C(_3663__43_), .Y(_1444_) );
OAI21X1 OAI21X1_241 ( .A(_1208_), .B(_1134__bF_buf14), .C(_1444_), .Y(_311_) );
OAI21X1 OAI21X1_242 ( .A(_1101__bF_buf0), .B(_1135__bF_buf8_bF_buf1), .C(_3663__42_), .Y(_1445_) );
OAI21X1 OAI21X1_243 ( .A(_1210_), .B(_1134__bF_buf7), .C(_1445_), .Y(_312_) );
OAI21X1 OAI21X1_244 ( .A(_1101__bF_buf17), .B(_1135__bF_buf7_bF_buf3), .C(_3663__41_), .Y(_1446_) );
OAI21X1 OAI21X1_245 ( .A(_1212_), .B(_1134__bF_buf6), .C(_1446_), .Y(_313_) );
OAI21X1 OAI21X1_246 ( .A(_1101__bF_buf7), .B(_1135__bF_buf6_bF_buf0), .C(_3663__40_), .Y(_1447_) );
OAI21X1 OAI21X1_247 ( .A(_1214_), .B(_1134__bF_buf2), .C(_1447_), .Y(_314_) );
OAI21X1 OAI21X1_248 ( .A(_1101__bF_buf15), .B(_1135__bF_buf5_bF_buf2), .C(_3663__39_), .Y(_1448_) );
OAI21X1 OAI21X1_249 ( .A(_1216_), .B(_1134__bF_buf12), .C(_1448_), .Y(_315_) );
OAI21X1 OAI21X1_250 ( .A(_1101__bF_buf41), .B(_1135__bF_buf4_bF_buf2), .C(_3663__38_), .Y(_1449_) );
OAI21X1 OAI21X1_251 ( .A(_1218_), .B(_1134__bF_buf11), .C(_1449_), .Y(_316_) );
OAI21X1 OAI21X1_252 ( .A(_1101__bF_buf31), .B(_1135__bF_buf3_bF_buf2), .C(_3663__37_), .Y(_1450_) );
OAI21X1 OAI21X1_253 ( .A(_1220_), .B(_1134__bF_buf11), .C(_1450_), .Y(_317_) );
OAI21X1 OAI21X1_254 ( .A(_1101__bF_buf14), .B(_1135__bF_buf2_bF_buf0), .C(_3663__36_), .Y(_1451_) );
OAI21X1 OAI21X1_255 ( .A(_1222_), .B(_1134__bF_buf10), .C(_1451_), .Y(_318_) );
OAI21X1 OAI21X1_256 ( .A(_1101__bF_buf21), .B(_1135__bF_buf1_bF_buf2), .C(_3663__35_), .Y(_1452_) );
OAI21X1 OAI21X1_257 ( .A(_1224_), .B(_1134__bF_buf0), .C(_1452_), .Y(_319_) );
OAI21X1 OAI21X1_258 ( .A(_1101__bF_buf13), .B(_1135__bF_buf5), .C(_3663__34_), .Y(_1453_) );
OAI21X1 OAI21X1_259 ( .A(_1226_), .B(_1134__bF_buf9), .C(_1453_), .Y(_320_) );
OAI21X1 OAI21X1_260 ( .A(_1101__bF_buf15), .B(_1135__bF_buf14_bF_buf3), .C(_3663__33_), .Y(_1454_) );
OAI21X1 OAI21X1_261 ( .A(_1228_), .B(_1134__bF_buf12), .C(_1454_), .Y(_321_) );
OAI21X1 OAI21X1_262 ( .A(_1101__bF_buf28), .B(_1135__bF_buf13_bF_buf3), .C(_3663__32_), .Y(_1455_) );
OAI21X1 OAI21X1_263 ( .A(_1230_), .B(_1134__bF_buf7), .C(_1455_), .Y(_322_) );
OAI21X1 OAI21X1_264 ( .A(_1101__bF_buf6), .B(_1135__bF_buf12_bF_buf2), .C(_3663__31_), .Y(_1456_) );
OAI21X1 OAI21X1_265 ( .A(_1232_), .B(_1134__bF_buf1), .C(_1456_), .Y(_323_) );
OAI21X1 OAI21X1_266 ( .A(_1101__bF_buf28), .B(_1135__bF_buf11_bF_buf0), .C(_3663__30_), .Y(_1457_) );
OAI21X1 OAI21X1_267 ( .A(_1234_), .B(_1134__bF_buf7), .C(_1457_), .Y(_324_) );
OAI21X1 OAI21X1_268 ( .A(_1101__bF_buf7), .B(_1135__bF_buf10_bF_buf0), .C(_3663__29_), .Y(_1458_) );
OAI21X1 OAI21X1_269 ( .A(_1236_), .B(_1134__bF_buf2), .C(_1458_), .Y(_325_) );
OAI21X1 OAI21X1_270 ( .A(_1101__bF_buf34), .B(_1135__bF_buf9_bF_buf0), .C(_3663__28_), .Y(_1459_) );
OAI21X1 OAI21X1_271 ( .A(_1238_), .B(_1134__bF_buf13), .C(_1459_), .Y(_326_) );
OAI21X1 OAI21X1_272 ( .A(_1101__bF_buf31), .B(_1135__bF_buf8_bF_buf3), .C(_3663__27_), .Y(_1460_) );
OAI21X1 OAI21X1_273 ( .A(_1240_), .B(_1134__bF_buf11), .C(_1460_), .Y(_327_) );
OAI21X1 OAI21X1_274 ( .A(_1101__bF_buf29), .B(_1135__bF_buf7_bF_buf2), .C(_3663__26_), .Y(_1461_) );
OAI21X1 OAI21X1_275 ( .A(_1242_), .B(_1134__bF_buf14), .C(_1461_), .Y(_328_) );
OAI21X1 OAI21X1_276 ( .A(_1101__bF_buf42), .B(_1135__bF_buf6_bF_buf3), .C(_3663__25_), .Y(_1462_) );
OAI21X1 OAI21X1_277 ( .A(_1244_), .B(_1134__bF_buf10), .C(_1462_), .Y(_329_) );
OAI21X1 OAI21X1_278 ( .A(_1101__bF_buf39), .B(_1135__bF_buf5_bF_buf1), .C(_3663__24_), .Y(_1463_) );
OAI21X1 OAI21X1_279 ( .A(_1246_), .B(_1134__bF_buf6), .C(_1463_), .Y(_330_) );
OAI21X1 OAI21X1_280 ( .A(_1101__bF_buf55), .B(_1135__bF_buf4_bF_buf2), .C(_3663__23_), .Y(_1464_) );
OAI21X1 OAI21X1_281 ( .A(_1248_), .B(_1134__bF_buf5), .C(_1464_), .Y(_331_) );
OAI21X1 OAI21X1_282 ( .A(_1101__bF_buf51), .B(_1135__bF_buf3_bF_buf0), .C(_3663__22_), .Y(_1465_) );
OAI21X1 OAI21X1_283 ( .A(_1250_), .B(_1134__bF_buf2), .C(_1465_), .Y(_332_) );
OAI21X1 OAI21X1_284 ( .A(_1101__bF_buf46), .B(_1135__bF_buf2_bF_buf3), .C(_3663__21_), .Y(_1466_) );
OAI21X1 OAI21X1_285 ( .A(_1252_), .B(_1134__bF_buf5), .C(_1466_), .Y(_333_) );
OAI21X1 OAI21X1_286 ( .A(_1101__bF_buf13), .B(_1135__bF_buf1_bF_buf3), .C(_3663__20_), .Y(_1467_) );
OAI21X1 OAI21X1_287 ( .A(_1254_), .B(_1134__bF_buf2), .C(_1467_), .Y(_334_) );
OAI21X1 OAI21X1_288 ( .A(_1101__bF_buf20), .B(_1135__bF_buf4), .C(_3663__19_), .Y(_1468_) );
OAI21X1 OAI21X1_289 ( .A(_1256_), .B(_1134__bF_buf11), .C(_1468_), .Y(_335_) );
OAI21X1 OAI21X1_290 ( .A(_1101__bF_buf15), .B(_1135__bF_buf14_bF_buf3), .C(_3663__18_), .Y(_1469_) );
OAI21X1 OAI21X1_291 ( .A(_1258_), .B(_1134__bF_buf12), .C(_1469_), .Y(_336_) );
OAI21X1 OAI21X1_292 ( .A(_1101__bF_buf45), .B(_1135__bF_buf13_bF_buf2), .C(_3663__17_), .Y(_1470_) );
OAI21X1 OAI21X1_293 ( .A(_1260_), .B(_1134__bF_buf1), .C(_1470_), .Y(_337_) );
OAI21X1 OAI21X1_294 ( .A(_1101__bF_buf20), .B(_1135__bF_buf12_bF_buf3), .C(_3663__16_), .Y(_1471_) );
OAI21X1 OAI21X1_295 ( .A(_1262_), .B(_1134__bF_buf11), .C(_1471_), .Y(_338_) );
OAI21X1 OAI21X1_296 ( .A(_1101__bF_buf41), .B(_1135__bF_buf11_bF_buf3), .C(_3663__15_), .Y(_1472_) );
OAI21X1 OAI21X1_297 ( .A(_1264_), .B(_1134__bF_buf11), .C(_1472_), .Y(_339_) );
OAI21X1 OAI21X1_298 ( .A(_1101__bF_buf42), .B(_1135__bF_buf10_bF_buf0), .C(_3663__14_), .Y(_1473_) );
OAI21X1 OAI21X1_299 ( .A(_1266_), .B(_1134__bF_buf10), .C(_1473_), .Y(_340_) );
OAI21X1 OAI21X1_300 ( .A(_1101__bF_buf14), .B(_1135__bF_buf9_bF_buf2), .C(_3663__13_), .Y(_1474_) );
OAI21X1 OAI21X1_301 ( .A(_1268_), .B(_1134__bF_buf10), .C(_1474_), .Y(_341_) );
OAI21X1 OAI21X1_302 ( .A(_1101__bF_buf35), .B(_1135__bF_buf8_bF_buf0), .C(_3663__12_), .Y(_1475_) );
OAI21X1 OAI21X1_303 ( .A(_1270_), .B(_1134__bF_buf0), .C(_1475_), .Y(_342_) );
OAI21X1 OAI21X1_304 ( .A(_1101__bF_buf49), .B(_1135__bF_buf7_bF_buf0), .C(_3663__11_), .Y(_1476_) );
OAI21X1 OAI21X1_305 ( .A(_1272_), .B(_1134__bF_buf8), .C(_1476_), .Y(_343_) );
OAI21X1 OAI21X1_306 ( .A(_1101__bF_buf1), .B(_1135__bF_buf6_bF_buf0), .C(_3663__10_), .Y(_1477_) );
OAI21X1 OAI21X1_307 ( .A(_1274_), .B(_1134__bF_buf2), .C(_1477_), .Y(_344_) );
OAI21X1 OAI21X1_308 ( .A(_1101__bF_buf28), .B(_1135__bF_buf5_bF_buf3), .C(_3663__9_), .Y(_1478_) );
OAI21X1 OAI21X1_309 ( .A(_1276_), .B(_1134__bF_buf13), .C(_1478_), .Y(_345_) );
OAI21X1 OAI21X1_310 ( .A(_1101__bF_buf45), .B(_1135__bF_buf4_bF_buf0), .C(_3663__8_), .Y(_1479_) );
OAI21X1 OAI21X1_311 ( .A(_1278_), .B(_1134__bF_buf1), .C(_1479_), .Y(_346_) );
OAI21X1 OAI21X1_312 ( .A(_1101__bF_buf11), .B(_1135__bF_buf3_bF_buf2), .C(_3663__7_), .Y(_1480_) );
OAI21X1 OAI21X1_313 ( .A(_1280_), .B(_1134__bF_buf12), .C(_1480_), .Y(_347_) );
OAI21X1 OAI21X1_314 ( .A(_1101__bF_buf32), .B(_1135__bF_buf2_bF_buf3), .C(_3663__6_), .Y(_1481_) );
OAI21X1 OAI21X1_315 ( .A(_1282_), .B(_1134__bF_buf8), .C(_1481_), .Y(_348_) );
OAI21X1 OAI21X1_316 ( .A(_1101__bF_buf48), .B(_1135__bF_buf1_bF_buf0), .C(_3663__5_), .Y(_1482_) );
OAI21X1 OAI21X1_317 ( .A(_1284_), .B(_1134__bF_buf4), .C(_1482_), .Y(_349_) );
OAI21X1 OAI21X1_318 ( .A(_1101__bF_buf10), .B(_1135__bF_buf3), .C(_3663__4_), .Y(_1483_) );
OAI21X1 OAI21X1_319 ( .A(_1286_), .B(_1134__bF_buf5), .C(_1483_), .Y(_350_) );
OAI21X1 OAI21X1_320 ( .A(_1101__bF_buf5), .B(_1135__bF_buf14_bF_buf3), .C(_3663__3_), .Y(_1484_) );
OAI21X1 OAI21X1_321 ( .A(_1288_), .B(_1134__bF_buf5), .C(_1484_), .Y(_351_) );
OAI21X1 OAI21X1_322 ( .A(_1101__bF_buf0), .B(_1135__bF_buf13_bF_buf3), .C(_3663__2_), .Y(_1485_) );
OAI21X1 OAI21X1_323 ( .A(_1290_), .B(_1134__bF_buf13), .C(_1485_), .Y(_352_) );
OAI21X1 OAI21X1_324 ( .A(_1101__bF_buf45), .B(_1135__bF_buf12_bF_buf2), .C(_3663__1_), .Y(_1486_) );
OAI21X1 OAI21X1_325 ( .A(_1292_), .B(_1134__bF_buf1), .C(_1486_), .Y(_353_) );
OAI21X1 OAI21X1_326 ( .A(_1101__bF_buf40), .B(_1135__bF_buf11_bF_buf2), .C(_3663__0_), .Y(_1487_) );
OAI21X1 OAI21X1_327 ( .A(_1294_), .B(_1134__bF_buf0), .C(_1487_), .Y(_354_) );
INVX4 INVX4_1 ( .A(bundleStartMajId_i[63]), .Y(_1488_) );
NAND2X1 NAND2X1_72 ( .A(_3652__63_), .B(_1031__bF_buf67), .Y(_1489_) );
OAI21X1 OAI21X1_328 ( .A(_1488_), .B(_1031__bF_buf67), .C(_1489_), .Y(_355_) );
INVX2 INVX2_8 ( .A(bundleStartMajId_i[62]), .Y(_1490_) );
NAND2X1 NAND2X1_73 ( .A(_3652__62_), .B(_1031__bF_buf67), .Y(_1491_) );
OAI21X1 OAI21X1_329 ( .A(_1490_), .B(_1031__bF_buf67), .C(_1491_), .Y(_356_) );
INVX2 INVX2_9 ( .A(bundleStartMajId_i[61]), .Y(_1492_) );
NAND2X1 NAND2X1_74 ( .A(_3652__61_), .B(_1031__bF_buf23), .Y(_1493_) );
OAI21X1 OAI21X1_330 ( .A(_1031__bF_buf23), .B(_1492_), .C(_1493_), .Y(_357_) );
INVX2 INVX2_10 ( .A(bundleStartMajId_i[60]), .Y(_1494_) );
NAND2X1 NAND2X1_75 ( .A(_3652__60_), .B(_1031__bF_buf67), .Y(_1495_) );
OAI21X1 OAI21X1_331 ( .A(_1031__bF_buf67), .B(_1494_), .C(_1495_), .Y(_358_) );
INVX2 INVX2_11 ( .A(bundleStartMajId_i[59]), .Y(_1496_) );
NAND2X1 NAND2X1_76 ( .A(_3652__59_), .B(_1031__bF_buf61), .Y(_1497_) );
OAI21X1 OAI21X1_332 ( .A(_1031__bF_buf68), .B(_1496_), .C(_1497_), .Y(_359_) );
INVX2 INVX2_12 ( .A(bundleStartMajId_i[58]), .Y(_1498_) );
NAND2X1 NAND2X1_77 ( .A(_3652__58_), .B(_1031__bF_buf33), .Y(_1499_) );
OAI21X1 OAI21X1_333 ( .A(_1031__bF_buf33), .B(_1498_), .C(_1499_), .Y(_360_) );
INVX4 INVX4_2 ( .A(bundleStartMajId_i[57]), .Y(_1500_) );
NAND2X1 NAND2X1_78 ( .A(_3652__57_), .B(_1031__bF_buf33), .Y(_1501_) );
OAI21X1 OAI21X1_334 ( .A(_1031__bF_buf33), .B(_1500_), .C(_1501_), .Y(_361_) );
INVX2 INVX2_13 ( .A(bundleStartMajId_i[56]), .Y(_1502_) );
NAND2X1 NAND2X1_79 ( .A(_3652__56_), .B(_1031__bF_buf33), .Y(_1503_) );
OAI21X1 OAI21X1_335 ( .A(_1031__bF_buf33), .B(_1502_), .C(_1503_), .Y(_362_) );
INVX2 INVX2_14 ( .A(bundleStartMajId_i[55]), .Y(_1504_) );
NAND2X1 NAND2X1_80 ( .A(_3652__55_), .B(_1031__bF_buf1), .Y(_1505_) );
OAI21X1 OAI21X1_336 ( .A(_1031__bF_buf1), .B(_1504_), .C(_1505_), .Y(_363_) );
INVX4 INVX4_3 ( .A(bundleStartMajId_i[54]), .Y(_1506_) );
NAND2X1 NAND2X1_81 ( .A(_3652__54_), .B(_1031__bF_buf1), .Y(_1507_) );
OAI21X1 OAI21X1_337 ( .A(_1031__bF_buf1), .B(_1506_), .C(_1507_), .Y(_364_) );
INVX2 INVX2_15 ( .A(bundleStartMajId_i[53]), .Y(_1508_) );
NAND2X1 NAND2X1_82 ( .A(_3652__53_), .B(_1031__bF_buf0), .Y(_1509_) );
OAI21X1 OAI21X1_338 ( .A(_1031__bF_buf0), .B(_1508_), .C(_1509_), .Y(_365_) );
INVX4 INVX4_4 ( .A(bundleStartMajId_i[52]), .Y(_1510_) );
NAND2X1 NAND2X1_83 ( .A(_3652__52_), .B(_1031__bF_buf1), .Y(_1511_) );
OAI21X1 OAI21X1_339 ( .A(_1031__bF_buf1), .B(_1510_), .C(_1511_), .Y(_366_) );
INVX4 INVX4_5 ( .A(bundleStartMajId_i[51]), .Y(_1512_) );
NAND2X1 NAND2X1_84 ( .A(_3652__51_), .B(_1031__bF_buf30), .Y(_1513_) );
OAI21X1 OAI21X1_340 ( .A(_1031__bF_buf30), .B(_1512_), .C(_1513_), .Y(_367_) );
INVX1 INVX1_1 ( .A(bundleStartMajId_i[50]), .Y(_1514_) );
NAND2X1 NAND2X1_85 ( .A(_3652__50_), .B(_1031__bF_buf43), .Y(_1515_) );
OAI21X1 OAI21X1_341 ( .A(_1031__bF_buf43), .B(_1514_), .C(_1515_), .Y(_368_) );
INVX2 INVX2_16 ( .A(bundleStartMajId_i[49]), .Y(_1516_) );
NAND2X1 NAND2X1_86 ( .A(_3652__49_), .B(_1031__bF_buf53), .Y(_1517_) );
OAI21X1 OAI21X1_342 ( .A(_1031__bF_buf53), .B(_1516_), .C(_1517_), .Y(_369_) );
INVX4 INVX4_6 ( .A(bundleStartMajId_i[48]), .Y(_1518_) );
NAND2X1 NAND2X1_87 ( .A(_3652__48_), .B(_1031__bF_buf0), .Y(_1519_) );
OAI21X1 OAI21X1_343 ( .A(_1031__bF_buf0), .B(_1518_), .C(_1519_), .Y(_370_) );
INVX2 INVX2_17 ( .A(bundleStartMajId_i[47]), .Y(_1520_) );
NAND2X1 NAND2X1_88 ( .A(_3652__47_), .B(_1031__bF_buf33), .Y(_1521_) );
OAI21X1 OAI21X1_344 ( .A(_1031__bF_buf33), .B(_1520_), .C(_1521_), .Y(_371_) );
INVX4 INVX4_7 ( .A(bundleStartMajId_i[46]), .Y(_1522_) );
NAND2X1 NAND2X1_89 ( .A(_3652__46_), .B(_1031__bF_buf1), .Y(_1523_) );
OAI21X1 OAI21X1_345 ( .A(_1031__bF_buf1), .B(_1522_), .C(_1523_), .Y(_372_) );
INVX2 INVX2_18 ( .A(bundleStartMajId_i[45]), .Y(_1524_) );
NAND2X1 NAND2X1_90 ( .A(_3652__45_), .B(_1031__bF_buf37), .Y(_1525_) );
OAI21X1 OAI21X1_346 ( .A(_1031__bF_buf37), .B(_1524_), .C(_1525_), .Y(_373_) );
INVX2 INVX2_19 ( .A(bundleStartMajId_i[44]), .Y(_1526_) );
NAND2X1 NAND2X1_91 ( .A(_3652__44_), .B(_1031__bF_buf37), .Y(_1527_) );
OAI21X1 OAI21X1_347 ( .A(_1031__bF_buf69), .B(_1526_), .C(_1527_), .Y(_374_) );
INVX2 INVX2_20 ( .A(bundleStartMajId_i[43]), .Y(_1528_) );
NAND2X1 NAND2X1_92 ( .A(_3652__43_), .B(_1031__bF_buf5), .Y(_1529_) );
OAI21X1 OAI21X1_348 ( .A(_1031__bF_buf5), .B(_1528_), .C(_1529_), .Y(_375_) );
INVX4 INVX4_8 ( .A(bundleStartMajId_i[42]), .Y(_1530_) );
NAND2X1 NAND2X1_93 ( .A(_3652__42_), .B(_1031__bF_buf51), .Y(_1531_) );
OAI21X1 OAI21X1_349 ( .A(_1031__bF_buf51), .B(_1530_), .C(_1531_), .Y(_376_) );
INVX2 INVX2_21 ( .A(bundleStartMajId_i[41]), .Y(_1532_) );
NAND2X1 NAND2X1_94 ( .A(_3652__41_), .B(_1031__bF_buf5), .Y(_1533_) );
OAI21X1 OAI21X1_350 ( .A(_1031__bF_buf51), .B(_1532_), .C(_1533_), .Y(_377_) );
INVX4 INVX4_9 ( .A(bundleStartMajId_i[40]), .Y(_1534_) );
NAND2X1 NAND2X1_95 ( .A(_3652__40_), .B(_1031__bF_buf51), .Y(_1535_) );
OAI21X1 OAI21X1_351 ( .A(_1031__bF_buf51), .B(_1534_), .C(_1535_), .Y(_378_) );
INVX4 INVX4_10 ( .A(bundleStartMajId_i[39]), .Y(_1536_) );
NAND2X1 NAND2X1_96 ( .A(_3652__39_), .B(_1031__bF_buf55), .Y(_1537_) );
OAI21X1 OAI21X1_352 ( .A(_1031__bF_buf55), .B(_1536_), .C(_1537_), .Y(_379_) );
INVX4 INVX4_11 ( .A(bundleStartMajId_i[38]), .Y(_1538_) );
NAND2X1 NAND2X1_97 ( .A(_3652__38_), .B(_1031__bF_buf10), .Y(_1539_) );
OAI21X1 OAI21X1_353 ( .A(_1031__bF_buf10), .B(_1538_), .C(_1539_), .Y(_380_) );
INVX2 INVX2_22 ( .A(bundleStartMajId_i[37]), .Y(_1540_) );
NAND2X1 NAND2X1_98 ( .A(_3652__37_), .B(_1031__bF_buf10), .Y(_1541_) );
OAI21X1 OAI21X1_354 ( .A(_1031__bF_buf10), .B(_1540_), .C(_1541_), .Y(_381_) );
INVX4 INVX4_12 ( .A(bundleStartMajId_i[36]), .Y(_1542_) );
NAND2X1 NAND2X1_99 ( .A(_3652__36_), .B(_1031__bF_buf5), .Y(_1543_) );
OAI21X1 OAI21X1_355 ( .A(_1031__bF_buf69), .B(_1542_), .C(_1543_), .Y(_382_) );
INVX4 INVX4_13 ( .A(bundleStartMajId_i[35]), .Y(_1544_) );
NAND2X1 NAND2X1_100 ( .A(_3652__35_), .B(_1031__bF_buf55), .Y(_1545_) );
OAI21X1 OAI21X1_356 ( .A(_1031__bF_buf55), .B(_1544_), .C(_1545_), .Y(_383_) );
INVX4 INVX4_14 ( .A(bundleStartMajId_i[34]), .Y(_1546_) );
NAND2X1 NAND2X1_101 ( .A(_3652__34_), .B(_1031__bF_buf74), .Y(_1547_) );
OAI21X1 OAI21X1_357 ( .A(_1031__bF_buf74), .B(_1546_), .C(_1547_), .Y(_384_) );
INVX2 INVX2_23 ( .A(bundleStartMajId_i[33]), .Y(_1548_) );
NAND2X1 NAND2X1_102 ( .A(_3652__33_), .B(_1031__bF_buf69), .Y(_1549_) );
OAI21X1 OAI21X1_358 ( .A(_1031__bF_buf74), .B(_1548_), .C(_1549_), .Y(_385_) );
INVX2 INVX2_24 ( .A(bundleStartMajId_i[32]), .Y(_1550_) );
NAND2X1 NAND2X1_103 ( .A(_3652__32_), .B(_1031__bF_buf74), .Y(_1551_) );
OAI21X1 OAI21X1_359 ( .A(_1031__bF_buf74), .B(_1550_), .C(_1551_), .Y(_386_) );
INVX2 INVX2_25 ( .A(bundleStartMajId_i[31]), .Y(_1552_) );
NAND2X1 NAND2X1_104 ( .A(_3652__31_), .B(_1031__bF_buf42), .Y(_1553_) );
OAI21X1 OAI21X1_360 ( .A(_1031__bF_buf42), .B(_1552_), .C(_1553_), .Y(_387_) );
INVX4 INVX4_15 ( .A(bundleStartMajId_i[30]), .Y(_1554_) );
NAND2X1 NAND2X1_105 ( .A(_3652__30_), .B(_1031__bF_buf53), .Y(_1555_) );
OAI21X1 OAI21X1_361 ( .A(_1031__bF_buf15), .B(_1554_), .C(_1555_), .Y(_388_) );
INVX1 INVX1_2 ( .A(bundleStartMajId_i[29]), .Y(_1556_) );
NAND2X1 NAND2X1_106 ( .A(_3652__29_), .B(_1031__bF_buf53), .Y(_1557_) );
OAI21X1 OAI21X1_362 ( .A(_1031__bF_buf15), .B(_1556_), .C(_1557_), .Y(_389_) );
INVX4 INVX4_16 ( .A(bundleStartMajId_i[28]), .Y(_1558_) );
NAND2X1 NAND2X1_107 ( .A(_3652__28_), .B(_1031__bF_buf15), .Y(_1559_) );
OAI21X1 OAI21X1_363 ( .A(_1031__bF_buf51), .B(_1558_), .C(_1559_), .Y(_390_) );
INVX4 INVX4_17 ( .A(bundleStartMajId_i[27]), .Y(_1560_) );
NAND2X1 NAND2X1_108 ( .A(_3652__27_), .B(_1031__bF_buf37), .Y(_1561_) );
OAI21X1 OAI21X1_364 ( .A(_1031__bF_buf37), .B(_1560_), .C(_1561_), .Y(_391_) );
INVX2 INVX2_26 ( .A(bundleStartMajId_i[26]), .Y(_1562_) );
NAND2X1 NAND2X1_109 ( .A(_3652__26_), .B(_1031__bF_buf69), .Y(_1563_) );
OAI21X1 OAI21X1_365 ( .A(_1031__bF_buf69), .B(_1562_), .C(_1563_), .Y(_392_) );
INVX2 INVX2_27 ( .A(bundleStartMajId_i[25]), .Y(_1564_) );
NAND2X1 NAND2X1_110 ( .A(_3652__25_), .B(_1031__bF_buf37), .Y(_1565_) );
OAI21X1 OAI21X1_366 ( .A(_1031__bF_buf37), .B(_1564_), .C(_1565_), .Y(_393_) );
INVX4 INVX4_18 ( .A(bundleStartMajId_i[24]), .Y(_1566_) );
NAND2X1 NAND2X1_111 ( .A(_3652__24_), .B(_1031__bF_buf63), .Y(_1567_) );
OAI21X1 OAI21X1_367 ( .A(_1031__bF_buf42), .B(_1566_), .C(_1567_), .Y(_394_) );
INVX4 INVX4_19 ( .A(bundleStartMajId_i[23]), .Y(_1568_) );
NAND2X1 NAND2X1_112 ( .A(_3652__23_), .B(_1031__bF_buf23), .Y(_1569_) );
OAI21X1 OAI21X1_368 ( .A(_1031__bF_buf30), .B(_1568_), .C(_1569_), .Y(_395_) );
INVX4 INVX4_20 ( .A(bundleStartMajId_i[22]), .Y(_1570_) );
NAND2X1 NAND2X1_113 ( .A(_3652__22_), .B(_1031__bF_buf26), .Y(_1571_) );
OAI21X1 OAI21X1_369 ( .A(_1031__bF_buf26), .B(_1570_), .C(_1571_), .Y(_396_) );
INVX2 INVX2_28 ( .A(bundleStartMajId_i[21]), .Y(_1572_) );
NAND2X1 NAND2X1_114 ( .A(_3652__21_), .B(_1031__bF_buf16), .Y(_1573_) );
OAI21X1 OAI21X1_370 ( .A(_1031__bF_buf63), .B(_1572_), .C(_1573_), .Y(_397_) );
INVX4 INVX4_21 ( .A(bundleStartMajId_i[20]), .Y(_1574_) );
NAND2X1 NAND2X1_115 ( .A(_3652__20_), .B(_1031__bF_buf63), .Y(_1575_) );
OAI21X1 OAI21X1_371 ( .A(_1031__bF_buf63), .B(_1574_), .C(_1575_), .Y(_398_) );
INVX2 INVX2_29 ( .A(bundleStartMajId_i[19]), .Y(_1576_) );
NAND2X1 NAND2X1_116 ( .A(_3652__19_), .B(_1031__bF_buf16), .Y(_1577_) );
OAI21X1 OAI21X1_372 ( .A(_1031__bF_buf16), .B(_1576_), .C(_1577_), .Y(_399_) );
INVX2 INVX2_30 ( .A(bundleStartMajId_i[18]), .Y(_1578_) );
NAND2X1 NAND2X1_117 ( .A(_3652__18_), .B(_1031__bF_buf43), .Y(_1579_) );
OAI21X1 OAI21X1_373 ( .A(_1031__bF_buf43), .B(_1578_), .C(_1579_), .Y(_400_) );
INVX2 INVX2_31 ( .A(bundleStartMajId_i[17]), .Y(_1580_) );
NAND2X1 NAND2X1_118 ( .A(_3652__17_), .B(_1031__bF_buf30), .Y(_1581_) );
OAI21X1 OAI21X1_374 ( .A(_1031__bF_buf30), .B(_1580_), .C(_1581_), .Y(_401_) );
INVX2 INVX2_32 ( .A(bundleStartMajId_i[16]), .Y(_1582_) );
NAND2X1 NAND2X1_119 ( .A(_3652__16_), .B(_1031__bF_buf26), .Y(_1583_) );
OAI21X1 OAI21X1_375 ( .A(_1031__bF_buf26), .B(_1582_), .C(_1583_), .Y(_402_) );
INVX4 INVX4_22 ( .A(bundleStartMajId_i[15]), .Y(_1584_) );
NAND2X1 NAND2X1_120 ( .A(_3652__15_), .B(_1031__bF_buf43), .Y(_1585_) );
OAI21X1 OAI21X1_376 ( .A(_1031__bF_buf43), .B(_1584_), .C(_1585_), .Y(_403_) );
INVX4 INVX4_23 ( .A(bundleStartMajId_i[14]), .Y(_1586_) );
NAND2X1 NAND2X1_121 ( .A(_3652__14_), .B(_1031__bF_buf65), .Y(_1587_) );
OAI21X1 OAI21X1_377 ( .A(_1031__bF_buf65), .B(_1586_), .C(_1587_), .Y(_404_) );
INVX2 INVX2_33 ( .A(bundleStartMajId_i[13]), .Y(_1588_) );
NAND2X1 NAND2X1_122 ( .A(_3652__13_), .B(_1031__bF_buf65), .Y(_1589_) );
OAI21X1 OAI21X1_378 ( .A(_1031__bF_buf65), .B(_1588_), .C(_1589_), .Y(_405_) );
INVX2 INVX2_34 ( .A(bundleStartMajId_i[12]), .Y(_1590_) );
NAND2X1 NAND2X1_123 ( .A(_3652__12_), .B(_1031__bF_buf65), .Y(_1591_) );
OAI21X1 OAI21X1_379 ( .A(_1031__bF_buf65), .B(_1590_), .C(_1591_), .Y(_406_) );
INVX2 INVX2_35 ( .A(bundleStartMajId_i[11]), .Y(_1592_) );
NAND2X1 NAND2X1_124 ( .A(_3652__11_), .B(_1031__bF_buf30), .Y(_1593_) );
OAI21X1 OAI21X1_380 ( .A(_1031__bF_buf16), .B(_1592_), .C(_1593_), .Y(_407_) );
INVX4 INVX4_24 ( .A(bundleStartMajId_i[10]), .Y(_1594_) );
NAND2X1 NAND2X1_125 ( .A(_3652__10_), .B(_1031__bF_buf63), .Y(_1595_) );
OAI21X1 OAI21X1_381 ( .A(_1031__bF_buf63), .B(_1594_), .C(_1595_), .Y(_408_) );
INVX1 INVX1_3 ( .A(bundleStartMajId_i[9]), .Y(_1596_) );
NAND2X1 NAND2X1_126 ( .A(_3652__9_), .B(_1031__bF_buf42), .Y(_1597_) );
OAI21X1 OAI21X1_382 ( .A(_1031__bF_buf42), .B(_1596_), .C(_1597_), .Y(_409_) );
INVX2 INVX2_36 ( .A(bundleStartMajId_i[8]), .Y(_1598_) );
NAND2X1 NAND2X1_127 ( .A(_3652__8_), .B(_1031__bF_buf53), .Y(_1599_) );
OAI21X1 OAI21X1_383 ( .A(_1031__bF_buf53), .B(_1598_), .C(_1599_), .Y(_410_) );
INVX2 INVX2_37 ( .A(bundleStartMajId_i[7]), .Y(_1600_) );
NAND2X1 NAND2X1_128 ( .A(_3652__7_), .B(_1031__bF_buf69), .Y(_1601_) );
OAI21X1 OAI21X1_384 ( .A(_1031__bF_buf69), .B(_1600_), .C(_1601_), .Y(_411_) );
INVX4 INVX4_25 ( .A(bundleStartMajId_i[6]), .Y(_1602_) );
NAND2X1 NAND2X1_129 ( .A(_3652__6_), .B(_1031__bF_buf32), .Y(_1603_) );
OAI21X1 OAI21X1_385 ( .A(_1031__bF_buf32), .B(_1602_), .C(_1603_), .Y(_412_) );
INVX4 INVX4_26 ( .A(bundleStartMajId_i[5]), .Y(_1604_) );
NAND2X1 NAND2X1_130 ( .A(_3652__5_), .B(_1031__bF_buf60), .Y(_1605_) );
OAI21X1 OAI21X1_386 ( .A(_1031__bF_buf60), .B(_1604_), .C(_1605_), .Y(_413_) );
INVX1 INVX1_4 ( .A(bundleStartMajId_i[4]), .Y(_1606_) );
NAND2X1 NAND2X1_131 ( .A(_3652__4_), .B(_1031__bF_buf72), .Y(_1607_) );
OAI21X1 OAI21X1_387 ( .A(_1031__bF_buf72), .B(_1606_), .C(_1607_), .Y(_414_) );
INVX2 INVX2_38 ( .A(bundleStartMajId_i[3]), .Y(_1608_) );
NAND2X1 NAND2X1_132 ( .A(_3652__3_), .B(_1031__bF_buf37), .Y(_1609_) );
OAI21X1 OAI21X1_388 ( .A(_1031__bF_buf37), .B(_1608_), .C(_1609_), .Y(_415_) );
INVX4 INVX4_27 ( .A(bundleStartMajId_i[2]), .Y(_1610_) );
NAND2X1 NAND2X1_133 ( .A(_3652__2_), .B(_1031__bF_buf51), .Y(_1611_) );
OAI21X1 OAI21X1_389 ( .A(_1031__bF_buf15), .B(_1610_), .C(_1611_), .Y(_416_) );
INVX1 INVX1_5 ( .A(bundleStartMajId_i[1]), .Y(_1612_) );
NAND2X1 NAND2X1_134 ( .A(_3652__1_), .B(_1031__bF_buf32), .Y(_1613_) );
OAI21X1 OAI21X1_390 ( .A(_1031__bF_buf32), .B(_1612_), .C(_1613_), .Y(_417_) );
INVX2 INVX2_39 ( .A(bundleStartMajId_i[0]), .Y(_1614_) );
NAND2X1 NAND2X1_135 ( .A(_3652__0_), .B(_1031__bF_buf15), .Y(_1615_) );
OAI21X1 OAI21X1_391 ( .A(_1031__bF_buf42), .B(_1614_), .C(_1615_), .Y(_418_) );
NAND2X1 NAND2X1_136 ( .A(_3653__63_), .B(_1039__bF_buf0), .Y(_1616_) );
OAI21X1 OAI21X1_392 ( .A(bundleStartMajId_i[63]), .B(_1039__bF_buf0), .C(_1616_), .Y(_419_) );
INVX1 INVX1_6 ( .A(_3653__62_), .Y(_1617_) );
INVX8 INVX8_1 ( .A(_1039__bF_buf25), .Y(_611_) );
NAND2X1 NAND2X1_137 ( .A(bundleStartMajId_i[63]), .B(bundleStartMajId_i[62]), .Y(_1618_) );
INVX1 INVX1_7 ( .A(_1618_), .Y(_1619_) );
NOR2X1 NOR2X1_1 ( .A(bundleStartMajId_i[63]), .B(bundleStartMajId_i[62]), .Y(_1620_) );
NOR2X1 NOR2X1_2 ( .A(_1620_), .B(_1619_), .Y(_1621_) );
NAND2X1 NAND2X1_138 ( .A(_611__bF_buf1), .B(_1621_), .Y(_1622_) );
OAI21X1 OAI21X1_393 ( .A(_1617_), .B(_611__bF_buf1), .C(_1622_), .Y(_420_) );
NAND2X1 NAND2X1_139 ( .A(bundleStartMajId_i[62]), .B(bundleStartMajId_i[61]), .Y(_1623_) );
OAI21X1 OAI21X1_394 ( .A(_1488_), .B(_1490_), .C(_1492_), .Y(_1624_) );
OAI21X1 OAI21X1_395 ( .A(_1488_), .B(_1623_), .C(_1624_), .Y(_1625_) );
NAND2X1 NAND2X1_140 ( .A(_3653__61_), .B(_1039__bF_buf57), .Y(_1626_) );
OAI21X1 OAI21X1_396 ( .A(_1625_), .B(_1039__bF_buf57), .C(_1626_), .Y(_421_) );
NAND2X1 NAND2X1_141 ( .A(bundleStartMajId_i[61]), .B(bundleStartMajId_i[60]), .Y(_1627_) );
OAI21X1 OAI21X1_397 ( .A(_1623_), .B(_1488_), .C(_1494_), .Y(_1628_) );
OAI21X1 OAI21X1_398 ( .A(_1618_), .B(_1627_), .C(_1628_), .Y(_1629_) );
NAND2X1 NAND2X1_142 ( .A(_3653__60_), .B(_1039__bF_buf15), .Y(_1630_) );
OAI21X1 OAI21X1_399 ( .A(_1629_), .B(_1039__bF_buf15), .C(_1630_), .Y(_422_) );
NOR2X1 NOR2X1_3 ( .A(_1618_), .B(_1627_), .Y(_1631_) );
NAND2X1 NAND2X1_143 ( .A(bundleStartMajId_i[59]), .B(_1631_), .Y(_1632_) );
INVX1 INVX1_8 ( .A(_1632_), .Y(_1633_) );
OAI21X1 OAI21X1_400 ( .A(_1631_), .B(bundleStartMajId_i[59]), .C(_611__bF_buf1), .Y(_1634_) );
NAND2X1 NAND2X1_144 ( .A(_3653__59_), .B(_1039__bF_buf38), .Y(_1635_) );
OAI21X1 OAI21X1_401 ( .A(_1633_), .B(_1634_), .C(_1635_), .Y(_423_) );
INVX2 INVX2_40 ( .A(_1631_), .Y(_1636_) );
NAND2X1 NAND2X1_145 ( .A(bundleStartMajId_i[59]), .B(bundleStartMajId_i[58]), .Y(_1637_) );
OAI21X1 OAI21X1_402 ( .A(_1636_), .B(_1496_), .C(_1498_), .Y(_1638_) );
OAI21X1 OAI21X1_403 ( .A(_1636_), .B(_1637_), .C(_1638_), .Y(_1639_) );
NAND2X1 NAND2X1_146 ( .A(_3653__58_), .B(_1039__bF_buf15), .Y(_1640_) );
OAI21X1 OAI21X1_404 ( .A(_1639_), .B(_1039__bF_buf15), .C(_1640_), .Y(_424_) );
NAND2X1 NAND2X1_147 ( .A(bundleStartMajId_i[58]), .B(bundleStartMajId_i[57]), .Y(_1641_) );
OAI21X1 OAI21X1_405 ( .A(_1636_), .B(_1637_), .C(_1500_), .Y(_1642_) );
OAI21X1 OAI21X1_406 ( .A(_1632_), .B(_1641_), .C(_1642_), .Y(_1643_) );
NAND2X1 NAND2X1_148 ( .A(_3653__57_), .B(_1039__bF_buf38), .Y(_1644_) );
OAI21X1 OAI21X1_407 ( .A(_1643_), .B(_1039__bF_buf38), .C(_1644_), .Y(_425_) );
OAI21X1 OAI21X1_408 ( .A(_1632_), .B(_1641_), .C(_1502_), .Y(_1645_) );
NAND2X1 NAND2X1_149 ( .A(bundleStartMajId_i[57]), .B(bundleStartMajId_i[56]), .Y(_1646_) );
NOR2X1 NOR2X1_4 ( .A(_1637_), .B(_1646_), .Y(_1647_) );
NAND2X1 NAND2X1_150 ( .A(_1631_), .B(_1647_), .Y(_1648_) );
NAND2X1 NAND2X1_151 ( .A(_1648_), .B(_1645_), .Y(_1649_) );
NAND2X1 NAND2X1_152 ( .A(_3653__56_), .B(_1039__bF_buf38), .Y(_1650_) );
OAI21X1 OAI21X1_409 ( .A(_1649_), .B(_1039__bF_buf38), .C(_1650_), .Y(_426_) );
NOR2X1 NOR2X1_5 ( .A(_1504_), .B(_1648_), .Y(_1651_) );
AND2X2 AND2X2_1 ( .A(_1631_), .B(_1647_), .Y(_1652_) );
OAI21X1 OAI21X1_410 ( .A(_1652_), .B(bundleStartMajId_i[55]), .C(_611__bF_buf1), .Y(_1653_) );
NAND2X1 NAND2X1_153 ( .A(_3653__55_), .B(_1039__bF_buf56), .Y(_1654_) );
OAI21X1 OAI21X1_411 ( .A(_1653_), .B(_1651_), .C(_1654_), .Y(_427_) );
XNOR2X1 XNOR2X1_1 ( .A(_1651_), .B(bundleStartMajId_i[54]), .Y(_1655_) );
NAND2X1 NAND2X1_154 ( .A(_3653__54_), .B(_1039__bF_buf56), .Y(_1656_) );
OAI21X1 OAI21X1_412 ( .A(_1655_), .B(_1039__bF_buf22), .C(_1656_), .Y(_428_) );
INVX2 INVX2_41 ( .A(_1651_), .Y(_1657_) );
OAI21X1 OAI21X1_413 ( .A(_1657_), .B(_1506_), .C(_1508_), .Y(_1658_) );
NAND2X1 NAND2X1_155 ( .A(bundleStartMajId_i[54]), .B(bundleStartMajId_i[53]), .Y(_1659_) );
OAI21X1 OAI21X1_414 ( .A(_1657_), .B(_1659_), .C(_1658_), .Y(_1660_) );
NAND2X1 NAND2X1_156 ( .A(_3653__53_), .B(_1039__bF_buf56), .Y(_1661_) );
OAI21X1 OAI21X1_415 ( .A(_1660_), .B(_1039__bF_buf56), .C(_1661_), .Y(_429_) );
INVX1 INVX1_9 ( .A(_1659_), .Y(_1662_) );
NAND2X1 NAND2X1_157 ( .A(_1662_), .B(_1651_), .Y(_1663_) );
XNOR2X1 XNOR2X1_2 ( .A(_1663_), .B(_1510_), .Y(_1664_) );
NAND2X1 NAND2X1_158 ( .A(_3653__52_), .B(_1039__bF_buf12), .Y(_1665_) );
OAI21X1 OAI21X1_416 ( .A(_1664_), .B(_1039__bF_buf12), .C(_1665_), .Y(_430_) );
OAI21X1 OAI21X1_417 ( .A(_1663_), .B(_1510_), .C(_1512_), .Y(_1666_) );
NAND2X1 NAND2X1_159 ( .A(bundleStartMajId_i[52]), .B(bundleStartMajId_i[51]), .Y(_1667_) );
OR2X2 OR2X2_1 ( .A(_1659_), .B(_1667_), .Y(_1668_) );
OAI21X1 OAI21X1_418 ( .A(_1657_), .B(_1668_), .C(_1666_), .Y(_1669_) );
NAND2X1 NAND2X1_160 ( .A(_3653__51_), .B(_1039__bF_buf56), .Y(_1670_) );
OAI21X1 OAI21X1_419 ( .A(_1669_), .B(_1039__bF_buf56), .C(_1670_), .Y(_431_) );
NOR2X1 NOR2X1_6 ( .A(_1668_), .B(_1657_), .Y(_1671_) );
XNOR2X1 XNOR2X1_3 ( .A(_1671_), .B(bundleStartMajId_i[50]), .Y(_1672_) );
NAND2X1 NAND2X1_161 ( .A(_3653__50_), .B(_1039__bF_buf12), .Y(_1673_) );
OAI21X1 OAI21X1_420 ( .A(_1672_), .B(_1039__bF_buf12), .C(_1673_), .Y(_432_) );
NAND2X1 NAND2X1_162 ( .A(bundleStartMajId_i[55]), .B(bundleStartMajId_i[52]), .Y(_1674_) );
NOR2X1 NOR2X1_7 ( .A(_1659_), .B(_1674_), .Y(_1675_) );
NOR2X1 NOR2X1_8 ( .A(_1512_), .B(_1514_), .Y(_1676_) );
NAND3X1 NAND3X1_1 ( .A(_1675_), .B(_1676_), .C(_1652_), .Y(_1677_) );
XNOR2X1 XNOR2X1_4 ( .A(_1677_), .B(_1516_), .Y(_1678_) );
NAND2X1 NAND2X1_163 ( .A(_3653__49_), .B(_1039__bF_buf22), .Y(_1679_) );
OAI21X1 OAI21X1_421 ( .A(_1678_), .B(_1039__bF_buf22), .C(_1679_), .Y(_433_) );
NAND2X1 NAND2X1_164 ( .A(_3653__48_), .B(_1039__bF_buf22), .Y(_1680_) );
NOR2X1 NOR2X1_9 ( .A(_1516_), .B(_1677_), .Y(_1681_) );
XNOR2X1 XNOR2X1_5 ( .A(_1681_), .B(bundleStartMajId_i[48]), .Y(_1682_) );
OAI21X1 OAI21X1_422 ( .A(_1682_), .B(_1039__bF_buf22), .C(_1680_), .Y(_434_) );
NAND2X1 NAND2X1_165 ( .A(bundleStartMajId_i[51]), .B(bundleStartMajId_i[48]), .Y(_1683_) );
NAND2X1 NAND2X1_166 ( .A(bundleStartMajId_i[50]), .B(bundleStartMajId_i[49]), .Y(_1684_) );
NOR2X1 NOR2X1_10 ( .A(_1683_), .B(_1684_), .Y(_1685_) );
NAND2X1 NAND2X1_167 ( .A(_1675_), .B(_1685_), .Y(_1686_) );
NOR2X1 NOR2X1_11 ( .A(_1648_), .B(_1686_), .Y(_1687_) );
NAND2X1 NAND2X1_168 ( .A(bundleStartMajId_i[47]), .B(_1687_), .Y(_1688_) );
INVX1 INVX1_10 ( .A(_1688_), .Y(_1689_) );
OAI21X1 OAI21X1_423 ( .A(_1687_), .B(bundleStartMajId_i[47]), .C(_611__bF_buf0), .Y(_1690_) );
NAND2X1 NAND2X1_169 ( .A(_3653__47_), .B(_1039__bF_buf1), .Y(_1691_) );
OAI21X1 OAI21X1_424 ( .A(_1689_), .B(_1690_), .C(_1691_), .Y(_435_) );
XNOR2X1 XNOR2X1_6 ( .A(_1688_), .B(_1522_), .Y(_1692_) );
NAND2X1 NAND2X1_170 ( .A(_3653__46_), .B(_1039__bF_buf1), .Y(_1693_) );
OAI21X1 OAI21X1_425 ( .A(_1692_), .B(_1039__bF_buf16), .C(_1693_), .Y(_436_) );
NAND2X1 NAND2X1_171 ( .A(bundleStartMajId_i[46]), .B(bundleStartMajId_i[45]), .Y(_1694_) );
NOR2X1 NOR2X1_12 ( .A(_1694_), .B(_1688_), .Y(_1695_) );
OAI21X1 OAI21X1_426 ( .A(_1688_), .B(_1522_), .C(_1524_), .Y(_1696_) );
NAND2X1 NAND2X1_172 ( .A(_611__bF_buf0), .B(_1696_), .Y(_1697_) );
NAND2X1 NAND2X1_173 ( .A(_3653__45_), .B(_1039__bF_buf1), .Y(_1698_) );
OAI21X1 OAI21X1_427 ( .A(_1697_), .B(_1695_), .C(_1698_), .Y(_437_) );
OAI21X1 OAI21X1_428 ( .A(_1688_), .B(_1694_), .C(_1526_), .Y(_1699_) );
NAND2X1 NAND2X1_174 ( .A(bundleStartMajId_i[44]), .B(_1695_), .Y(_1700_) );
NAND2X1 NAND2X1_175 ( .A(_1699_), .B(_1700_), .Y(_1701_) );
NAND2X1 NAND2X1_176 ( .A(_3653__44_), .B(_1039__bF_buf13), .Y(_1702_) );
OAI21X1 OAI21X1_429 ( .A(_1701_), .B(_1039__bF_buf13), .C(_1702_), .Y(_438_) );
NAND2X1 NAND2X1_177 ( .A(_1528_), .B(_1700_), .Y(_1703_) );
NAND2X1 NAND2X1_178 ( .A(bundleStartMajId_i[44]), .B(bundleStartMajId_i[43]), .Y(_1704_) );
OR2X2 OR2X2_2 ( .A(_1694_), .B(_1704_), .Y(_1705_) );
OAI21X1 OAI21X1_430 ( .A(_1688_), .B(_1705_), .C(_1703_), .Y(_1706_) );
NAND2X1 NAND2X1_179 ( .A(_3653__43_), .B(_1039__bF_buf43), .Y(_1707_) );
OAI21X1 OAI21X1_431 ( .A(_1706_), .B(_1039__bF_buf43), .C(_1707_), .Y(_439_) );
NOR2X1 NOR2X1_13 ( .A(_1705_), .B(_1688_), .Y(_1708_) );
XNOR2X1 XNOR2X1_7 ( .A(_1708_), .B(bundleStartMajId_i[42]), .Y(_1709_) );
NAND2X1 NAND2X1_180 ( .A(_3653__42_), .B(_1039__bF_buf1), .Y(_1710_) );
OAI21X1 OAI21X1_432 ( .A(_1709_), .B(_1039__bF_buf1), .C(_1710_), .Y(_440_) );
AND2X2 AND2X2_2 ( .A(_1675_), .B(_1685_), .Y(_1711_) );
NAND2X1 NAND2X1_181 ( .A(_1711_), .B(_1652_), .Y(_1712_) );
NAND2X1 NAND2X1_182 ( .A(bundleStartMajId_i[47]), .B(bundleStartMajId_i[44]), .Y(_1713_) );
OR2X2 OR2X2_3 ( .A(_1694_), .B(_1713_), .Y(_1714_) );
NOR2X1 NOR2X1_14 ( .A(_1714_), .B(_1712_), .Y(_1715_) );
NOR2X1 NOR2X1_15 ( .A(_1528_), .B(_1530_), .Y(_1716_) );
AND2X2 AND2X2_3 ( .A(_1715_), .B(_1716_), .Y(_1717_) );
XNOR2X1 XNOR2X1_8 ( .A(_1717_), .B(bundleStartMajId_i[41]), .Y(_1718_) );
NAND2X1 NAND2X1_183 ( .A(_3653__41_), .B(_1039__bF_buf43), .Y(_1719_) );
OAI21X1 OAI21X1_433 ( .A(_1718_), .B(_1039__bF_buf43), .C(_1719_), .Y(_441_) );
NAND2X1 NAND2X1_184 ( .A(_3653__40_), .B(_1039__bF_buf4), .Y(_1720_) );
NAND2X1 NAND2X1_185 ( .A(bundleStartMajId_i[41]), .B(_1717_), .Y(_1721_) );
XNOR2X1 XNOR2X1_9 ( .A(_1721_), .B(_1534_), .Y(_1722_) );
OAI21X1 OAI21X1_434 ( .A(_1722_), .B(_1039__bF_buf43), .C(_1720_), .Y(_442_) );
AND2X2 AND2X2_4 ( .A(bundleStartMajId_i[43]), .B(bundleStartMajId_i[40]), .Y(_1723_) );
AND2X2 AND2X2_5 ( .A(bundleStartMajId_i[42]), .B(bundleStartMajId_i[41]), .Y(_1724_) );
NAND2X1 NAND2X1_186 ( .A(_1723_), .B(_1724_), .Y(_1725_) );
NOR2X1 NOR2X1_16 ( .A(_1725_), .B(_1714_), .Y(_1726_) );
NAND2X1 NAND2X1_187 ( .A(_1726_), .B(_1687_), .Y(_1727_) );
NOR2X1 NOR2X1_17 ( .A(_1536_), .B(_1727_), .Y(_1728_) );
INVX1 INVX1_11 ( .A(_1727_), .Y(_1729_) );
OAI21X1 OAI21X1_435 ( .A(_1729_), .B(bundleStartMajId_i[39]), .C(_611__bF_buf0), .Y(_1730_) );
NAND2X1 NAND2X1_188 ( .A(_3653__39_), .B(_1039__bF_buf23), .Y(_1731_) );
OAI21X1 OAI21X1_436 ( .A(_1730_), .B(_1728_), .C(_1731_), .Y(_443_) );
XNOR2X1 XNOR2X1_10 ( .A(_1728_), .B(bundleStartMajId_i[38]), .Y(_1732_) );
NAND2X1 NAND2X1_189 ( .A(_3653__38_), .B(_1039__bF_buf28), .Y(_1733_) );
OAI21X1 OAI21X1_437 ( .A(_1732_), .B(_1039__bF_buf28), .C(_1733_), .Y(_444_) );
NOR2X1 NOR2X1_18 ( .A(_1536_), .B(_1538_), .Y(_1734_) );
NAND3X1 NAND3X1_2 ( .A(bundleStartMajId_i[37]), .B(_1734_), .C(_1729_), .Y(_1735_) );
INVX1 INVX1_12 ( .A(_1734_), .Y(_1736_) );
OAI21X1 OAI21X1_438 ( .A(_1727_), .B(_1736_), .C(_1540_), .Y(_1737_) );
NAND2X1 NAND2X1_190 ( .A(_1737_), .B(_1735_), .Y(_1738_) );
NAND2X1 NAND2X1_191 ( .A(_3653__37_), .B(_1039__bF_buf23), .Y(_1739_) );
OAI21X1 OAI21X1_439 ( .A(_1738_), .B(_1039__bF_buf23), .C(_1739_), .Y(_445_) );
NAND2X1 NAND2X1_192 ( .A(bundleStartMajId_i[38]), .B(bundleStartMajId_i[37]), .Y(_1740_) );
INVX2 INVX2_42 ( .A(_1740_), .Y(_1741_) );
AOI21X1 AOI21X1_1 ( .A(_1741_), .B(_1728_), .C(bundleStartMajId_i[36]), .Y(_1742_) );
OAI21X1 OAI21X1_440 ( .A(_1735_), .B(_1542_), .C(_611__bF_buf0), .Y(_1743_) );
NAND2X1 NAND2X1_193 ( .A(_3653__36_), .B(_1039__bF_buf23), .Y(_1744_) );
OAI21X1 OAI21X1_441 ( .A(_1743_), .B(_1742_), .C(_1744_), .Y(_446_) );
NAND2X1 NAND2X1_194 ( .A(bundleStartMajId_i[36]), .B(bundleStartMajId_i[35]), .Y(_1745_) );
NOR2X1 NOR2X1_19 ( .A(_1740_), .B(_1745_), .Y(_1746_) );
NAND2X1 NAND2X1_195 ( .A(_1746_), .B(_1728_), .Y(_1747_) );
OAI21X1 OAI21X1_442 ( .A(_1735_), .B(_1542_), .C(_1544_), .Y(_1748_) );
NAND2X1 NAND2X1_196 ( .A(_1747_), .B(_1748_), .Y(_1749_) );
NAND2X1 NAND2X1_197 ( .A(_3653__35_), .B(_1039__bF_buf23), .Y(_1750_) );
OAI21X1 OAI21X1_443 ( .A(_1749_), .B(_1039__bF_buf23), .C(_1750_), .Y(_447_) );
XNOR2X1 XNOR2X1_11 ( .A(_1747_), .B(_1546_), .Y(_1751_) );
NAND2X1 NAND2X1_198 ( .A(_3653__34_), .B(_1039__bF_buf23), .Y(_1752_) );
OAI21X1 OAI21X1_444 ( .A(_1751_), .B(_1039__bF_buf23), .C(_1752_), .Y(_448_) );
NAND2X1 NAND2X1_199 ( .A(bundleStartMajId_i[39]), .B(bundleStartMajId_i[36]), .Y(_1753_) );
OR2X2 OR2X2_4 ( .A(_1740_), .B(_1753_), .Y(_1754_) );
NOR2X1 NOR2X1_20 ( .A(_1544_), .B(_1546_), .Y(_1755_) );
INVX1 INVX1_13 ( .A(_1755_), .Y(_1756_) );
NOR3X1 NOR3X1_1 ( .A(_1754_), .B(_1756_), .C(_1727_), .Y(_1757_) );
XNOR2X1 XNOR2X1_12 ( .A(_1757_), .B(bundleStartMajId_i[33]), .Y(_1758_) );
NAND2X1 NAND2X1_200 ( .A(_3653__33_), .B(_1039__bF_buf28), .Y(_1759_) );
OAI21X1 OAI21X1_445 ( .A(_1758_), .B(_1039__bF_buf28), .C(_1759_), .Y(_449_) );
INVX1 INVX1_14 ( .A(_3653__32_), .Y(_1760_) );
AOI21X1 AOI21X1_2 ( .A(bundleStartMajId_i[33]), .B(_1757_), .C(_1550_), .Y(_1761_) );
NAND2X1 NAND2X1_201 ( .A(bundleStartMajId_i[33]), .B(_1757_), .Y(_1762_) );
NOR2X1 NOR2X1_21 ( .A(bundleStartMajId_i[32]), .B(_1762_), .Y(_1763_) );
OAI21X1 OAI21X1_446 ( .A(_1763_), .B(_1761_), .C(_611__bF_buf0), .Y(_1764_) );
OAI21X1 OAI21X1_447 ( .A(_1760_), .B(_611__bF_buf0), .C(_1764_), .Y(_450_) );
AND2X2 AND2X2_6 ( .A(bundleStartMajId_i[34]), .B(bundleStartMajId_i[33]), .Y(_1765_) );
NAND3X1 NAND3X1_3 ( .A(bundleStartMajId_i[35]), .B(bundleStartMajId_i[32]), .C(_1765_), .Y(_1766_) );
NOR2X1 NOR2X1_22 ( .A(_1754_), .B(_1766_), .Y(_1767_) );
NAND2X1 NAND2X1_202 ( .A(_1726_), .B(_1767_), .Y(_1768_) );
NOR2X1 NOR2X1_23 ( .A(_1712_), .B(_1768_), .Y(_1769_) );
NAND2X1 NAND2X1_203 ( .A(bundleStartMajId_i[31]), .B(_1769_), .Y(_1770_) );
INVX1 INVX1_15 ( .A(_1770_), .Y(_1771_) );
OAI21X1 OAI21X1_448 ( .A(_1769_), .B(bundleStartMajId_i[31]), .C(_611__bF_buf0), .Y(_1772_) );
NAND2X1 NAND2X1_204 ( .A(_3653__31_), .B(_1039__bF_buf43), .Y(_1773_) );
OAI21X1 OAI21X1_449 ( .A(_1771_), .B(_1772_), .C(_1773_), .Y(_451_) );
XNOR2X1 XNOR2X1_13 ( .A(_1770_), .B(_1554_), .Y(_1774_) );
NAND2X1 NAND2X1_205 ( .A(_3653__30_), .B(_1039__bF_buf55), .Y(_1775_) );
OAI21X1 OAI21X1_450 ( .A(_1774_), .B(_1039__bF_buf43), .C(_1775_), .Y(_452_) );
NAND2X1 NAND2X1_206 ( .A(bundleStartMajId_i[30]), .B(bundleStartMajId_i[29]), .Y(_1776_) );
NOR2X1 NOR2X1_24 ( .A(_1776_), .B(_1770_), .Y(_1777_) );
INVX1 INVX1_16 ( .A(_1769_), .Y(_1778_) );
NOR2X1 NOR2X1_25 ( .A(_1552_), .B(_1554_), .Y(_1779_) );
INVX2 INVX2_43 ( .A(_1779_), .Y(_1780_) );
NOR2X1 NOR2X1_26 ( .A(_1780_), .B(_1778_), .Y(_1781_) );
OAI21X1 OAI21X1_451 ( .A(_1781_), .B(bundleStartMajId_i[29]), .C(_611__bF_buf0), .Y(_1782_) );
NAND2X1 NAND2X1_207 ( .A(_3653__29_), .B(_1039__bF_buf43), .Y(_1783_) );
OAI21X1 OAI21X1_452 ( .A(_1782_), .B(_1777_), .C(_1783_), .Y(_453_) );
XNOR2X1 XNOR2X1_14 ( .A(_1777_), .B(bundleStartMajId_i[28]), .Y(_1784_) );
NAND2X1 NAND2X1_208 ( .A(_3653__28_), .B(_1039__bF_buf1), .Y(_1785_) );
OAI21X1 OAI21X1_453 ( .A(_1784_), .B(_1039__bF_buf1), .C(_1785_), .Y(_454_) );
NOR2X1 NOR2X1_27 ( .A(_1694_), .B(_1713_), .Y(_1786_) );
NAND3X1 NAND3X1_4 ( .A(_1723_), .B(_1724_), .C(_1786_), .Y(_1787_) );
NOR2X1 NOR2X1_28 ( .A(_1740_), .B(_1753_), .Y(_1788_) );
NOR2X1 NOR2X1_29 ( .A(_1544_), .B(_1550_), .Y(_1789_) );
NAND3X1 NAND3X1_5 ( .A(_1789_), .B(_1765_), .C(_1788_), .Y(_1790_) );
NOR2X1 NOR2X1_30 ( .A(_1787_), .B(_1790_), .Y(_1791_) );
NAND2X1 NAND2X1_209 ( .A(bundleStartMajId_i[31]), .B(bundleStartMajId_i[28]), .Y(_1792_) );
NOR2X1 NOR2X1_31 ( .A(_1776_), .B(_1792_), .Y(_1793_) );
NAND3X1 NAND3X1_6 ( .A(_1793_), .B(_1687_), .C(_1791_), .Y(_1794_) );
XNOR2X1 XNOR2X1_15 ( .A(_1794_), .B(_1560_), .Y(_1795_) );
NAND2X1 NAND2X1_210 ( .A(_3653__27_), .B(_1039__bF_buf13), .Y(_1796_) );
OAI21X1 OAI21X1_454 ( .A(_1795_), .B(_1039__bF_buf13), .C(_1796_), .Y(_455_) );
NOR2X1 NOR2X1_32 ( .A(_1560_), .B(_1794_), .Y(_1797_) );
XNOR2X1 XNOR2X1_16 ( .A(_1797_), .B(bundleStartMajId_i[26]), .Y(_1798_) );
NAND2X1 NAND2X1_211 ( .A(_3653__26_), .B(_1039__bF_buf16), .Y(_1799_) );
OAI21X1 OAI21X1_455 ( .A(_1798_), .B(_1039__bF_buf16), .C(_1799_), .Y(_456_) );
NAND2X1 NAND2X1_212 ( .A(bundleStartMajId_i[27]), .B(bundleStartMajId_i[26]), .Y(_1800_) );
NOR2X1 NOR2X1_33 ( .A(_1800_), .B(_1794_), .Y(_1801_) );
XNOR2X1 XNOR2X1_17 ( .A(_1801_), .B(bundleStartMajId_i[25]), .Y(_1802_) );
NAND2X1 NAND2X1_213 ( .A(_3653__25_), .B(_1039__bF_buf24), .Y(_1803_) );
OAI21X1 OAI21X1_456 ( .A(_1802_), .B(_1039__bF_buf24), .C(_1803_), .Y(_457_) );
NAND2X1 NAND2X1_214 ( .A(_3653__24_), .B(_1039__bF_buf24), .Y(_1804_) );
NAND2X1 NAND2X1_215 ( .A(bundleStartMajId_i[25]), .B(_1801_), .Y(_1805_) );
XNOR2X1 XNOR2X1_18 ( .A(_1805_), .B(_1566_), .Y(_1806_) );
OAI21X1 OAI21X1_457 ( .A(_1806_), .B(_1039__bF_buf24), .C(_1804_), .Y(_458_) );
NAND2X1 NAND2X1_216 ( .A(bundleStartMajId_i[25]), .B(bundleStartMajId_i[24]), .Y(_1807_) );
NOR2X1 NOR2X1_34 ( .A(_1800_), .B(_1807_), .Y(_1808_) );
AND2X2 AND2X2_7 ( .A(_1793_), .B(_1808_), .Y(_1809_) );
NAND3X1 NAND3X1_7 ( .A(_1809_), .B(_1687_), .C(_1791_), .Y(_1810_) );
NOR2X1 NOR2X1_35 ( .A(_1568_), .B(_1810_), .Y(_1811_) );
INVX1 INVX1_17 ( .A(_1810_), .Y(_1812_) );
OAI21X1 OAI21X1_458 ( .A(_1812_), .B(bundleStartMajId_i[23]), .C(_611__bF_buf4), .Y(_1813_) );
NAND2X1 NAND2X1_217 ( .A(_3653__23_), .B(_1039__bF_buf33), .Y(_1814_) );
OAI21X1 OAI21X1_459 ( .A(_1813_), .B(_1811_), .C(_1814_), .Y(_459_) );
NAND2X1 NAND2X1_218 ( .A(bundleStartMajId_i[22]), .B(_1811_), .Y(_1815_) );
OAI21X1 OAI21X1_460 ( .A(_1810_), .B(_1568_), .C(_1570_), .Y(_1816_) );
NAND2X1 NAND2X1_219 ( .A(_1816_), .B(_1815_), .Y(_1817_) );
NAND2X1 NAND2X1_220 ( .A(_3653__22_), .B(_1039__bF_buf33), .Y(_1818_) );
OAI21X1 OAI21X1_461 ( .A(_1817_), .B(_1039__bF_buf33), .C(_1818_), .Y(_460_) );
NAND2X1 NAND2X1_221 ( .A(bundleStartMajId_i[23]), .B(bundleStartMajId_i[22]), .Y(_1819_) );
NOR2X1 NOR2X1_36 ( .A(_1819_), .B(_1810_), .Y(_1820_) );
NOR2X1 NOR2X1_37 ( .A(bundleStartMajId_i[21]), .B(_1820_), .Y(_1821_) );
OAI21X1 OAI21X1_462 ( .A(_1815_), .B(_1572_), .C(_611__bF_buf4), .Y(_1822_) );
NAND2X1 NAND2X1_222 ( .A(_3653__21_), .B(_1039__bF_buf33), .Y(_1823_) );
OAI21X1 OAI21X1_463 ( .A(_1822_), .B(_1821_), .C(_1823_), .Y(_461_) );
NAND2X1 NAND2X1_223 ( .A(_3653__20_), .B(_1039__bF_buf54), .Y(_1824_) );
NAND2X1 NAND2X1_224 ( .A(bundleStartMajId_i[21]), .B(_1820_), .Y(_1825_) );
XNOR2X1 XNOR2X1_19 ( .A(_1825_), .B(_1574_), .Y(_1826_) );
OAI21X1 OAI21X1_464 ( .A(_1826_), .B(_1039__bF_buf54), .C(_1824_), .Y(_462_) );
NAND3X1 NAND3X1_8 ( .A(bundleStartMajId_i[23]), .B(bundleStartMajId_i[22]), .C(bundleStartMajId_i[21]), .Y(_1827_) );
NOR2X1 NOR2X1_38 ( .A(_1574_), .B(_1827_), .Y(_1828_) );
INVX2 INVX2_44 ( .A(_1828_), .Y(_1829_) );
NOR3X1 NOR3X1_2 ( .A(_1576_), .B(_1829_), .C(_1810_), .Y(_1830_) );
OAI21X1 OAI21X1_465 ( .A(_1810_), .B(_1829_), .C(_1576_), .Y(_1831_) );
NAND2X1 NAND2X1_225 ( .A(_611__bF_buf1), .B(_1831_), .Y(_1832_) );
NAND2X1 NAND2X1_226 ( .A(_3653__19_), .B(_1039__bF_buf55), .Y(_1833_) );
OAI21X1 OAI21X1_466 ( .A(_1832_), .B(_1830_), .C(_1833_), .Y(_463_) );
XNOR2X1 XNOR2X1_20 ( .A(_1830_), .B(bundleStartMajId_i[18]), .Y(_1834_) );
NAND2X1 NAND2X1_227 ( .A(_3653__18_), .B(_1039__bF_buf12), .Y(_1835_) );
OAI21X1 OAI21X1_467 ( .A(_1834_), .B(_1039__bF_buf38), .C(_1835_), .Y(_464_) );
NAND2X1 NAND2X1_228 ( .A(_3653__17_), .B(_1039__bF_buf22), .Y(_1836_) );
NOR2X1 NOR2X1_39 ( .A(_1578_), .B(_1580_), .Y(_1837_) );
AND2X2 AND2X2_8 ( .A(_1830_), .B(_1837_), .Y(_1838_) );
AND2X2 AND2X2_9 ( .A(_1830_), .B(bundleStartMajId_i[18]), .Y(_1839_) );
OAI21X1 OAI21X1_468 ( .A(_1839_), .B(bundleStartMajId_i[17]), .C(_611__bF_buf1), .Y(_1840_) );
OAI21X1 OAI21X1_469 ( .A(_1840_), .B(_1838_), .C(_1836_), .Y(_465_) );
NAND2X1 NAND2X1_229 ( .A(_3653__16_), .B(_1039__bF_buf55), .Y(_1841_) );
NOR2X1 NOR2X1_40 ( .A(bundleStartMajId_i[16]), .B(_1838_), .Y(_1842_) );
NAND3X1 NAND3X1_9 ( .A(bundleStartMajId_i[18]), .B(bundleStartMajId_i[17]), .C(bundleStartMajId_i[16]), .Y(_1843_) );
NAND2X1 NAND2X1_230 ( .A(bundleStartMajId_i[20]), .B(bundleStartMajId_i[19]), .Y(_1844_) );
NOR3X1 NOR3X1_3 ( .A(_1827_), .B(_1844_), .C(_1843_), .Y(_1845_) );
NAND2X1 NAND2X1_231 ( .A(_1845_), .B(_1809_), .Y(_1846_) );
OAI21X1 OAI21X1_470 ( .A(_1778_), .B(_1846_), .C(_611__bF_buf1), .Y(_1847_) );
OAI21X1 OAI21X1_471 ( .A(_1842_), .B(_1847_), .C(_1841_), .Y(_466_) );
NAND2X1 NAND2X1_232 ( .A(_1793_), .B(_1808_), .Y(_1848_) );
INVX1 INVX1_18 ( .A(_1843_), .Y(_1849_) );
NOR2X1 NOR2X1_41 ( .A(_1844_), .B(_1827_), .Y(_1850_) );
NAND2X1 NAND2X1_233 ( .A(_1849_), .B(_1850_), .Y(_1851_) );
NOR2X1 NOR2X1_42 ( .A(_1848_), .B(_1851_), .Y(_1852_) );
NAND3X1 NAND3X1_10 ( .A(_1687_), .B(_1852_), .C(_1791_), .Y(_1853_) );
NOR2X1 NOR2X1_43 ( .A(_1584_), .B(_1853_), .Y(_1854_) );
INVX1 INVX1_19 ( .A(_1853_), .Y(_1855_) );
OAI21X1 OAI21X1_472 ( .A(_1855_), .B(bundleStartMajId_i[15]), .C(_611__bF_buf4), .Y(_1856_) );
NAND2X1 NAND2X1_234 ( .A(_3653__15_), .B(_1039__bF_buf33), .Y(_1857_) );
OAI21X1 OAI21X1_473 ( .A(_1856_), .B(_1854_), .C(_1857_), .Y(_467_) );
NAND2X1 NAND2X1_235 ( .A(bundleStartMajId_i[14]), .B(_1854_), .Y(_1858_) );
OAI21X1 OAI21X1_474 ( .A(_1853_), .B(_1584_), .C(_1586_), .Y(_1859_) );
NAND2X1 NAND2X1_236 ( .A(_1859_), .B(_1858_), .Y(_1860_) );
NAND2X1 NAND2X1_237 ( .A(_3653__14_), .B(_1039__bF_buf37), .Y(_1861_) );
OAI21X1 OAI21X1_475 ( .A(_1860_), .B(_1039__bF_buf54), .C(_1861_), .Y(_468_) );
NAND2X1 NAND2X1_238 ( .A(bundleStartMajId_i[15]), .B(bundleStartMajId_i[14]), .Y(_1862_) );
NOR2X1 NOR2X1_44 ( .A(_1862_), .B(_1853_), .Y(_1863_) );
NOR2X1 NOR2X1_45 ( .A(bundleStartMajId_i[13]), .B(_1863_), .Y(_1864_) );
OAI21X1 OAI21X1_476 ( .A(_1858_), .B(_1588_), .C(_611__bF_buf4), .Y(_1865_) );
NAND2X1 NAND2X1_239 ( .A(_3653__13_), .B(_1039__bF_buf33), .Y(_1866_) );
OAI21X1 OAI21X1_477 ( .A(_1865_), .B(_1864_), .C(_1866_), .Y(_469_) );
NAND2X1 NAND2X1_240 ( .A(_3653__12_), .B(_1039__bF_buf37), .Y(_1867_) );
NAND2X1 NAND2X1_241 ( .A(bundleStartMajId_i[13]), .B(_1863_), .Y(_1868_) );
XNOR2X1 XNOR2X1_21 ( .A(_1868_), .B(_1590_), .Y(_1869_) );
OAI21X1 OAI21X1_478 ( .A(_1869_), .B(_1039__bF_buf37), .C(_1867_), .Y(_470_) );
NOR2X1 NOR2X1_46 ( .A(_1586_), .B(_1588_), .Y(_1870_) );
NAND2X1 NAND2X1_242 ( .A(bundleStartMajId_i[15]), .B(_1870_), .Y(_1871_) );
INVX2 INVX2_45 ( .A(_1871_), .Y(_1872_) );
NAND2X1 NAND2X1_243 ( .A(bundleStartMajId_i[12]), .B(_1872_), .Y(_1873_) );
NOR2X1 NOR2X1_47 ( .A(_1873_), .B(_1853_), .Y(_1874_) );
NAND2X1 NAND2X1_244 ( .A(bundleStartMajId_i[11]), .B(_1874_), .Y(_1875_) );
INVX1 INVX1_20 ( .A(_1875_), .Y(_1876_) );
OAI21X1 OAI21X1_479 ( .A(_1874_), .B(bundleStartMajId_i[11]), .C(_611__bF_buf5), .Y(_1877_) );
NAND2X1 NAND2X1_245 ( .A(_3653__11_), .B(_1039__bF_buf55), .Y(_1878_) );
OAI21X1 OAI21X1_480 ( .A(_1876_), .B(_1877_), .C(_1878_), .Y(_471_) );
XNOR2X1 XNOR2X1_22 ( .A(_1875_), .B(_1594_), .Y(_1879_) );
NAND2X1 NAND2X1_246 ( .A(_3653__10_), .B(_1039__bF_buf55), .Y(_1880_) );
OAI21X1 OAI21X1_481 ( .A(_1879_), .B(_1039__bF_buf55), .C(_1880_), .Y(_472_) );
NAND2X1 NAND2X1_247 ( .A(_3653__9_), .B(_1039__bF_buf55), .Y(_1881_) );
NOR2X1 NOR2X1_48 ( .A(_1594_), .B(_1596_), .Y(_1882_) );
INVX2 INVX2_46 ( .A(_1882_), .Y(_1883_) );
NOR2X1 NOR2X1_49 ( .A(_1883_), .B(_1875_), .Y(_1884_) );
NOR2X1 NOR2X1_50 ( .A(_1592_), .B(_1594_), .Y(_1885_) );
AND2X2 AND2X2_10 ( .A(_1874_), .B(_1885_), .Y(_1886_) );
OAI21X1 OAI21X1_482 ( .A(_1886_), .B(bundleStartMajId_i[9]), .C(_611__bF_buf5), .Y(_1887_) );
OAI21X1 OAI21X1_483 ( .A(_1887_), .B(_1884_), .C(_1881_), .Y(_473_) );
NAND2X1 NAND2X1_248 ( .A(_3653__8_), .B(_1039__bF_buf55), .Y(_1888_) );
AOI21X1 AOI21X1_3 ( .A(_1882_), .B(_1876_), .C(bundleStartMajId_i[8]), .Y(_1889_) );
NAND2X1 NAND2X1_249 ( .A(bundleStartMajId_i[8]), .B(_1882_), .Y(_1890_) );
OAI21X1 OAI21X1_484 ( .A(_1875_), .B(_1890_), .C(_611__bF_buf1), .Y(_1891_) );
OAI21X1 OAI21X1_485 ( .A(_1889_), .B(_1891_), .C(_1888_), .Y(_474_) );
INVX1 INVX1_21 ( .A(_1890_), .Y(_1892_) );
NOR2X1 NOR2X1_51 ( .A(_1590_), .B(_1592_), .Y(_1893_) );
NAND3X1 NAND3X1_11 ( .A(_1893_), .B(_1872_), .C(_1892_), .Y(_1894_) );
NOR2X1 NOR2X1_52 ( .A(_1894_), .B(_1853_), .Y(_1895_) );
NAND2X1 NAND2X1_250 ( .A(bundleStartMajId_i[7]), .B(_1895_), .Y(_1896_) );
INVX1 INVX1_22 ( .A(_1896_), .Y(_1897_) );
OAI21X1 OAI21X1_486 ( .A(_1895_), .B(bundleStartMajId_i[7]), .C(_611__bF_buf5), .Y(_1898_) );
NAND2X1 NAND2X1_251 ( .A(_3653__7_), .B(_1039__bF_buf16), .Y(_1899_) );
OAI21X1 OAI21X1_487 ( .A(_1897_), .B(_1898_), .C(_1899_), .Y(_475_) );
NOR2X1 NOR2X1_53 ( .A(_1600_), .B(_1602_), .Y(_1900_) );
NAND2X1 NAND2X1_252 ( .A(_1900_), .B(_1895_), .Y(_1901_) );
INVX2 INVX2_47 ( .A(_1894_), .Y(_1902_) );
NAND2X1 NAND2X1_253 ( .A(_1902_), .B(_1855_), .Y(_1903_) );
OAI21X1 OAI21X1_488 ( .A(_1903_), .B(_1600_), .C(_1602_), .Y(_1904_) );
NAND2X1 NAND2X1_254 ( .A(_1901_), .B(_1904_), .Y(_1905_) );
NAND2X1 NAND2X1_255 ( .A(_3653__6_), .B(_1039__bF_buf16), .Y(_1906_) );
OAI21X1 OAI21X1_489 ( .A(_1905_), .B(_1039__bF_buf24), .C(_1906_), .Y(_476_) );
XNOR2X1 XNOR2X1_23 ( .A(_1901_), .B(_1604_), .Y(_1907_) );
NAND2X1 NAND2X1_256 ( .A(_3653__5_), .B(_1039__bF_buf6), .Y(_1908_) );
OAI21X1 OAI21X1_490 ( .A(_1907_), .B(_1039__bF_buf6), .C(_1908_), .Y(_477_) );
NAND2X1 NAND2X1_257 ( .A(_3653__4_), .B(_1039__bF_buf24), .Y(_1909_) );
NOR2X1 NOR2X1_54 ( .A(_1602_), .B(_1604_), .Y(_1910_) );
AOI21X1 AOI21X1_4 ( .A(_1910_), .B(_1897_), .C(bundleStartMajId_i[4]), .Y(_1911_) );
NAND2X1 NAND2X1_258 ( .A(bundleStartMajId_i[4]), .B(_1910_), .Y(_1912_) );
OAI21X1 OAI21X1_491 ( .A(_1896_), .B(_1912_), .C(_611__bF_buf5), .Y(_1913_) );
OAI21X1 OAI21X1_492 ( .A(_1911_), .B(_1913_), .C(_1909_), .Y(_478_) );
NAND2X1 NAND2X1_259 ( .A(_3653__3_), .B(_1039__bF_buf16), .Y(_1914_) );
NOR2X1 NOR2X1_55 ( .A(_1600_), .B(_1912_), .Y(_1915_) );
AOI21X1 AOI21X1_5 ( .A(_1915_), .B(_1895_), .C(bundleStartMajId_i[3]), .Y(_1916_) );
NAND2X1 NAND2X1_260 ( .A(bundleStartMajId_i[3]), .B(_1915_), .Y(_1917_) );
OAI21X1 OAI21X1_493 ( .A(_1903_), .B(_1917_), .C(_611__bF_buf5), .Y(_1918_) );
OAI21X1 OAI21X1_494 ( .A(_1918_), .B(_1916_), .C(_1914_), .Y(_479_) );
NAND2X1 NAND2X1_261 ( .A(_3653__2_), .B(_1039__bF_buf16), .Y(_1919_) );
NOR3X1 NOR3X1_4 ( .A(_1894_), .B(_1917_), .C(_1853_), .Y(_1920_) );
NOR2X1 NOR2X1_56 ( .A(bundleStartMajId_i[2]), .B(_1920_), .Y(_1921_) );
INVX1 INVX1_23 ( .A(_1917_), .Y(_1922_) );
NAND2X1 NAND2X1_262 ( .A(_1922_), .B(_1895_), .Y(_1923_) );
OAI21X1 OAI21X1_495 ( .A(_1923_), .B(_1610_), .C(_611__bF_buf5), .Y(_1924_) );
OAI21X1 OAI21X1_496 ( .A(_1924_), .B(_1921_), .C(_1919_), .Y(_480_) );
NAND2X1 NAND2X1_263 ( .A(_3653__1_), .B(_1039__bF_buf16), .Y(_1925_) );
AOI21X1 AOI21X1_6 ( .A(bundleStartMajId_i[2]), .B(_1920_), .C(bundleStartMajId_i[1]), .Y(_1926_) );
NOR2X1 NOR2X1_57 ( .A(_1610_), .B(_1612_), .Y(_1927_) );
INVX4 INVX4_28 ( .A(_1927_), .Y(_1928_) );
OAI21X1 OAI21X1_497 ( .A(_1923_), .B(_1928_), .C(_611__bF_buf5), .Y(_1929_) );
OAI21X1 OAI21X1_498 ( .A(_1929_), .B(_1926_), .C(_1925_), .Y(_481_) );
NAND2X1 NAND2X1_264 ( .A(_3653__0_), .B(_1039__bF_buf2), .Y(_1930_) );
NAND3X1 NAND3X1_12 ( .A(bundleStartMajId_i[0]), .B(_1927_), .C(_1920_), .Y(_1931_) );
OAI21X1 OAI21X1_499 ( .A(_1923_), .B(_1928_), .C(_1614_), .Y(_1932_) );
NAND3X1 NAND3X1_13 ( .A(_611__bF_buf5), .B(_1931_), .C(_1932_), .Y(_1933_) );
NAND2X1 NAND2X1_265 ( .A(_1930_), .B(_1933_), .Y(_482_) );
OAI21X1 OAI21X1_500 ( .A(_1100__bF_buf10_bF_buf3), .B(_1031__bF_buf26), .C(_3654__63_), .Y(_1934_) );
OAI21X1 OAI21X1_501 ( .A(_1101__bF_buf3), .B(_1488_), .C(_1934_), .Y(_483_) );
OAI21X1 OAI21X1_502 ( .A(_1100__bF_buf9_bF_buf3), .B(_1031__bF_buf23), .C(_3654__62_), .Y(_1935_) );
OAI21X1 OAI21X1_503 ( .A(_1101__bF_buf44), .B(bundleStartMajId_i[62]), .C(_1935_), .Y(_484_) );
NAND2X1 NAND2X1_266 ( .A(_1490_), .B(_1492_), .Y(_1936_) );
NAND2X1 NAND2X1_267 ( .A(_1623_), .B(_1936_), .Y(_1937_) );
OAI21X1 OAI21X1_504 ( .A(_1100__bF_buf8_bF_buf1), .B(_1031__bF_buf23), .C(_3654__61_), .Y(_1938_) );
OAI21X1 OAI21X1_505 ( .A(_1937_), .B(_1101__bF_buf44), .C(_1938_), .Y(_485_) );
INVX1 INVX1_24 ( .A(_1623_), .Y(_1939_) );
NAND2X1 NAND2X1_268 ( .A(bundleStartMajId_i[60]), .B(_1939_), .Y(_1940_) );
INVX1 INVX1_25 ( .A(_1940_), .Y(_1941_) );
OAI21X1 OAI21X1_506 ( .A(_1939_), .B(bundleStartMajId_i[60]), .C(_612__bF_buf6), .Y(_1942_) );
OAI21X1 OAI21X1_507 ( .A(_1100__bF_buf7_bF_buf2), .B(_1031__bF_buf68), .C(_3654__60_), .Y(_1943_) );
OAI21X1 OAI21X1_508 ( .A(_1941_), .B(_1942_), .C(_1943_), .Y(_486_) );
NAND2X1 NAND2X1_269 ( .A(bundleStartMajId_i[60]), .B(bundleStartMajId_i[59]), .Y(_1944_) );
OAI21X1 OAI21X1_509 ( .A(_1623_), .B(_1494_), .C(_1496_), .Y(_1945_) );
OAI21X1 OAI21X1_510 ( .A(_1623_), .B(_1944_), .C(_1945_), .Y(_1946_) );
OAI21X1 OAI21X1_511 ( .A(_1100__bF_buf6), .B(_1031__bF_buf33), .C(_3654__59_), .Y(_1947_) );
OAI21X1 OAI21X1_512 ( .A(_1946_), .B(_1101__bF_buf16), .C(_1947_), .Y(_487_) );
NOR2X1 NOR2X1_58 ( .A(_1637_), .B(_1940_), .Y(_1948_) );
NOR2X1 NOR2X1_59 ( .A(_1623_), .B(_1944_), .Y(_1949_) );
OAI21X1 OAI21X1_513 ( .A(_1949_), .B(bundleStartMajId_i[58]), .C(_612__bF_buf6), .Y(_1950_) );
OAI21X1 OAI21X1_514 ( .A(_1100__bF_buf6), .B(_1031__bF_buf23), .C(_3654__58_), .Y(_1951_) );
OAI21X1 OAI21X1_515 ( .A(_1948_), .B(_1950_), .C(_1951_), .Y(_488_) );
INVX4 INVX4_29 ( .A(_1948_), .Y(_1952_) );
XNOR2X1 XNOR2X1_24 ( .A(_1952_), .B(_1500_), .Y(_1953_) );
OAI21X1 OAI21X1_516 ( .A(_1100__bF_buf6), .B(_1031__bF_buf0), .C(_3654__57_), .Y(_1954_) );
OAI21X1 OAI21X1_517 ( .A(_1953_), .B(_1101__bF_buf16), .C(_1954_), .Y(_489_) );
OAI21X1 OAI21X1_518 ( .A(_1952_), .B(_1500_), .C(_1502_), .Y(_1955_) );
OAI21X1 OAI21X1_519 ( .A(_1646_), .B(_1952_), .C(_1955_), .Y(_1956_) );
OAI21X1 OAI21X1_520 ( .A(_1100__bF_buf6), .B(_1031__bF_buf30), .C(_3654__56_), .Y(_1957_) );
OAI21X1 OAI21X1_521 ( .A(_1956_), .B(_1101__bF_buf16), .C(_1957_), .Y(_490_) );
NAND2X1 NAND2X1_270 ( .A(bundleStartMajId_i[56]), .B(bundleStartMajId_i[55]), .Y(_1958_) );
NOR2X1 NOR2X1_60 ( .A(_1641_), .B(_1958_), .Y(_1959_) );
AND2X2 AND2X2_11 ( .A(_1949_), .B(_1959_), .Y(_1960_) );
INVX4 INVX4_30 ( .A(_1960_), .Y(_1961_) );
OAI21X1 OAI21X1_522 ( .A(_1952_), .B(_1646_), .C(_1504_), .Y(_1962_) );
NAND2X1 NAND2X1_271 ( .A(_1961_), .B(_1962_), .Y(_1963_) );
OAI21X1 OAI21X1_523 ( .A(_1100__bF_buf6), .B(_1031__bF_buf0), .C(_3654__55_), .Y(_1964_) );
OAI21X1 OAI21X1_524 ( .A(_1963_), .B(_1101__bF_buf12), .C(_1964_), .Y(_491_) );
XNOR2X1 XNOR2X1_25 ( .A(_1960_), .B(bundleStartMajId_i[54]), .Y(_1965_) );
OAI21X1 OAI21X1_525 ( .A(_1100__bF_buf4), .B(_1031__bF_buf65), .C(_3654__54_), .Y(_1966_) );
OAI21X1 OAI21X1_526 ( .A(_1965_), .B(_1101__bF_buf18), .C(_1966_), .Y(_492_) );
OAI21X1 OAI21X1_527 ( .A(_1961_), .B(_1506_), .C(_1508_), .Y(_1967_) );
OAI21X1 OAI21X1_528 ( .A(_1659_), .B(_1961_), .C(_1967_), .Y(_1968_) );
OAI21X1 OAI21X1_529 ( .A(_1100__bF_buf6), .B(_1031__bF_buf0), .C(_3654__53_), .Y(_1969_) );
OAI21X1 OAI21X1_530 ( .A(_1968_), .B(_1101__bF_buf16), .C(_1969_), .Y(_493_) );
NAND2X1 NAND2X1_272 ( .A(bundleStartMajId_i[52]), .B(_1662_), .Y(_1970_) );
OAI21X1 OAI21X1_531 ( .A(_1961_), .B(_1659_), .C(_1510_), .Y(_1971_) );
OAI21X1 OAI21X1_532 ( .A(_1970_), .B(_1961_), .C(_1971_), .Y(_1972_) );
OAI21X1 OAI21X1_533 ( .A(_1100__bF_buf14_bF_buf0), .B(_1031__bF_buf16), .C(_3654__52_), .Y(_1973_) );
OAI21X1 OAI21X1_534 ( .A(_1972_), .B(_1101__bF_buf57), .C(_1973_), .Y(_494_) );
NAND3X1 NAND3X1_14 ( .A(bundleStartMajId_i[52]), .B(_1662_), .C(_1960_), .Y(_1974_) );
XNOR2X1 XNOR2X1_26 ( .A(_1974_), .B(_1512_), .Y(_1975_) );
OAI21X1 OAI21X1_535 ( .A(_1100__bF_buf13_bF_buf1), .B(_1031__bF_buf43), .C(_3654__51_), .Y(_1976_) );
OAI21X1 OAI21X1_536 ( .A(_1975_), .B(_1101__bF_buf57), .C(_1976_), .Y(_495_) );
INVX1 INVX1_26 ( .A(_1676_), .Y(_1977_) );
NOR2X1 NOR2X1_61 ( .A(_1512_), .B(_1974_), .Y(_1978_) );
OAI22X1 OAI22X1_1 ( .A(_1977_), .B(_1974_), .C(_1978_), .D(bundleStartMajId_i[50]), .Y(_1979_) );
OAI21X1 OAI21X1_537 ( .A(_1100__bF_buf12_bF_buf3), .B(_1031__bF_buf30), .C(_3654__50_), .Y(_1980_) );
OAI21X1 OAI21X1_538 ( .A(_1979_), .B(_1101__bF_buf12), .C(_1980_), .Y(_496_) );
AND2X2 AND2X2_12 ( .A(bundleStartMajId_i[50]), .B(bundleStartMajId_i[49]), .Y(_1981_) );
NAND2X1 NAND2X1_273 ( .A(_1981_), .B(_1978_), .Y(_1982_) );
OAI21X1 OAI21X1_539 ( .A(_1974_), .B(_1977_), .C(_1516_), .Y(_1983_) );
NAND2X1 NAND2X1_274 ( .A(_1983_), .B(_1982_), .Y(_1984_) );
OAI21X1 OAI21X1_540 ( .A(_1100__bF_buf11_bF_buf2), .B(_1031__bF_buf23), .C(_3654__49_), .Y(_1985_) );
OAI21X1 OAI21X1_541 ( .A(_1984_), .B(_1101__bF_buf44), .C(_1985_), .Y(_497_) );
XNOR2X1 XNOR2X1_27 ( .A(_1982_), .B(_1518_), .Y(_1986_) );
OAI21X1 OAI21X1_542 ( .A(_1100__bF_buf10_bF_buf3), .B(_1031__bF_buf16), .C(_3654__48_), .Y(_1987_) );
OAI21X1 OAI21X1_543 ( .A(_1986_), .B(_1101__bF_buf12), .C(_1987_), .Y(_498_) );
OAI21X1 OAI21X1_544 ( .A(_1100__bF_buf9_bF_buf3), .B(_1031__bF_buf43), .C(_3654__47_), .Y(_1988_) );
OAI21X1 OAI21X1_545 ( .A(_1982_), .B(_1518_), .C(_1520_), .Y(_1989_) );
NAND3X1 NAND3X1_15 ( .A(bundleStartMajId_i[48]), .B(bundleStartMajId_i[47]), .C(_1981_), .Y(_1990_) );
NOR2X1 NOR2X1_62 ( .A(_1668_), .B(_1990_), .Y(_1991_) );
NAND2X1 NAND2X1_275 ( .A(_1960_), .B(_1991_), .Y(_1992_) );
NAND2X1 NAND2X1_276 ( .A(_1992_), .B(_1989_), .Y(_1993_) );
OAI21X1 OAI21X1_546 ( .A(_1993_), .B(_1101__bF_buf57), .C(_1988_), .Y(_499_) );
XNOR2X1 XNOR2X1_28 ( .A(_1992_), .B(_1522_), .Y(_1994_) );
OAI21X1 OAI21X1_547 ( .A(_1100__bF_buf8_bF_buf1), .B(_1031__bF_buf30), .C(_3654__46_), .Y(_1995_) );
OAI21X1 OAI21X1_548 ( .A(_1994_), .B(_1101__bF_buf44), .C(_1995_), .Y(_500_) );
OAI21X1 OAI21X1_549 ( .A(_1992_), .B(_1522_), .C(_1524_), .Y(_1996_) );
OAI21X1 OAI21X1_550 ( .A(_1694_), .B(_1992_), .C(_1996_), .Y(_1997_) );
OAI21X1 OAI21X1_551 ( .A(_1100__bF_buf7_bF_buf0), .B(_1031__bF_buf74), .C(_3654__45_), .Y(_1998_) );
OAI21X1 OAI21X1_552 ( .A(_1997_), .B(_1101__bF_buf49), .C(_1998_), .Y(_501_) );
OR2X2 OR2X2_5 ( .A(_1694_), .B(_1526_), .Y(_1999_) );
OAI21X1 OAI21X1_553 ( .A(_1992_), .B(_1694_), .C(_1526_), .Y(_2000_) );
OAI21X1 OAI21X1_554 ( .A(_1999_), .B(_1992_), .C(_2000_), .Y(_2001_) );
OAI21X1 OAI21X1_555 ( .A(_1100__bF_buf0), .B(_1031__bF_buf69), .C(_3654__44_), .Y(_2002_) );
OAI21X1 OAI21X1_556 ( .A(_2001_), .B(_1101__bF_buf4), .C(_2002_), .Y(_502_) );
NOR2X1 NOR2X1_63 ( .A(_1999_), .B(_1992_), .Y(_2003_) );
NOR2X1 NOR2X1_64 ( .A(bundleStartMajId_i[43]), .B(_2003_), .Y(_2004_) );
OAI21X1 OAI21X1_557 ( .A(_1992_), .B(_1705_), .C(_612__bF_buf1), .Y(_2005_) );
OAI21X1 OAI21X1_558 ( .A(_1100__bF_buf0), .B(_1031__bF_buf69), .C(_3654__43_), .Y(_2006_) );
OAI21X1 OAI21X1_559 ( .A(_2004_), .B(_2005_), .C(_2006_), .Y(_503_) );
NOR2X1 NOR2X1_65 ( .A(bundleStartMajId_i[42]), .B(_2005_), .Y(_2007_) );
NAND2X1 NAND2X1_277 ( .A(_1716_), .B(_2003_), .Y(_2008_) );
MUX2X1 MUX2X1_1 ( .A(_2008_), .B(_3654__42_), .S(_612__bF_buf1), .Y(_2009_) );
NOR2X1 NOR2X1_66 ( .A(_2007_), .B(_2009_), .Y(_504_) );
XNOR2X1 XNOR2X1_29 ( .A(_2008_), .B(_1532_), .Y(_2010_) );
OAI21X1 OAI21X1_560 ( .A(_1100__bF_buf0), .B(_1031__bF_buf51), .C(_3654__41_), .Y(_2011_) );
OAI21X1 OAI21X1_561 ( .A(_2010_), .B(_1101__bF_buf2), .C(_2011_), .Y(_505_) );
OAI21X1 OAI21X1_562 ( .A(_1100__bF_buf0), .B(_1031__bF_buf5), .C(_3654__40_), .Y(_2012_) );
NAND2X1 NAND2X1_278 ( .A(bundleStartMajId_i[42]), .B(bundleStartMajId_i[41]), .Y(_2013_) );
NOR2X1 NOR2X1_67 ( .A(_1694_), .B(_1704_), .Y(_2014_) );
AND2X2 AND2X2_13 ( .A(_1991_), .B(_1960_), .Y(_2015_) );
NAND2X1 NAND2X1_279 ( .A(_2014_), .B(_2015_), .Y(_2016_) );
NOR2X1 NOR2X1_68 ( .A(_2013_), .B(_2016_), .Y(_2017_) );
XNOR2X1 XNOR2X1_30 ( .A(_2017_), .B(bundleStartMajId_i[40]), .Y(_2018_) );
OAI21X1 OAI21X1_563 ( .A(_2018_), .B(_1101__bF_buf49), .C(_2012_), .Y(_506_) );
NAND2X1 NAND2X1_280 ( .A(bundleStartMajId_i[40]), .B(_2017_), .Y(_2019_) );
XNOR2X1 XNOR2X1_31 ( .A(_2019_), .B(_1536_), .Y(_2020_) );
OAI21X1 OAI21X1_564 ( .A(_1100__bF_buf0), .B(_1031__bF_buf5), .C(_3654__39_), .Y(_2021_) );
OAI21X1 OAI21X1_565 ( .A(_2020_), .B(_1101__bF_buf49), .C(_2021_), .Y(_507_) );
INVX1 INVX1_27 ( .A(_2016_), .Y(_2022_) );
NAND2X1 NAND2X1_281 ( .A(bundleStartMajId_i[40]), .B(bundleStartMajId_i[39]), .Y(_2023_) );
NOR2X1 NOR2X1_69 ( .A(_2013_), .B(_2023_), .Y(_2024_) );
NAND2X1 NAND2X1_282 ( .A(_2024_), .B(_2022_), .Y(_2025_) );
XNOR2X1 XNOR2X1_32 ( .A(_2025_), .B(_1538_), .Y(_2026_) );
OAI21X1 OAI21X1_566 ( .A(_1100__bF_buf0), .B(_1031__bF_buf10), .C(_3654__38_), .Y(_2027_) );
OAI21X1 OAI21X1_567 ( .A(_2026_), .B(_1101__bF_buf32), .C(_2027_), .Y(_508_) );
OAI21X1 OAI21X1_568 ( .A(_1100__bF_buf0), .B(_1031__bF_buf54), .C(_3654__37_), .Y(_2028_) );
OAI21X1 OAI21X1_569 ( .A(_2025_), .B(_1538_), .C(_1540_), .Y(_2029_) );
OAI21X1 OAI21X1_570 ( .A(_1740_), .B(_2025_), .C(_2029_), .Y(_2030_) );
OAI21X1 OAI21X1_571 ( .A(_2030_), .B(_1101__bF_buf32), .C(_2028_), .Y(_509_) );
OAI21X1 OAI21X1_572 ( .A(_1100__bF_buf14_bF_buf3), .B(_1031__bF_buf74), .C(_3654__36_), .Y(_2031_) );
NOR2X1 NOR2X1_70 ( .A(_1740_), .B(_2025_), .Y(_2032_) );
NOR2X1 NOR2X1_71 ( .A(bundleStartMajId_i[36]), .B(_2032_), .Y(_2033_) );
NAND2X1 NAND2X1_283 ( .A(bundleStartMajId_i[36]), .B(_1741_), .Y(_2034_) );
OAI21X1 OAI21X1_573 ( .A(_2025_), .B(_2034_), .C(_612__bF_buf1), .Y(_2035_) );
OAI21X1 OAI21X1_574 ( .A(_2033_), .B(_2035_), .C(_2031_), .Y(_510_) );
INVX1 INVX1_28 ( .A(_3654__35_), .Y(_2036_) );
OAI21X1 OAI21X1_575 ( .A(_2025_), .B(_2034_), .C(_1544_), .Y(_2037_) );
NAND2X1 NAND2X1_284 ( .A(_1746_), .B(_2024_), .Y(_2038_) );
OR2X2 OR2X2_6 ( .A(_2016_), .B(_2038_), .Y(_2039_) );
NAND3X1 NAND3X1_16 ( .A(_612__bF_buf1), .B(_2039_), .C(_2037_), .Y(_2040_) );
OAI21X1 OAI21X1_576 ( .A(_2036_), .B(_612__bF_buf1), .C(_2040_), .Y(_511_) );
NOR2X1 NOR2X1_72 ( .A(_2038_), .B(_2016_), .Y(_2041_) );
XNOR2X1 XNOR2X1_33 ( .A(_2041_), .B(bundleStartMajId_i[34]), .Y(_2042_) );
OAI21X1 OAI21X1_577 ( .A(_1100__bF_buf13_bF_buf0), .B(_1031__bF_buf10), .C(_3654__34_), .Y(_2043_) );
OAI21X1 OAI21X1_578 ( .A(_2042_), .B(_1101__bF_buf5), .C(_2043_), .Y(_512_) );
OAI21X1 OAI21X1_579 ( .A(_1100__bF_buf12_bF_buf0), .B(_1031__bF_buf10), .C(_3654__33_), .Y(_2044_) );
AOI21X1 AOI21X1_7 ( .A(bundleStartMajId_i[34]), .B(_2041_), .C(bundleStartMajId_i[33]), .Y(_2045_) );
NAND2X1 NAND2X1_285 ( .A(bundleStartMajId_i[34]), .B(bundleStartMajId_i[33]), .Y(_2046_) );
OAI21X1 OAI21X1_580 ( .A(_2039_), .B(_2046_), .C(_612__bF_buf1), .Y(_2047_) );
OAI21X1 OAI21X1_581 ( .A(_2047_), .B(_2045_), .C(_2044_), .Y(_513_) );
OAI21X1 OAI21X1_582 ( .A(_2039_), .B(_2046_), .C(_1550_), .Y(_2048_) );
NAND3X1 NAND3X1_17 ( .A(bundleStartMajId_i[32]), .B(_1765_), .C(_2041_), .Y(_2049_) );
NAND2X1 NAND2X1_286 ( .A(_2049_), .B(_2048_), .Y(_2050_) );
OAI21X1 OAI21X1_583 ( .A(_1100__bF_buf11_bF_buf3), .B(_1031__bF_buf54), .C(_3654__32_), .Y(_2051_) );
OAI21X1 OAI21X1_584 ( .A(_2050_), .B(_1101__bF_buf30), .C(_2051_), .Y(_514_) );
NOR2X1 NOR2X1_73 ( .A(_3654__31_), .B(_612__bF_buf1), .Y(_2052_) );
OR2X2 OR2X2_7 ( .A(_2049_), .B(bundleStartMajId_i[31]), .Y(_2053_) );
AOI21X1 AOI21X1_8 ( .A(bundleStartMajId_i[31]), .B(_2049_), .C(_1101__bF_buf4), .Y(_2054_) );
AOI21X1 AOI21X1_9 ( .A(_2054_), .B(_2053_), .C(_2052_), .Y(_515_) );
NAND2X1 NAND2X1_287 ( .A(bundleStartMajId_i[32]), .B(bundleStartMajId_i[31]), .Y(_2055_) );
NOR2X1 NOR2X1_74 ( .A(_2046_), .B(_2055_), .Y(_2056_) );
AND2X2 AND2X2_14 ( .A(_1746_), .B(_2056_), .Y(_2057_) );
NAND3X1 NAND3X1_18 ( .A(_2014_), .B(_2024_), .C(_2057_), .Y(_2058_) );
NOR2X1 NOR2X1_75 ( .A(_1992_), .B(_2058_), .Y(_2059_) );
XNOR2X1 XNOR2X1_34 ( .A(_2059_), .B(bundleStartMajId_i[30]), .Y(_2060_) );
OAI21X1 OAI21X1_585 ( .A(_1100__bF_buf10_bF_buf3), .B(_1031__bF_buf53), .C(_3654__30_), .Y(_2061_) );
OAI21X1 OAI21X1_586 ( .A(_2060_), .B(_1101__bF_buf48), .C(_2061_), .Y(_516_) );
NAND2X1 NAND2X1_288 ( .A(_2014_), .B(_2056_), .Y(_2062_) );
NOR2X1 NOR2X1_76 ( .A(_2038_), .B(_2062_), .Y(_2063_) );
NAND2X1 NAND2X1_289 ( .A(_2063_), .B(_2015_), .Y(_2064_) );
OAI21X1 OAI21X1_587 ( .A(_2064_), .B(_1554_), .C(_1556_), .Y(_2065_) );
OAI21X1 OAI21X1_588 ( .A(_1776_), .B(_2064_), .C(_2065_), .Y(_2066_) );
OAI21X1 OAI21X1_589 ( .A(_1100__bF_buf9_bF_buf3), .B(_1031__bF_buf53), .C(_3654__29_), .Y(_2067_) );
OAI21X1 OAI21X1_590 ( .A(_2066_), .B(_1101__bF_buf48), .C(_2067_), .Y(_517_) );
OR2X2 OR2X2_8 ( .A(_1776_), .B(_1558_), .Y(_2068_) );
OAI21X1 OAI21X1_591 ( .A(_2064_), .B(_1776_), .C(_1558_), .Y(_2069_) );
OAI21X1 OAI21X1_592 ( .A(_2068_), .B(_2064_), .C(_2069_), .Y(_2070_) );
OAI21X1 OAI21X1_593 ( .A(_1100__bF_buf8_bF_buf1), .B(_1031__bF_buf16), .C(_3654__28_), .Y(_2071_) );
OAI21X1 OAI21X1_594 ( .A(_2070_), .B(_1101__bF_buf57), .C(_2071_), .Y(_518_) );
NAND2X1 NAND2X1_290 ( .A(bundleStartMajId_i[28]), .B(bundleStartMajId_i[27]), .Y(_2072_) );
NOR2X1 NOR2X1_77 ( .A(_1776_), .B(_2072_), .Y(_2073_) );
INVX2 INVX2_48 ( .A(_2073_), .Y(_2074_) );
NOR2X1 NOR2X1_78 ( .A(_2068_), .B(_2064_), .Y(_2075_) );
OAI22X1 OAI22X1_2 ( .A(_2074_), .B(_2064_), .C(_2075_), .D(bundleStartMajId_i[27]), .Y(_2076_) );
OAI21X1 OAI21X1_595 ( .A(_1100__bF_buf7_bF_buf1), .B(_1031__bF_buf42), .C(_3654__27_), .Y(_2077_) );
OAI21X1 OAI21X1_596 ( .A(_2076_), .B(_1101__bF_buf24), .C(_2077_), .Y(_519_) );
OR2X2 OR2X2_9 ( .A(_2064_), .B(_2068_), .Y(_2078_) );
OAI21X1 OAI21X1_597 ( .A(_2064_), .B(_2074_), .C(_1562_), .Y(_2079_) );
OAI21X1 OAI21X1_598 ( .A(_2078_), .B(_1800_), .C(_2079_), .Y(_2080_) );
OAI21X1 OAI21X1_599 ( .A(_1100__bF_buf0), .B(_1031__bF_buf42), .C(_3654__26_), .Y(_2081_) );
OAI21X1 OAI21X1_600 ( .A(_2080_), .B(_1101__bF_buf24), .C(_2081_), .Y(_520_) );
OAI21X1 OAI21X1_601 ( .A(_1100__bF_buf0), .B(_1031__bF_buf5), .C(_3654__25_), .Y(_2082_) );
NAND2X1 NAND2X1_291 ( .A(_2073_), .B(_2059_), .Y(_2083_) );
NOR2X1 NOR2X1_79 ( .A(_1562_), .B(_2083_), .Y(_2084_) );
XNOR2X1 XNOR2X1_35 ( .A(_2084_), .B(bundleStartMajId_i[25]), .Y(_2085_) );
OAI21X1 OAI21X1_602 ( .A(_2085_), .B(_1101__bF_buf49), .C(_2082_), .Y(_521_) );
INVX1 INVX1_29 ( .A(_3654__24_), .Y(_2086_) );
NAND2X1 NAND2X1_292 ( .A(bundleStartMajId_i[26]), .B(bundleStartMajId_i[25]), .Y(_2087_) );
INVX1 INVX1_30 ( .A(_2087_), .Y(_2088_) );
OR2X2 OR2X2_10 ( .A(_2058_), .B(_1992_), .Y(_2089_) );
NOR2X1 NOR2X1_80 ( .A(_2074_), .B(_2089_), .Y(_2090_) );
AOI21X1 AOI21X1_10 ( .A(_2088_), .B(_2090_), .C(_1566_), .Y(_2091_) );
NOR3X1 NOR3X1_5 ( .A(bundleStartMajId_i[24]), .B(_2087_), .C(_2083_), .Y(_2092_) );
OAI21X1 OAI21X1_603 ( .A(_2091_), .B(_2092_), .C(_612__bF_buf6), .Y(_2093_) );
OAI21X1 OAI21X1_604 ( .A(_2086_), .B(_612__bF_buf6), .C(_2093_), .Y(_522_) );
NOR2X1 NOR2X1_81 ( .A(_3654__23_), .B(_612__bF_buf6), .Y(_2094_) );
NOR3X1 NOR3X1_6 ( .A(_1564_), .B(_1800_), .C(_2078_), .Y(_2095_) );
NAND3X1 NAND3X1_19 ( .A(bundleStartMajId_i[24]), .B(_1568_), .C(_2095_), .Y(_2096_) );
NAND3X1 NAND3X1_20 ( .A(bundleStartMajId_i[24]), .B(_2088_), .C(_2090_), .Y(_2097_) );
AOI21X1 AOI21X1_11 ( .A(bundleStartMajId_i[23]), .B(_2097_), .C(_1101__bF_buf24), .Y(_2098_) );
AOI21X1 AOI21X1_12 ( .A(_2098_), .B(_2096_), .C(_2094_), .Y(_523_) );
NAND3X1 NAND3X1_21 ( .A(_1746_), .B(_2024_), .C(_2056_), .Y(_2099_) );
NOR2X1 NOR2X1_82 ( .A(_1705_), .B(_2099_), .Y(_2100_) );
NAND2X1 NAND2X1_293 ( .A(bundleStartMajId_i[24]), .B(bundleStartMajId_i[23]), .Y(_2101_) );
NOR2X1 NOR2X1_83 ( .A(_2087_), .B(_2101_), .Y(_2102_) );
NAND2X1 NAND2X1_294 ( .A(_2073_), .B(_2102_), .Y(_2103_) );
INVX1 INVX1_31 ( .A(_2103_), .Y(_2104_) );
NAND3X1 NAND3X1_22 ( .A(_2100_), .B(_2104_), .C(_2015_), .Y(_2105_) );
XNOR2X1 XNOR2X1_36 ( .A(_2105_), .B(_1570_), .Y(_2106_) );
OAI21X1 OAI21X1_605 ( .A(_1100__bF_buf4), .B(_1031__bF_buf65), .C(_3654__22_), .Y(_2107_) );
OAI21X1 OAI21X1_606 ( .A(_2106_), .B(_1101__bF_buf18), .C(_2107_), .Y(_524_) );
OAI21X1 OAI21X1_607 ( .A(_1100__bF_buf8), .B(_1031__bF_buf63), .C(_3654__21_), .Y(_2108_) );
NOR2X1 NOR2X1_84 ( .A(_2103_), .B(_2064_), .Y(_2109_) );
AOI21X1 AOI21X1_13 ( .A(bundleStartMajId_i[22]), .B(_2109_), .C(bundleStartMajId_i[21]), .Y(_2110_) );
NAND2X1 NAND2X1_295 ( .A(bundleStartMajId_i[22]), .B(bundleStartMajId_i[21]), .Y(_2111_) );
INVX1 INVX1_32 ( .A(_2111_), .Y(_2112_) );
NAND2X1 NAND2X1_296 ( .A(_2112_), .B(_2109_), .Y(_2113_) );
NAND2X1 NAND2X1_297 ( .A(_612__bF_buf4), .B(_2113_), .Y(_2114_) );
OAI21X1 OAI21X1_608 ( .A(_2114_), .B(_2110_), .C(_2108_), .Y(_525_) );
OAI21X1 OAI21X1_609 ( .A(_1100__bF_buf4), .B(_1031__bF_buf26), .C(_3654__20_), .Y(_2115_) );
AND2X2 AND2X2_15 ( .A(_2109_), .B(_2112_), .Y(_2116_) );
NOR2X1 NOR2X1_85 ( .A(bundleStartMajId_i[20]), .B(_2116_), .Y(_2117_) );
OAI21X1 OAI21X1_610 ( .A(_2113_), .B(_1574_), .C(_612__bF_buf4), .Y(_2118_) );
OAI21X1 OAI21X1_611 ( .A(_2117_), .B(_2118_), .C(_2115_), .Y(_526_) );
OAI21X1 OAI21X1_612 ( .A(_1100__bF_buf4), .B(_1031__bF_buf26), .C(_3654__19_), .Y(_2119_) );
AOI21X1 AOI21X1_14 ( .A(bundleStartMajId_i[20]), .B(_2116_), .C(bundleStartMajId_i[19]), .Y(_2120_) );
NOR2X1 NOR2X1_86 ( .A(_2111_), .B(_1844_), .Y(_2121_) );
INVX2 INVX2_49 ( .A(_2121_), .Y(_2122_) );
OAI21X1 OAI21X1_613 ( .A(_2105_), .B(_2122_), .C(_612__bF_buf4), .Y(_2123_) );
OAI21X1 OAI21X1_614 ( .A(_2120_), .B(_2123_), .C(_2119_), .Y(_527_) );
OAI21X1 OAI21X1_615 ( .A(_1100__bF_buf0), .B(_1031__bF_buf43), .C(_3654__18_), .Y(_2124_) );
NOR2X1 NOR2X1_87 ( .A(_2122_), .B(_2105_), .Y(_2125_) );
NOR2X1 NOR2X1_88 ( .A(bundleStartMajId_i[18]), .B(_2125_), .Y(_2126_) );
INVX2 INVX2_50 ( .A(_2125_), .Y(_2127_) );
OAI21X1 OAI21X1_616 ( .A(_2127_), .B(_1578_), .C(_612__bF_buf6), .Y(_2128_) );
OAI21X1 OAI21X1_617 ( .A(_2128_), .B(_2126_), .C(_2124_), .Y(_528_) );
OAI21X1 OAI21X1_618 ( .A(_1100__bF_buf14_bF_buf0), .B(_1031__bF_buf16), .C(_3654__17_), .Y(_2129_) );
AOI21X1 AOI21X1_15 ( .A(bundleStartMajId_i[18]), .B(_2125_), .C(bundleStartMajId_i[17]), .Y(_2130_) );
INVX1 INVX1_33 ( .A(_1837_), .Y(_2131_) );
OAI21X1 OAI21X1_619 ( .A(_2127_), .B(_2131_), .C(_612__bF_buf6), .Y(_2132_) );
OAI21X1 OAI21X1_620 ( .A(_2132_), .B(_2130_), .C(_2129_), .Y(_529_) );
OAI21X1 OAI21X1_621 ( .A(_1100__bF_buf13_bF_buf1), .B(_1031__bF_buf16), .C(_3654__16_), .Y(_2133_) );
AOI21X1 AOI21X1_16 ( .A(_1837_), .B(_2125_), .C(bundleStartMajId_i[16]), .Y(_2134_) );
OAI21X1 OAI21X1_622 ( .A(_2127_), .B(_1843_), .C(_612__bF_buf6), .Y(_2135_) );
OAI21X1 OAI21X1_623 ( .A(_2135_), .B(_2134_), .C(_2133_), .Y(_530_) );
NOR2X1 NOR2X1_89 ( .A(_3654__15_), .B(_612__bF_buf6), .Y(_2136_) );
NAND2X1 NAND2X1_298 ( .A(_1849_), .B(_2125_), .Y(_2137_) );
OR2X2 OR2X2_11 ( .A(_2137_), .B(bundleStartMajId_i[15]), .Y(_2138_) );
AOI21X1 AOI21X1_17 ( .A(bundleStartMajId_i[15]), .B(_2137_), .C(_1101__bF_buf57), .Y(_2139_) );
AOI21X1 AOI21X1_18 ( .A(_2139_), .B(_2138_), .C(_2136_), .Y(_531_) );
NOR2X1 NOR2X1_90 ( .A(_1582_), .B(_1584_), .Y(_2140_) );
NAND3X1 NAND3X1_23 ( .A(_1837_), .B(_2140_), .C(_2121_), .Y(_2141_) );
NOR2X1 NOR2X1_91 ( .A(_2103_), .B(_2141_), .Y(_2142_) );
NAND3X1 NAND3X1_24 ( .A(_2063_), .B(_2142_), .C(_2015_), .Y(_2143_) );
XNOR2X1 XNOR2X1_37 ( .A(_2143_), .B(_1586_), .Y(_2144_) );
OAI21X1 OAI21X1_624 ( .A(_1100__bF_buf12_bF_buf2), .B(_1031__bF_buf21), .C(_3654__14_), .Y(_2145_) );
OAI21X1 OAI21X1_625 ( .A(_2144_), .B(_1101__bF_buf45), .C(_2145_), .Y(_532_) );
OAI21X1 OAI21X1_626 ( .A(_1100__bF_buf11_bF_buf0), .B(_1031__bF_buf41), .C(_3654__13_), .Y(_2146_) );
NOR2X1 NOR2X1_92 ( .A(_1586_), .B(_2143_), .Y(_2147_) );
NOR2X1 NOR2X1_93 ( .A(bundleStartMajId_i[13]), .B(_2147_), .Y(_2148_) );
INVX2 INVX2_51 ( .A(_1870_), .Y(_2149_) );
OAI21X1 OAI21X1_627 ( .A(_2143_), .B(_2149_), .C(_612__bF_buf4), .Y(_2150_) );
OAI21X1 OAI21X1_628 ( .A(_2148_), .B(_2150_), .C(_2146_), .Y(_533_) );
OAI21X1 OAI21X1_629 ( .A(_1100__bF_buf10_bF_buf3), .B(_1031__bF_buf65), .C(_3654__12_), .Y(_2151_) );
NOR2X1 NOR2X1_94 ( .A(_2149_), .B(_2143_), .Y(_2152_) );
XNOR2X1 XNOR2X1_38 ( .A(_2152_), .B(bundleStartMajId_i[12]), .Y(_2153_) );
OAI21X1 OAI21X1_630 ( .A(_2153_), .B(_1101__bF_buf34), .C(_2151_), .Y(_534_) );
OAI21X1 OAI21X1_631 ( .A(_1100__bF_buf9_bF_buf3), .B(_1031__bF_buf63), .C(_3654__11_), .Y(_2154_) );
AOI21X1 AOI21X1_19 ( .A(bundleStartMajId_i[12]), .B(_2152_), .C(bundleStartMajId_i[11]), .Y(_2155_) );
NAND2X1 NAND2X1_299 ( .A(_1870_), .B(_1893_), .Y(_2156_) );
OAI21X1 OAI21X1_632 ( .A(_2143_), .B(_2156_), .C(_612__bF_buf4), .Y(_2157_) );
OAI21X1 OAI21X1_633 ( .A(_2155_), .B(_2157_), .C(_2154_), .Y(_535_) );
OAI21X1 OAI21X1_634 ( .A(_1100__bF_buf8_bF_buf0), .B(_1031__bF_buf41), .C(_3654__10_), .Y(_2158_) );
NOR2X1 NOR2X1_95 ( .A(_2156_), .B(_2143_), .Y(_2159_) );
XNOR2X1 XNOR2X1_39 ( .A(_2159_), .B(bundleStartMajId_i[10]), .Y(_2160_) );
OAI21X1 OAI21X1_635 ( .A(_2160_), .B(_1101__bF_buf0), .C(_2158_), .Y(_536_) );
OAI21X1 OAI21X1_636 ( .A(_1100__bF_buf7_bF_buf1), .B(_1031__bF_buf42), .C(_3654__9_), .Y(_2161_) );
AOI21X1 AOI21X1_20 ( .A(bundleStartMajId_i[10]), .B(_2159_), .C(bundleStartMajId_i[9]), .Y(_2162_) );
NAND2X1 NAND2X1_300 ( .A(_1882_), .B(_2159_), .Y(_2163_) );
NAND2X1 NAND2X1_301 ( .A(_612__bF_buf4), .B(_2163_), .Y(_2164_) );
OAI21X1 OAI21X1_637 ( .A(_2164_), .B(_2162_), .C(_2161_), .Y(_537_) );
OAI21X1 OAI21X1_638 ( .A(_1100__bF_buf4), .B(_1031__bF_buf63), .C(_3654__8_), .Y(_2165_) );
AOI21X1 AOI21X1_21 ( .A(_1882_), .B(_2159_), .C(bundleStartMajId_i[8]), .Y(_2166_) );
OAI21X1 OAI21X1_639 ( .A(_2163_), .B(_1598_), .C(_612__bF_buf4), .Y(_2167_) );
OAI21X1 OAI21X1_640 ( .A(_2167_), .B(_2166_), .C(_2165_), .Y(_538_) );
NOR2X1 NOR2X1_96 ( .A(_3654__7_), .B(_612__bF_buf4), .Y(_2168_) );
NAND2X1 NAND2X1_302 ( .A(_1892_), .B(_2159_), .Y(_2169_) );
OR2X2 OR2X2_12 ( .A(_2169_), .B(bundleStartMajId_i[7]), .Y(_2170_) );
AOI21X1 AOI21X1_22 ( .A(bundleStartMajId_i[7]), .B(_2169_), .C(_1101__bF_buf24), .Y(_2171_) );
AOI21X1 AOI21X1_23 ( .A(_2171_), .B(_2170_), .C(_2168_), .Y(_539_) );
OAI21X1 OAI21X1_641 ( .A(_1100__bF_buf9), .B(_1031__bF_buf60), .C(_3654__6_), .Y(_2172_) );
NAND3X1 NAND3X1_25 ( .A(bundleStartMajId_i[8]), .B(bundleStartMajId_i[7]), .C(_1882_), .Y(_2173_) );
OR2X2 OR2X2_13 ( .A(_2173_), .B(_2156_), .Y(_2174_) );
OAI21X1 OAI21X1_642 ( .A(_2143_), .B(_2174_), .C(_1602_), .Y(_2175_) );
NOR2X1 NOR2X1_97 ( .A(_2174_), .B(_2143_), .Y(_2176_) );
NAND2X1 NAND2X1_303 ( .A(bundleStartMajId_i[6]), .B(_2176_), .Y(_2177_) );
NAND2X1 NAND2X1_304 ( .A(_2175_), .B(_2177_), .Y(_2178_) );
OAI21X1 OAI21X1_643 ( .A(_2178_), .B(_1101__bF_buf33), .C(_2172_), .Y(_540_) );
OAI21X1 OAI21X1_644 ( .A(_1100__bF_buf9), .B(_1031__bF_buf60), .C(_3654__5_), .Y(_2179_) );
AOI21X1 AOI21X1_24 ( .A(bundleStartMajId_i[6]), .B(_2176_), .C(bundleStartMajId_i[5]), .Y(_2180_) );
OAI21X1 OAI21X1_645 ( .A(_2177_), .B(_1604_), .C(_612__bF_buf5), .Y(_2181_) );
OAI21X1 OAI21X1_646 ( .A(_2181_), .B(_2180_), .C(_2179_), .Y(_541_) );
AND2X2 AND2X2_16 ( .A(_2176_), .B(_1910_), .Y(_2182_) );
NOR2X1 NOR2X1_98 ( .A(bundleStartMajId_i[4]), .B(_2182_), .Y(_2183_) );
OAI21X1 OAI21X1_647 ( .A(_1100__bF_buf14), .B(_1031__bF_buf2), .C(_3654__4_), .Y(_2184_) );
NAND2X1 NAND2X1_305 ( .A(_1910_), .B(_2176_), .Y(_2185_) );
OAI21X1 OAI21X1_648 ( .A(_2185_), .B(_1606_), .C(_612__bF_buf5), .Y(_2186_) );
OAI21X1 OAI21X1_649 ( .A(_2183_), .B(_2186_), .C(_2184_), .Y(_542_) );
OAI21X1 OAI21X1_650 ( .A(_1100__bF_buf14), .B(_1031__bF_buf32), .C(_3654__3_), .Y(_2187_) );
AOI21X1 AOI21X1_25 ( .A(bundleStartMajId_i[4]), .B(_2182_), .C(bundleStartMajId_i[3]), .Y(_2188_) );
NOR2X1 NOR2X1_99 ( .A(_1608_), .B(_1912_), .Y(_2189_) );
NAND2X1 NAND2X1_306 ( .A(_2189_), .B(_2176_), .Y(_2190_) );
NAND2X1 NAND2X1_307 ( .A(_612__bF_buf5), .B(_2190_), .Y(_2191_) );
OAI21X1 OAI21X1_651 ( .A(_2188_), .B(_2191_), .C(_2187_), .Y(_543_) );
OAI21X1 OAI21X1_652 ( .A(_1100__bF_buf14), .B(_1031__bF_buf2), .C(_3654__2_), .Y(_2192_) );
AND2X2 AND2X2_17 ( .A(_2176_), .B(_2189_), .Y(_2193_) );
NOR2X1 NOR2X1_100 ( .A(bundleStartMajId_i[2]), .B(_2193_), .Y(_2194_) );
OAI21X1 OAI21X1_653 ( .A(_2190_), .B(_1610_), .C(_612__bF_buf5), .Y(_2195_) );
OAI21X1 OAI21X1_654 ( .A(_2194_), .B(_2195_), .C(_2192_), .Y(_544_) );
OAI21X1 OAI21X1_655 ( .A(_1100__bF_buf10), .B(_1031__bF_buf48), .C(_3654__1_), .Y(_2196_) );
AOI21X1 AOI21X1_26 ( .A(bundleStartMajId_i[2]), .B(_2193_), .C(bundleStartMajId_i[1]), .Y(_2197_) );
OAI21X1 OAI21X1_656 ( .A(_2190_), .B(_1928_), .C(_612__bF_buf5), .Y(_2198_) );
OAI21X1 OAI21X1_657 ( .A(_2197_), .B(_2198_), .C(_2196_), .Y(_545_) );
NOR2X1 NOR2X1_101 ( .A(_3654__0_), .B(_612__bF_buf4), .Y(_2199_) );
NAND3X1 NAND3X1_26 ( .A(_1927_), .B(_2189_), .C(_2176_), .Y(_2200_) );
OR2X2 OR2X2_14 ( .A(_2200_), .B(bundleStartMajId_i[0]), .Y(_2201_) );
AOI21X1 AOI21X1_27 ( .A(bundleStartMajId_i[0]), .B(_2200_), .C(_1101__bF_buf23), .Y(_2202_) );
AOI21X1 AOI21X1_28 ( .A(_2202_), .B(_2201_), .C(_2199_), .Y(_546_) );
OAI21X1 OAI21X1_658 ( .A(_1101__bF_buf34), .B(_1135__bF_buf10_bF_buf3), .C(_3655__63_), .Y(_2203_) );
OAI21X1 OAI21X1_659 ( .A(bundleStartMajId_i[63]), .B(_1134__bF_buf13), .C(_2203_), .Y(_547_) );
OAI21X1 OAI21X1_660 ( .A(_1101__bF_buf48), .B(_1135__bF_buf9_bF_buf1), .C(_3655__62_), .Y(_2204_) );
OAI21X1 OAI21X1_661 ( .A(_1134__bF_buf4), .B(_1621_), .C(_2204_), .Y(_548_) );
OAI21X1 OAI21X1_662 ( .A(bundleStartMajId_i[63]), .B(bundleStartMajId_i[62]), .C(bundleStartMajId_i[61]), .Y(_2205_) );
OAI21X1 OAI21X1_663 ( .A(_1936_), .B(bundleStartMajId_i[63]), .C(_2205_), .Y(_2206_) );
OAI21X1 OAI21X1_664 ( .A(_1101__bF_buf3), .B(_1135__bF_buf8_bF_buf1), .C(_3655__61_), .Y(_2207_) );
OAI21X1 OAI21X1_665 ( .A(_2206_), .B(_1134__bF_buf1), .C(_2207_), .Y(_549_) );
OAI21X1 OAI21X1_666 ( .A(_1620_), .B(_1492_), .C(_1494_), .Y(_2208_) );
OAI21X1 OAI21X1_667 ( .A(_1620_), .B(_1627_), .C(_2208_), .Y(_2209_) );
OAI21X1 OAI21X1_668 ( .A(_1101__bF_buf3), .B(_1135__bF_buf7_bF_buf2), .C(_3655__60_), .Y(_2210_) );
OAI21X1 OAI21X1_669 ( .A(_2209_), .B(_1134__bF_buf7), .C(_2210_), .Y(_550_) );
AOI21X1 AOI21X1_29 ( .A(_1488_), .B(_1490_), .C(_1627_), .Y(_2211_) );
XNOR2X1 XNOR2X1_40 ( .A(_2211_), .B(bundleStartMajId_i[59]), .Y(_2212_) );
OAI21X1 OAI21X1_670 ( .A(_1101__bF_buf44), .B(_1135__bF_buf6_bF_buf1), .C(_3655__59_), .Y(_2213_) );
OAI21X1 OAI21X1_671 ( .A(_2212_), .B(_1134__bF_buf1), .C(_2213_), .Y(_551_) );
INVX2 INVX2_52 ( .A(_2211_), .Y(_2214_) );
OAI21X1 OAI21X1_672 ( .A(_2214_), .B(_1496_), .C(_1498_), .Y(_2215_) );
OAI21X1 OAI21X1_673 ( .A(_1637_), .B(_2214_), .C(_2215_), .Y(_2216_) );
OAI21X1 OAI21X1_674 ( .A(_1101__bF_buf6), .B(_1135__bF_buf5_bF_buf0), .C(_3655__58_), .Y(_2217_) );
OAI21X1 OAI21X1_675 ( .A(_2216_), .B(_1134__bF_buf1), .C(_2217_), .Y(_552_) );
NOR2X1 NOR2X1_102 ( .A(_1637_), .B(_2214_), .Y(_2218_) );
INVX1 INVX1_34 ( .A(_2218_), .Y(_2219_) );
NOR2X1 NOR2X1_103 ( .A(_1500_), .B(_2219_), .Y(_2220_) );
INVX8 INVX8_2 ( .A(_1134__bF_buf5), .Y(_613_) );
OAI21X1 OAI21X1_676 ( .A(_2218_), .B(bundleStartMajId_i[57]), .C(_613__bF_buf3), .Y(_2221_) );
OAI21X1 OAI21X1_677 ( .A(_1101__bF_buf16), .B(_1135__bF_buf4_bF_buf0), .C(_3655__57_), .Y(_2222_) );
OAI21X1 OAI21X1_678 ( .A(_2220_), .B(_2221_), .C(_2222_), .Y(_553_) );
OAI21X1 OAI21X1_679 ( .A(_2219_), .B(_1500_), .C(_1502_), .Y(_2223_) );
NAND2X1 NAND2X1_308 ( .A(_2211_), .B(_1647_), .Y(_2224_) );
NAND2X1 NAND2X1_309 ( .A(_2224_), .B(_2223_), .Y(_2225_) );
OAI21X1 OAI21X1_680 ( .A(_1101__bF_buf34), .B(_1135__bF_buf3_bF_buf1), .C(_3655__56_), .Y(_2226_) );
OAI21X1 OAI21X1_681 ( .A(_2225_), .B(_1134__bF_buf13), .C(_2226_), .Y(_554_) );
AND2X2 AND2X2_18 ( .A(_1647_), .B(_2211_), .Y(_2227_) );
NAND2X1 NAND2X1_310 ( .A(bundleStartMajId_i[55]), .B(_2227_), .Y(_2228_) );
NAND2X1 NAND2X1_311 ( .A(_1504_), .B(_2224_), .Y(_2229_) );
NAND2X1 NAND2X1_312 ( .A(_2229_), .B(_2228_), .Y(_2230_) );
OAI21X1 OAI21X1_682 ( .A(_1101__bF_buf12), .B(_1135__bF_buf2_bF_buf1), .C(_3655__55_), .Y(_2231_) );
OAI21X1 OAI21X1_683 ( .A(_2230_), .B(_1134__bF_buf4), .C(_2231_), .Y(_555_) );
XNOR2X1 XNOR2X1_41 ( .A(_2228_), .B(_1506_), .Y(_2232_) );
OAI21X1 OAI21X1_684 ( .A(_1101__bF_buf12), .B(_1135__bF_buf1_bF_buf0), .C(_3655__54_), .Y(_2233_) );
OAI21X1 OAI21X1_685 ( .A(_2232_), .B(_1134__bF_buf4), .C(_2233_), .Y(_556_) );
INVX1 INVX1_35 ( .A(_2228_), .Y(_2234_) );
AOI21X1 AOI21X1_30 ( .A(bundleStartMajId_i[54]), .B(_2234_), .C(bundleStartMajId_i[53]), .Y(_2235_) );
OAI21X1 OAI21X1_686 ( .A(_2228_), .B(_1659_), .C(_613__bF_buf3), .Y(_2236_) );
OAI21X1 OAI21X1_687 ( .A(_1101__bF_buf12), .B(_1135__bF_buf0), .C(_3655__53_), .Y(_2237_) );
OAI21X1 OAI21X1_688 ( .A(_2235_), .B(_2236_), .C(_2237_), .Y(_557_) );
OAI21X1 OAI21X1_689 ( .A(_2228_), .B(_1659_), .C(_1510_), .Y(_2238_) );
OAI21X1 OAI21X1_690 ( .A(_1970_), .B(_2228_), .C(_2238_), .Y(_2239_) );
OAI21X1 OAI21X1_691 ( .A(_1101__bF_buf3), .B(_1135__bF_buf14_bF_buf1), .C(_3655__52_), .Y(_2240_) );
OAI21X1 OAI21X1_692 ( .A(_2239_), .B(_1134__bF_buf1), .C(_2240_), .Y(_558_) );
NOR2X1 NOR2X1_104 ( .A(_1970_), .B(_2228_), .Y(_2241_) );
AND2X2 AND2X2_19 ( .A(_2241_), .B(bundleStartMajId_i[51]), .Y(_2242_) );
OAI21X1 OAI21X1_693 ( .A(_2241_), .B(bundleStartMajId_i[51]), .C(_613__bF_buf3), .Y(_2243_) );
OAI21X1 OAI21X1_694 ( .A(_1101__bF_buf57), .B(_1135__bF_buf13_bF_buf2), .C(_3655__51_), .Y(_2244_) );
OAI21X1 OAI21X1_695 ( .A(_2242_), .B(_2243_), .C(_2244_), .Y(_559_) );
XNOR2X1 XNOR2X1_42 ( .A(_2242_), .B(bundleStartMajId_i[50]), .Y(_2245_) );
OAI21X1 OAI21X1_696 ( .A(_1101__bF_buf12), .B(_1135__bF_buf12_bF_buf2), .C(_3655__50_), .Y(_2246_) );
OAI21X1 OAI21X1_697 ( .A(_2245_), .B(_1134__bF_buf4), .C(_2246_), .Y(_560_) );
AND2X2 AND2X2_20 ( .A(_2242_), .B(bundleStartMajId_i[50]), .Y(_2247_) );
NAND2X1 NAND2X1_313 ( .A(_1981_), .B(_2242_), .Y(_2248_) );
OAI21X1 OAI21X1_698 ( .A(_2247_), .B(bundleStartMajId_i[49]), .C(_2248_), .Y(_2249_) );
OAI21X1 OAI21X1_699 ( .A(_1101__bF_buf12), .B(_1135__bF_buf11_bF_buf1), .C(_3655__49_), .Y(_2250_) );
OAI21X1 OAI21X1_700 ( .A(_2249_), .B(_1134__bF_buf4), .C(_2250_), .Y(_561_) );
NAND2X1 NAND2X1_314 ( .A(_1518_), .B(_2248_), .Y(_2251_) );
OAI21X1 OAI21X1_701 ( .A(_1686_), .B(_2224_), .C(_2251_), .Y(_2252_) );
OAI21X1 OAI21X1_702 ( .A(_1101__bF_buf34), .B(_1135__bF_buf10_bF_buf3), .C(_3655__48_), .Y(_2253_) );
OAI21X1 OAI21X1_703 ( .A(_2252_), .B(_1134__bF_buf13), .C(_2253_), .Y(_562_) );
NOR2X1 NOR2X1_105 ( .A(_2224_), .B(_1686_), .Y(_2254_) );
NAND2X1 NAND2X1_315 ( .A(bundleStartMajId_i[47]), .B(_2254_), .Y(_2255_) );
OAI21X1 OAI21X1_704 ( .A(_1686_), .B(_2224_), .C(_1520_), .Y(_2256_) );
NAND2X1 NAND2X1_316 ( .A(_2256_), .B(_2255_), .Y(_2257_) );
OAI21X1 OAI21X1_705 ( .A(_1101__bF_buf48), .B(_1135__bF_buf9_bF_buf1), .C(_3655__47_), .Y(_2258_) );
OAI21X1 OAI21X1_706 ( .A(_2257_), .B(_1134__bF_buf4), .C(_2258_), .Y(_563_) );
XNOR2X1 XNOR2X1_43 ( .A(_2255_), .B(_1522_), .Y(_2259_) );
OAI21X1 OAI21X1_707 ( .A(_1101__bF_buf4), .B(_1135__bF_buf8_bF_buf2), .C(_3655__46_), .Y(_2260_) );
OAI21X1 OAI21X1_708 ( .A(_2259_), .B(_1134__bF_buf3), .C(_2260_), .Y(_564_) );
INVX1 INVX1_36 ( .A(_2255_), .Y(_2261_) );
AOI21X1 AOI21X1_31 ( .A(bundleStartMajId_i[46]), .B(_2261_), .C(bundleStartMajId_i[45]), .Y(_2262_) );
OAI21X1 OAI21X1_709 ( .A(_2255_), .B(_1694_), .C(_613__bF_buf1), .Y(_2263_) );
OAI21X1 OAI21X1_710 ( .A(_1101__bF_buf4), .B(_1135__bF_buf7_bF_buf0), .C(_3655__45_), .Y(_2264_) );
OAI21X1 OAI21X1_711 ( .A(_2262_), .B(_2263_), .C(_2264_), .Y(_565_) );
OAI21X1 OAI21X1_712 ( .A(_2255_), .B(_1694_), .C(_1526_), .Y(_2265_) );
OAI21X1 OAI21X1_713 ( .A(_1999_), .B(_2255_), .C(_2265_), .Y(_2266_) );
OAI21X1 OAI21X1_714 ( .A(_1101__bF_buf8), .B(_1135__bF_buf6_bF_buf2), .C(_3655__44_), .Y(_2267_) );
OAI21X1 OAI21X1_715 ( .A(_2266_), .B(_1134__bF_buf14), .C(_2267_), .Y(_566_) );
NOR2X1 NOR2X1_106 ( .A(_1999_), .B(_2255_), .Y(_2268_) );
NAND2X1 NAND2X1_317 ( .A(bundleStartMajId_i[43]), .B(_2268_), .Y(_2269_) );
INVX1 INVX1_37 ( .A(_2269_), .Y(_2270_) );
OAI21X1 OAI21X1_716 ( .A(_2268_), .B(bundleStartMajId_i[43]), .C(_613__bF_buf1), .Y(_2271_) );
OAI21X1 OAI21X1_717 ( .A(_1101__bF_buf37), .B(_1135__bF_buf5_bF_buf3), .C(_3655__43_), .Y(_2272_) );
OAI21X1 OAI21X1_718 ( .A(_2270_), .B(_2271_), .C(_2272_), .Y(_567_) );
XNOR2X1 XNOR2X1_44 ( .A(_2269_), .B(_1530_), .Y(_2273_) );
OAI21X1 OAI21X1_719 ( .A(_1101__bF_buf2), .B(_1135__bF_buf4_bF_buf1), .C(_3655__42_), .Y(_2274_) );
OAI21X1 OAI21X1_720 ( .A(_2273_), .B(_1134__bF_buf3), .C(_2274_), .Y(_568_) );
OAI21X1 OAI21X1_721 ( .A(_2269_), .B(_1530_), .C(_1532_), .Y(_2275_) );
OAI21X1 OAI21X1_722 ( .A(_2013_), .B(_2269_), .C(_2275_), .Y(_2276_) );
OAI21X1 OAI21X1_723 ( .A(_1101__bF_buf37), .B(_1135__bF_buf3_bF_buf1), .C(_3655__41_), .Y(_2277_) );
OAI21X1 OAI21X1_724 ( .A(_2276_), .B(_1134__bF_buf3), .C(_2277_), .Y(_569_) );
NAND2X1 NAND2X1_318 ( .A(_2227_), .B(_1711_), .Y(_2278_) );
NOR2X1 NOR2X1_107 ( .A(_1714_), .B(_2278_), .Y(_2279_) );
NAND3X1 NAND3X1_27 ( .A(bundleStartMajId_i[41]), .B(_1716_), .C(_2279_), .Y(_2280_) );
XNOR2X1 XNOR2X1_45 ( .A(_2280_), .B(_1534_), .Y(_2281_) );
OAI21X1 OAI21X1_725 ( .A(_1101__bF_buf2), .B(_1135__bF_buf2_bF_buf1), .C(_3655__40_), .Y(_2282_) );
OAI21X1 OAI21X1_726 ( .A(_2281_), .B(_1134__bF_buf3), .C(_2282_), .Y(_570_) );
NAND2X1 NAND2X1_319 ( .A(_1726_), .B(_2254_), .Y(_2283_) );
NOR2X1 NOR2X1_108 ( .A(_1536_), .B(_2283_), .Y(_2284_) );
INVX1 INVX1_38 ( .A(_2284_), .Y(_2285_) );
OAI21X1 OAI21X1_727 ( .A(_2278_), .B(_1787_), .C(_1536_), .Y(_2286_) );
NAND2X1 NAND2X1_320 ( .A(_2286_), .B(_2285_), .Y(_2287_) );
OAI21X1 OAI21X1_728 ( .A(_1101__bF_buf46), .B(_1135__bF_buf1_bF_buf3), .C(_3655__39_), .Y(_2288_) );
OAI21X1 OAI21X1_729 ( .A(_2287_), .B(_1134__bF_buf8), .C(_2288_), .Y(_571_) );
OAI21X1 OAI21X1_730 ( .A(_2283_), .B(_1536_), .C(_1538_), .Y(_2289_) );
OAI21X1 OAI21X1_731 ( .A(_1736_), .B(_2283_), .C(_2289_), .Y(_2290_) );
OAI21X1 OAI21X1_732 ( .A(_1101__bF_buf46), .B(_1135__bF_buf8), .C(_3655__38_), .Y(_2291_) );
OAI21X1 OAI21X1_733 ( .A(_2290_), .B(_1134__bF_buf8), .C(_2291_), .Y(_572_) );
NOR2X1 NOR2X1_109 ( .A(_1787_), .B(_2278_), .Y(_2292_) );
AOI21X1 AOI21X1_32 ( .A(_1734_), .B(_2292_), .C(bundleStartMajId_i[37]), .Y(_2293_) );
OAI21X1 OAI21X1_734 ( .A(_2285_), .B(_1740_), .C(_613__bF_buf1), .Y(_2294_) );
OAI21X1 OAI21X1_735 ( .A(_1101__bF_buf5), .B(_1135__bF_buf14_bF_buf3), .C(_3655__37_), .Y(_2295_) );
OAI21X1 OAI21X1_736 ( .A(_2294_), .B(_2293_), .C(_2295_), .Y(_573_) );
NAND2X1 NAND2X1_321 ( .A(_1741_), .B(_2284_), .Y(_2296_) );
XNOR2X1 XNOR2X1_46 ( .A(_2296_), .B(_1542_), .Y(_2297_) );
OAI21X1 OAI21X1_737 ( .A(_1101__bF_buf32), .B(_1135__bF_buf13_bF_buf1), .C(_3655__36_), .Y(_2298_) );
OAI21X1 OAI21X1_738 ( .A(_2297_), .B(_1134__bF_buf8), .C(_2298_), .Y(_574_) );
OAI21X1 OAI21X1_739 ( .A(_2296_), .B(_1542_), .C(_1544_), .Y(_2299_) );
NAND2X1 NAND2X1_322 ( .A(_1746_), .B(_2284_), .Y(_2300_) );
NAND2X1 NAND2X1_323 ( .A(_2300_), .B(_2299_), .Y(_2301_) );
OAI21X1 OAI21X1_740 ( .A(_1101__bF_buf4), .B(_1135__bF_buf12_bF_buf3), .C(_3655__35_), .Y(_2302_) );
OAI21X1 OAI21X1_741 ( .A(_2301_), .B(_1134__bF_buf8), .C(_2302_), .Y(_575_) );
XNOR2X1 XNOR2X1_47 ( .A(_2300_), .B(_1546_), .Y(_2303_) );
OAI21X1 OAI21X1_742 ( .A(_1101__bF_buf49), .B(_1135__bF_buf11_bF_buf3), .C(_3655__34_), .Y(_2304_) );
OAI21X1 OAI21X1_743 ( .A(_2303_), .B(_1134__bF_buf8), .C(_2304_), .Y(_576_) );
OAI21X1 OAI21X1_744 ( .A(_1101__bF_buf52), .B(_1135__bF_buf10_bF_buf2), .C(_3655__33_), .Y(_2305_) );
NAND3X1 NAND3X1_28 ( .A(_1788_), .B(_1755_), .C(_2292_), .Y(_2306_) );
XNOR2X1 XNOR2X1_48 ( .A(_2306_), .B(_1548_), .Y(_2307_) );
OAI21X1 OAI21X1_745 ( .A(_2307_), .B(_1134__bF_buf8), .C(_2305_), .Y(_577_) );
INVX1 INVX1_39 ( .A(_3655__32_), .Y(_2308_) );
NOR3X1 NOR3X1_7 ( .A(_1548_), .B(bundleStartMajId_i[32]), .C(_2306_), .Y(_2309_) );
INVX1 INVX1_40 ( .A(_2306_), .Y(_2310_) );
AOI21X1 AOI21X1_33 ( .A(bundleStartMajId_i[33]), .B(_2310_), .C(_1550_), .Y(_2311_) );
OAI21X1 OAI21X1_746 ( .A(_2311_), .B(_2309_), .C(_613__bF_buf1), .Y(_2312_) );
OAI21X1 OAI21X1_747 ( .A(_2308_), .B(_613__bF_buf2), .C(_2312_), .Y(_578_) );
NAND2X1 NAND2X1_324 ( .A(_2254_), .B(_1791_), .Y(_2313_) );
OR2X2 OR2X2_15 ( .A(_2313_), .B(_1552_), .Y(_2314_) );
OAI21X1 OAI21X1_748 ( .A(_1768_), .B(_2278_), .C(_1552_), .Y(_2315_) );
NAND2X1 NAND2X1_325 ( .A(_2315_), .B(_2314_), .Y(_2316_) );
OAI21X1 OAI21X1_749 ( .A(_1101__bF_buf24), .B(_1135__bF_buf9_bF_buf1), .C(_3655__31_), .Y(_2317_) );
OAI21X1 OAI21X1_750 ( .A(_2316_), .B(_1134__bF_buf4), .C(_2317_), .Y(_579_) );
OAI21X1 OAI21X1_751 ( .A(_2313_), .B(_1552_), .C(_1554_), .Y(_2318_) );
OAI21X1 OAI21X1_752 ( .A(_1780_), .B(_2313_), .C(_2318_), .Y(_2319_) );
OAI21X1 OAI21X1_753 ( .A(_1101__bF_buf2), .B(_1135__bF_buf8_bF_buf2), .C(_3655__30_), .Y(_2320_) );
OAI21X1 OAI21X1_754 ( .A(_2319_), .B(_1134__bF_buf3), .C(_2320_), .Y(_580_) );
NOR2X1 NOR2X1_110 ( .A(_1780_), .B(_2313_), .Y(_2321_) );
NAND2X1 NAND2X1_326 ( .A(bundleStartMajId_i[29]), .B(_2321_), .Y(_2322_) );
INVX1 INVX1_41 ( .A(_2322_), .Y(_2323_) );
OAI21X1 OAI21X1_755 ( .A(_2321_), .B(bundleStartMajId_i[29]), .C(_613__bF_buf3), .Y(_2324_) );
OAI21X1 OAI21X1_756 ( .A(_1101__bF_buf37), .B(_1135__bF_buf7_bF_buf0), .C(_3655__29_), .Y(_2325_) );
OAI21X1 OAI21X1_757 ( .A(_2323_), .B(_2324_), .C(_2325_), .Y(_581_) );
XNOR2X1 XNOR2X1_49 ( .A(_2322_), .B(_1558_), .Y(_2326_) );
OAI21X1 OAI21X1_758 ( .A(_1101__bF_buf8), .B(_1135__bF_buf6_bF_buf2), .C(_3655__28_), .Y(_2327_) );
OAI21X1 OAI21X1_759 ( .A(_2326_), .B(_1134__bF_buf3), .C(_2327_), .Y(_582_) );
OAI21X1 OAI21X1_760 ( .A(_2322_), .B(_1558_), .C(_1560_), .Y(_2328_) );
OAI21X1 OAI21X1_761 ( .A(_2074_), .B(_2314_), .C(_2328_), .Y(_2329_) );
OAI21X1 OAI21X1_762 ( .A(_1101__bF_buf37), .B(_1135__bF_buf5_bF_buf3), .C(_3655__27_), .Y(_2330_) );
OAI21X1 OAI21X1_763 ( .A(_2329_), .B(_1134__bF_buf3), .C(_2330_), .Y(_583_) );
NAND3X1 NAND3X1_29 ( .A(_1793_), .B(_2254_), .C(_1791_), .Y(_2331_) );
NOR2X1 NOR2X1_111 ( .A(_1560_), .B(_2331_), .Y(_2332_) );
XNOR2X1 XNOR2X1_50 ( .A(_2332_), .B(bundleStartMajId_i[26]), .Y(_2333_) );
OAI21X1 OAI21X1_764 ( .A(_1101__bF_buf52), .B(_1135__bF_buf4_bF_buf1), .C(_3655__26_), .Y(_2334_) );
OAI21X1 OAI21X1_765 ( .A(_2333_), .B(_1134__bF_buf12), .C(_2334_), .Y(_584_) );
INVX1 INVX1_42 ( .A(_3655__25_), .Y(_2335_) );
NOR2X1 NOR2X1_112 ( .A(_1800_), .B(_2331_), .Y(_2336_) );
NOR2X1 NOR2X1_113 ( .A(_1564_), .B(_2336_), .Y(_2337_) );
AND2X2 AND2X2_21 ( .A(_2336_), .B(_1564_), .Y(_2338_) );
OAI21X1 OAI21X1_766 ( .A(_2338_), .B(_2337_), .C(_613__bF_buf1), .Y(_2339_) );
OAI21X1 OAI21X1_767 ( .A(_2335_), .B(_613__bF_buf1), .C(_2339_), .Y(_585_) );
NAND2X1 NAND2X1_327 ( .A(bundleStartMajId_i[25]), .B(_2336_), .Y(_2340_) );
XNOR2X1 XNOR2X1_51 ( .A(_2340_), .B(_1566_), .Y(_2341_) );
OAI21X1 OAI21X1_768 ( .A(_1101__bF_buf37), .B(_1135__bF_buf3_bF_buf1), .C(_3655__24_), .Y(_2342_) );
OAI21X1 OAI21X1_769 ( .A(_2341_), .B(_1134__bF_buf3), .C(_2342_), .Y(_586_) );
NAND3X1 NAND3X1_30 ( .A(_1809_), .B(_2254_), .C(_1791_), .Y(_2343_) );
NOR2X1 NOR2X1_114 ( .A(_1568_), .B(_2343_), .Y(_2344_) );
INVX4 INVX4_31 ( .A(_2344_), .Y(_2345_) );
OAI21X1 OAI21X1_770 ( .A(_2313_), .B(_1848_), .C(_1568_), .Y(_2346_) );
NAND2X1 NAND2X1_328 ( .A(_2346_), .B(_2345_), .Y(_2347_) );
OAI21X1 OAI21X1_771 ( .A(_1101__bF_buf4), .B(_1135__bF_buf2_bF_buf3), .C(_3655__23_), .Y(_2348_) );
OAI21X1 OAI21X1_772 ( .A(_2347_), .B(_1134__bF_buf3), .C(_2348_), .Y(_587_) );
XNOR2X1 XNOR2X1_52 ( .A(_2344_), .B(bundleStartMajId_i[22]), .Y(_2349_) );
OAI21X1 OAI21X1_773 ( .A(_1101__bF_buf57), .B(_1135__bF_buf1_bF_buf1), .C(_3655__22_), .Y(_2350_) );
OAI21X1 OAI21X1_774 ( .A(_2349_), .B(_1134__bF_buf4), .C(_2350_), .Y(_588_) );
OAI21X1 OAI21X1_775 ( .A(_2345_), .B(_1570_), .C(_1572_), .Y(_2351_) );
OAI21X1 OAI21X1_776 ( .A(_1827_), .B(_2343_), .C(_2351_), .Y(_2352_) );
OAI21X1 OAI21X1_777 ( .A(_1101__bF_buf44), .B(_1135__bF_buf9), .C(_3655__21_), .Y(_2353_) );
OAI21X1 OAI21X1_778 ( .A(_2352_), .B(_1134__bF_buf4), .C(_2353_), .Y(_589_) );
OAI21X1 OAI21X1_779 ( .A(_2343_), .B(_1827_), .C(_1574_), .Y(_2354_) );
OAI21X1 OAI21X1_780 ( .A(_1829_), .B(_2343_), .C(_2354_), .Y(_2355_) );
OAI21X1 OAI21X1_781 ( .A(_1101__bF_buf18), .B(_1135__bF_buf14_bF_buf0), .C(_3655__20_), .Y(_2356_) );
OAI21X1 OAI21X1_782 ( .A(_2355_), .B(_1134__bF_buf14), .C(_2356_), .Y(_590_) );
OAI21X1 OAI21X1_783 ( .A(_2343_), .B(_1829_), .C(_1576_), .Y(_2357_) );
OAI21X1 OAI21X1_784 ( .A(_2345_), .B(_2122_), .C(_2357_), .Y(_2358_) );
OAI21X1 OAI21X1_785 ( .A(_1101__bF_buf34), .B(_1135__bF_buf13_bF_buf2), .C(_3655__19_), .Y(_2359_) );
OAI21X1 OAI21X1_786 ( .A(_2358_), .B(_1134__bF_buf4), .C(_2359_), .Y(_591_) );
OAI21X1 OAI21X1_787 ( .A(_2345_), .B(_2122_), .C(_1578_), .Y(_2360_) );
NAND3X1 NAND3X1_31 ( .A(bundleStartMajId_i[18]), .B(_2121_), .C(_2344_), .Y(_2361_) );
NAND2X1 NAND2X1_329 ( .A(_2361_), .B(_2360_), .Y(_2362_) );
OAI21X1 OAI21X1_788 ( .A(_1101__bF_buf37), .B(_1135__bF_buf12_bF_buf0), .C(_3655__18_), .Y(_2363_) );
OAI21X1 OAI21X1_789 ( .A(_2362_), .B(_1134__bF_buf3), .C(_2363_), .Y(_592_) );
OAI21X1 OAI21X1_790 ( .A(_1101__bF_buf57), .B(_1135__bF_buf11_bF_buf1), .C(_3655__17_), .Y(_2364_) );
AND2X2 AND2X2_22 ( .A(_2361_), .B(_1580_), .Y(_2365_) );
NAND2X1 NAND2X1_330 ( .A(_1837_), .B(_2121_), .Y(_2366_) );
OAI21X1 OAI21X1_791 ( .A(_2345_), .B(_2366_), .C(_613__bF_buf3), .Y(_2367_) );
OAI21X1 OAI21X1_792 ( .A(_2365_), .B(_2367_), .C(_2364_), .Y(_593_) );
OAI21X1 OAI21X1_793 ( .A(_2345_), .B(_2366_), .C(_1582_), .Y(_2368_) );
OAI21X1 OAI21X1_794 ( .A(_1846_), .B(_2313_), .C(_2368_), .Y(_2369_) );
OAI21X1 OAI21X1_795 ( .A(_1101__bF_buf18), .B(_1135__bF_buf10_bF_buf3), .C(_3655__16_), .Y(_2370_) );
OAI21X1 OAI21X1_796 ( .A(_2369_), .B(_1134__bF_buf14), .C(_2370_), .Y(_594_) );
NAND3X1 NAND3X1_32 ( .A(_2254_), .B(_1852_), .C(_1791_), .Y(_2371_) );
NOR2X1 NOR2X1_115 ( .A(_1584_), .B(_2371_), .Y(_2372_) );
INVX2 INVX2_53 ( .A(_2372_), .Y(_2373_) );
OAI21X1 OAI21X1_797 ( .A(_2313_), .B(_1846_), .C(_1584_), .Y(_2374_) );
NAND2X1 NAND2X1_331 ( .A(_2374_), .B(_2373_), .Y(_2375_) );
OAI21X1 OAI21X1_798 ( .A(_1101__bF_buf18), .B(_1135__bF_buf9_bF_buf0), .C(_3655__15_), .Y(_2376_) );
OAI21X1 OAI21X1_799 ( .A(_2375_), .B(_1134__bF_buf13), .C(_2376_), .Y(_595_) );
XNOR2X1 XNOR2X1_53 ( .A(_2372_), .B(bundleStartMajId_i[14]), .Y(_2377_) );
OAI21X1 OAI21X1_800 ( .A(_1101__bF_buf24), .B(_1135__bF_buf8_bF_buf1), .C(_3655__14_), .Y(_2378_) );
OAI21X1 OAI21X1_801 ( .A(_2377_), .B(_1134__bF_buf4), .C(_2378_), .Y(_596_) );
OAI21X1 OAI21X1_802 ( .A(_2373_), .B(_1586_), .C(_1588_), .Y(_2379_) );
OAI21X1 OAI21X1_803 ( .A(_2149_), .B(_2373_), .C(_2379_), .Y(_2380_) );
OAI21X1 OAI21X1_804 ( .A(_1101__bF_buf18), .B(_1135__bF_buf7_bF_buf2), .C(_3655__13_), .Y(_2381_) );
OAI21X1 OAI21X1_805 ( .A(_2380_), .B(_1134__bF_buf13), .C(_2381_), .Y(_597_) );
OAI21X1 OAI21X1_806 ( .A(_2371_), .B(_1871_), .C(_1590_), .Y(_2382_) );
OAI21X1 OAI21X1_807 ( .A(_1873_), .B(_2371_), .C(_2382_), .Y(_2383_) );
OAI21X1 OAI21X1_808 ( .A(_1101__bF_buf23), .B(_1135__bF_buf6_bF_buf2), .C(_3655__12_), .Y(_2384_) );
OAI21X1 OAI21X1_809 ( .A(_2383_), .B(_1134__bF_buf14), .C(_2384_), .Y(_598_) );
OAI21X1 OAI21X1_810 ( .A(_2371_), .B(_1873_), .C(_1592_), .Y(_2385_) );
OAI21X1 OAI21X1_811 ( .A(_2373_), .B(_2156_), .C(_2385_), .Y(_2386_) );
OAI21X1 OAI21X1_812 ( .A(_1101__bF_buf18), .B(_1135__bF_buf5_bF_buf3), .C(_3655__11_), .Y(_2387_) );
OAI21X1 OAI21X1_813 ( .A(_2386_), .B(_1134__bF_buf14), .C(_2387_), .Y(_599_) );
NOR3X1 NOR3X1_8 ( .A(_1592_), .B(_1873_), .C(_2371_), .Y(_2388_) );
XNOR2X1 XNOR2X1_54 ( .A(_2388_), .B(bundleStartMajId_i[10]), .Y(_2389_) );
OAI21X1 OAI21X1_814 ( .A(_1101__bF_buf37), .B(_1135__bF_buf4_bF_buf1), .C(_3655__10_), .Y(_2390_) );
OAI21X1 OAI21X1_815 ( .A(_2389_), .B(_1134__bF_buf3), .C(_2390_), .Y(_600_) );
AOI21X1 AOI21X1_34 ( .A(bundleStartMajId_i[10]), .B(_2388_), .C(bundleStartMajId_i[9]), .Y(_2391_) );
OAI21X1 OAI21X1_816 ( .A(_1101__bF_buf24), .B(_1135__bF_buf3_bF_buf1), .C(_3655__9_), .Y(_2392_) );
NOR3X1 NOR3X1_9 ( .A(_2278_), .B(_1846_), .C(_1768_), .Y(_2393_) );
NAND3X1 NAND3X1_33 ( .A(_1872_), .B(_1893_), .C(_2393_), .Y(_2394_) );
OAI21X1 OAI21X1_817 ( .A(_2394_), .B(_1883_), .C(_613__bF_buf3), .Y(_2395_) );
OAI21X1 OAI21X1_818 ( .A(_2395_), .B(_2391_), .C(_2392_), .Y(_601_) );
OAI21X1 OAI21X1_819 ( .A(_1101__bF_buf46), .B(_1135__bF_buf2_bF_buf3), .C(_3655__8_), .Y(_2396_) );
OAI21X1 OAI21X1_820 ( .A(_2394_), .B(_1883_), .C(_1598_), .Y(_2397_) );
NAND3X1 NAND3X1_34 ( .A(bundleStartMajId_i[8]), .B(_1882_), .C(_2388_), .Y(_2398_) );
NAND2X1 NAND2X1_332 ( .A(_2398_), .B(_2397_), .Y(_2399_) );
OAI21X1 OAI21X1_821 ( .A(_2399_), .B(_1134__bF_buf8), .C(_2396_), .Y(_602_) );
NAND3X1 NAND3X1_35 ( .A(bundleStartMajId_i[7]), .B(_1902_), .C(_2393_), .Y(_2400_) );
OAI21X1 OAI21X1_822 ( .A(_2371_), .B(_1894_), .C(_1600_), .Y(_2401_) );
NAND2X1 NAND2X1_333 ( .A(_2401_), .B(_2400_), .Y(_2402_) );
OAI21X1 OAI21X1_823 ( .A(_1101__bF_buf52), .B(_1135__bF_buf1_bF_buf3), .C(_3655__7_), .Y(_2403_) );
OAI21X1 OAI21X1_824 ( .A(_2402_), .B(_1134__bF_buf8), .C(_2403_), .Y(_603_) );
XNOR2X1 XNOR2X1_55 ( .A(_2400_), .B(_1602_), .Y(_2404_) );
OAI21X1 OAI21X1_825 ( .A(_1101__bF_buf8), .B(_1135__bF_buf2), .C(_3655__6_), .Y(_2405_) );
OAI21X1 OAI21X1_826 ( .A(_2404_), .B(_1134__bF_buf14), .C(_2405_), .Y(_604_) );
INVX1 INVX1_43 ( .A(_1910_), .Y(_2406_) );
OAI21X1 OAI21X1_827 ( .A(_2400_), .B(_1602_), .C(_1604_), .Y(_2407_) );
OAI21X1 OAI21X1_828 ( .A(_2406_), .B(_2400_), .C(_2407_), .Y(_2408_) );
OAI21X1 OAI21X1_829 ( .A(_1101__bF_buf23), .B(_1135__bF_buf14_bF_buf0), .C(_3655__5_), .Y(_2409_) );
OAI21X1 OAI21X1_830 ( .A(_2408_), .B(_1134__bF_buf14), .C(_2409_), .Y(_605_) );
OAI21X1 OAI21X1_831 ( .A(_1101__bF_buf8), .B(_1135__bF_buf13_bF_buf1), .C(_3655__4_), .Y(_2410_) );
NOR2X1 NOR2X1_116 ( .A(_2406_), .B(_2400_), .Y(_2411_) );
NOR2X1 NOR2X1_117 ( .A(bundleStartMajId_i[4]), .B(_2411_), .Y(_2412_) );
NAND3X1 NAND3X1_36 ( .A(_1902_), .B(_1915_), .C(_2393_), .Y(_2413_) );
NAND2X1 NAND2X1_334 ( .A(_613__bF_buf0), .B(_2413_), .Y(_2414_) );
OAI21X1 OAI21X1_832 ( .A(_2412_), .B(_2414_), .C(_2410_), .Y(_606_) );
INVX1 INVX1_44 ( .A(_1915_), .Y(_2415_) );
NOR3X1 NOR3X1_10 ( .A(_1894_), .B(_2415_), .C(_2371_), .Y(_2416_) );
NAND2X1 NAND2X1_335 ( .A(bundleStartMajId_i[3]), .B(_2416_), .Y(_2417_) );
NAND2X1 NAND2X1_336 ( .A(_1608_), .B(_2413_), .Y(_2418_) );
NAND2X1 NAND2X1_337 ( .A(_2417_), .B(_2418_), .Y(_2419_) );
OAI21X1 OAI21X1_833 ( .A(_1101__bF_buf2), .B(_1135__bF_buf12_bF_buf0), .C(_3655__3_), .Y(_2420_) );
OAI21X1 OAI21X1_834 ( .A(_2419_), .B(_1134__bF_buf4), .C(_2420_), .Y(_607_) );
OAI21X1 OAI21X1_835 ( .A(_1101__bF_buf23), .B(_1135__bF_buf11_bF_buf0), .C(_3655__2_), .Y(_2421_) );
NOR2X1 NOR2X1_118 ( .A(_1608_), .B(_2413_), .Y(_2422_) );
NOR2X1 NOR2X1_119 ( .A(bundleStartMajId_i[2]), .B(_2422_), .Y(_2423_) );
OAI21X1 OAI21X1_836 ( .A(_2417_), .B(_1610_), .C(_613__bF_buf0), .Y(_2424_) );
OAI21X1 OAI21X1_837 ( .A(_2423_), .B(_2424_), .C(_2421_), .Y(_608_) );
OAI21X1 OAI21X1_838 ( .A(_1101__bF_buf23), .B(_1135__bF_buf10_bF_buf3), .C(_3655__1_), .Y(_2425_) );
AOI21X1 AOI21X1_35 ( .A(bundleStartMajId_i[2]), .B(_2422_), .C(bundleStartMajId_i[1]), .Y(_2426_) );
OAI21X1 OAI21X1_839 ( .A(_2417_), .B(_1928_), .C(_613__bF_buf0), .Y(_2427_) );
OAI21X1 OAI21X1_840 ( .A(_2426_), .B(_2427_), .C(_2425_), .Y(_609_) );
OAI21X1 OAI21X1_841 ( .A(_1101__bF_buf24), .B(_1135__bF_buf9_bF_buf1), .C(_3655__0_), .Y(_2428_) );
NAND3X1 NAND3X1_37 ( .A(bundleStartMajId_i[3]), .B(_1927_), .C(_2416_), .Y(_2429_) );
NOR2X1 NOR2X1_120 ( .A(_1614_), .B(_2429_), .Y(_2430_) );
NOR3X1 NOR3X1_11 ( .A(_1608_), .B(_1928_), .C(_2413_), .Y(_2431_) );
OAI21X1 OAI21X1_842 ( .A(_2431_), .B(bundleStartMajId_i[0]), .C(_613__bF_buf0), .Y(_2432_) );
OAI21X1 OAI21X1_843 ( .A(_2432_), .B(_2430_), .C(_2428_), .Y(_610_) );
INVX1 INVX1_45 ( .A(_3644__31_), .Y(_2433_) );
NAND2X1 NAND2X1_338 ( .A(enable_i_bF_buf4), .B(bundle_i[31]), .Y(_2434_) );
OAI21X1 OAI21X1_844 ( .A(_2433_), .B(enable_i_bF_buf4), .C(_2434_), .Y(_614_) );
INVX1 INVX1_46 ( .A(_3644__30_), .Y(_2435_) );
NAND2X1 NAND2X1_339 ( .A(enable_i_bF_buf0), .B(bundle_i[30]), .Y(_2436_) );
OAI21X1 OAI21X1_845 ( .A(_2435_), .B(enable_i_bF_buf3), .C(_2436_), .Y(_615_) );
INVX1 INVX1_47 ( .A(_3644__29_), .Y(_2437_) );
NAND2X1 NAND2X1_340 ( .A(enable_i_bF_buf1), .B(bundle_i[29]), .Y(_2438_) );
OAI21X1 OAI21X1_846 ( .A(_2437_), .B(enable_i_bF_buf1), .C(_2438_), .Y(_616_) );
INVX1 INVX1_48 ( .A(_3644__28_), .Y(_2439_) );
NAND2X1 NAND2X1_341 ( .A(enable_i_bF_buf2), .B(bundle_i[28]), .Y(_2440_) );
OAI21X1 OAI21X1_847 ( .A(_2439_), .B(enable_i_bF_buf2), .C(_2440_), .Y(_617_) );
INVX1 INVX1_49 ( .A(_3644__27_), .Y(_2441_) );
NAND2X1 NAND2X1_342 ( .A(enable_i_bF_buf0), .B(bundle_i[27]), .Y(_2442_) );
OAI21X1 OAI21X1_848 ( .A(_2441_), .B(enable_i_bF_buf6), .C(_2442_), .Y(_618_) );
INVX1 INVX1_50 ( .A(_3644__26_), .Y(_2443_) );
NAND2X1 NAND2X1_343 ( .A(enable_i_bF_buf3), .B(bundle_i[26]), .Y(_2444_) );
OAI21X1 OAI21X1_849 ( .A(_2443_), .B(enable_i_bF_buf3), .C(_2444_), .Y(_619_) );
INVX1 INVX1_51 ( .A(_3644__25_), .Y(_2445_) );
NAND2X1 NAND2X1_344 ( .A(enable_i_bF_buf2), .B(bundle_i[25]), .Y(_2446_) );
OAI21X1 OAI21X1_850 ( .A(_2445_), .B(enable_i_bF_buf2), .C(_2446_), .Y(_620_) );
INVX1 INVX1_52 ( .A(_3644__24_), .Y(_2447_) );
NAND2X1 NAND2X1_345 ( .A(enable_i_bF_buf7), .B(bundle_i[24]), .Y(_2448_) );
OAI21X1 OAI21X1_851 ( .A(_2447_), .B(enable_i_bF_buf7), .C(_2448_), .Y(_621_) );
INVX1 INVX1_53 ( .A(_3644__23_), .Y(_2449_) );
NAND2X1 NAND2X1_346 ( .A(enable_i_bF_buf5), .B(bundle_i[23]), .Y(_2450_) );
OAI21X1 OAI21X1_852 ( .A(_2449_), .B(enable_i_bF_buf3), .C(_2450_), .Y(_622_) );
INVX1 INVX1_54 ( .A(_3644__22_), .Y(_2451_) );
NAND2X1 NAND2X1_347 ( .A(enable_i_bF_buf6), .B(bundle_i[22]), .Y(_2452_) );
OAI21X1 OAI21X1_853 ( .A(_2451_), .B(enable_i_bF_buf2), .C(_2452_), .Y(_623_) );
INVX1 INVX1_55 ( .A(_3644__21_), .Y(_2453_) );
NAND2X1 NAND2X1_348 ( .A(enable_i_bF_buf0), .B(bundle_i[21]), .Y(_2454_) );
OAI21X1 OAI21X1_854 ( .A(_2453_), .B(enable_i_bF_buf0), .C(_2454_), .Y(_624_) );
INVX1 INVX1_56 ( .A(_3644__20_), .Y(_2455_) );
NAND2X1 NAND2X1_349 ( .A(enable_i_bF_buf1), .B(bundle_i[20]), .Y(_2456_) );
OAI21X1 OAI21X1_855 ( .A(_2455_), .B(enable_i_bF_buf1), .C(_2456_), .Y(_625_) );
INVX1 INVX1_57 ( .A(_3644__19_), .Y(_2457_) );
NAND2X1 NAND2X1_350 ( .A(enable_i_bF_buf4), .B(bundle_i[19]), .Y(_2458_) );
OAI21X1 OAI21X1_856 ( .A(_2457_), .B(enable_i_bF_buf4), .C(_2458_), .Y(_626_) );
INVX1 INVX1_58 ( .A(_3644__18_), .Y(_2459_) );
NAND2X1 NAND2X1_351 ( .A(enable_i_bF_buf7), .B(bundle_i[18]), .Y(_2460_) );
OAI21X1 OAI21X1_857 ( .A(_2459_), .B(enable_i_bF_buf7), .C(_2460_), .Y(_627_) );
INVX1 INVX1_59 ( .A(_3644__17_), .Y(_2461_) );
NAND2X1 NAND2X1_352 ( .A(enable_i_bF_buf5), .B(bundle_i[17]), .Y(_2462_) );
OAI21X1 OAI21X1_858 ( .A(_2461_), .B(enable_i_bF_buf5), .C(_2462_), .Y(_628_) );
INVX1 INVX1_60 ( .A(_3644__16_), .Y(_2463_) );
NAND2X1 NAND2X1_353 ( .A(enable_i_bF_buf6), .B(bundle_i[16]), .Y(_2464_) );
OAI21X1 OAI21X1_859 ( .A(_2463_), .B(enable_i_bF_buf6), .C(_2464_), .Y(_629_) );
INVX1 INVX1_61 ( .A(_3644__15_), .Y(_2465_) );
NAND2X1 NAND2X1_354 ( .A(enable_i_bF_buf3), .B(bundle_i[15]), .Y(_2466_) );
OAI21X1 OAI21X1_860 ( .A(_2465_), .B(enable_i_bF_buf3), .C(_2466_), .Y(_630_) );
INVX1 INVX1_62 ( .A(_3644__14_), .Y(_2467_) );
NAND2X1 NAND2X1_355 ( .A(enable_i_bF_buf3), .B(bundle_i[14]), .Y(_2468_) );
OAI21X1 OAI21X1_861 ( .A(_2467_), .B(enable_i_bF_buf3), .C(_2468_), .Y(_631_) );
INVX1 INVX1_63 ( .A(_3644__13_), .Y(_2469_) );
NAND2X1 NAND2X1_356 ( .A(enable_i_bF_buf2), .B(bundle_i[13]), .Y(_2470_) );
OAI21X1 OAI21X1_862 ( .A(_2469_), .B(enable_i_bF_buf1), .C(_2470_), .Y(_632_) );
INVX1 INVX1_64 ( .A(_3644__12_), .Y(_2471_) );
NAND2X1 NAND2X1_357 ( .A(enable_i_bF_buf7), .B(bundle_i[12]), .Y(_2472_) );
OAI21X1 OAI21X1_863 ( .A(_2471_), .B(enable_i_bF_buf1), .C(_2472_), .Y(_633_) );
INVX1 INVX1_65 ( .A(_3644__11_), .Y(_2473_) );
NAND2X1 NAND2X1_358 ( .A(enable_i_bF_buf5), .B(bundle_i[11]), .Y(_2474_) );
OAI21X1 OAI21X1_864 ( .A(_2473_), .B(enable_i_bF_buf5), .C(_2474_), .Y(_634_) );
INVX1 INVX1_66 ( .A(_3644__10_), .Y(_2475_) );
NAND2X1 NAND2X1_359 ( .A(enable_i_bF_buf6), .B(bundle_i[10]), .Y(_2476_) );
OAI21X1 OAI21X1_865 ( .A(_2475_), .B(enable_i_bF_buf6), .C(_2476_), .Y(_635_) );
INVX1 INVX1_67 ( .A(_3644__9_), .Y(_2477_) );
NAND2X1 NAND2X1_360 ( .A(enable_i_bF_buf7), .B(bundle_i[9]), .Y(_2478_) );
OAI21X1 OAI21X1_866 ( .A(_2477_), .B(enable_i_bF_buf7), .C(_2478_), .Y(_636_) );
INVX1 INVX1_68 ( .A(_3644__8_), .Y(_2479_) );
NAND2X1 NAND2X1_361 ( .A(enable_i_bF_buf5), .B(bundle_i[8]), .Y(_2480_) );
OAI21X1 OAI21X1_867 ( .A(_2479_), .B(enable_i_bF_buf5), .C(_2480_), .Y(_637_) );
INVX1 INVX1_69 ( .A(_3644__7_), .Y(_2481_) );
NAND2X1 NAND2X1_362 ( .A(enable_i_bF_buf1), .B(bundle_i[7]), .Y(_2482_) );
OAI21X1 OAI21X1_868 ( .A(_2481_), .B(enable_i_bF_buf1), .C(_2482_), .Y(_638_) );
INVX1 INVX1_70 ( .A(_3644__6_), .Y(_2483_) );
NAND2X1 NAND2X1_363 ( .A(enable_i_bF_buf4), .B(bundle_i[6]), .Y(_2484_) );
OAI21X1 OAI21X1_869 ( .A(_2483_), .B(enable_i_bF_buf4), .C(_2484_), .Y(_639_) );
INVX1 INVX1_71 ( .A(_3644__5_), .Y(_2485_) );
NAND2X1 NAND2X1_364 ( .A(enable_i_bF_buf7), .B(bundle_i[5]), .Y(_2486_) );
OAI21X1 OAI21X1_870 ( .A(_2485_), .B(enable_i_bF_buf7), .C(_2486_), .Y(_640_) );
INVX1 INVX1_72 ( .A(_3644__4_), .Y(_2487_) );
NAND2X1 NAND2X1_365 ( .A(enable_i_bF_buf4), .B(bundle_i[4]), .Y(_2488_) );
OAI21X1 OAI21X1_871 ( .A(_2487_), .B(enable_i_bF_buf4), .C(_2488_), .Y(_641_) );
INVX1 INVX1_73 ( .A(_3644__3_), .Y(_2489_) );
NAND2X1 NAND2X1_366 ( .A(enable_i_bF_buf6), .B(bundle_i[3]), .Y(_2490_) );
OAI21X1 OAI21X1_872 ( .A(_2489_), .B(enable_i_bF_buf6), .C(_2490_), .Y(_642_) );
INVX1 INVX1_74 ( .A(_3644__2_), .Y(_2491_) );
NAND2X1 NAND2X1_367 ( .A(enable_i_bF_buf5), .B(bundle_i[2]), .Y(_2492_) );
OAI21X1 OAI21X1_873 ( .A(_2491_), .B(enable_i_bF_buf5), .C(_2492_), .Y(_643_) );
INVX1 INVX1_75 ( .A(_3644__1_), .Y(_2493_) );
NAND2X1 NAND2X1_368 ( .A(enable_i_bF_buf0), .B(bundle_i[1]), .Y(_2494_) );
OAI21X1 OAI21X1_874 ( .A(_2493_), .B(enable_i_bF_buf0), .C(_2494_), .Y(_644_) );
INVX1 INVX1_76 ( .A(_3644__0_), .Y(_2495_) );
NAND2X1 NAND2X1_369 ( .A(enable_i_bF_buf0), .B(bundle_i[0]), .Y(_2496_) );
OAI21X1 OAI21X1_875 ( .A(_2495_), .B(enable_i_bF_buf0), .C(_2496_), .Y(_645_) );
INVX1 INVX1_77 ( .A(bundle_i[63]), .Y(_2497_) );
NAND2X1 NAND2X1_370 ( .A(_3645__31_), .B(_1039__bF_buf57), .Y(_2498_) );
OAI21X1 OAI21X1_876 ( .A(_2497_), .B(_1039__bF_buf57), .C(_2498_), .Y(_646_) );
INVX1 INVX1_78 ( .A(bundle_i[62]), .Y(_2499_) );
NAND2X1 NAND2X1_371 ( .A(_3645__30_), .B(_1039__bF_buf26), .Y(_2500_) );
OAI21X1 OAI21X1_877 ( .A(_2499_), .B(_1039__bF_buf26), .C(_2500_), .Y(_647_) );
INVX1 INVX1_79 ( .A(bundle_i[61]), .Y(_2501_) );
NAND2X1 NAND2X1_372 ( .A(_3645__29_), .B(_1039__bF_buf26), .Y(_2502_) );
OAI21X1 OAI21X1_878 ( .A(_2501_), .B(_1039__bF_buf26), .C(_2502_), .Y(_648_) );
INVX1 INVX1_80 ( .A(bundle_i[60]), .Y(_2503_) );
NAND2X1 NAND2X1_373 ( .A(_3645__28_), .B(_1039__bF_buf32), .Y(_2504_) );
OAI21X1 OAI21X1_879 ( .A(_2503_), .B(_1039__bF_buf32), .C(_2504_), .Y(_649_) );
INVX1 INVX1_81 ( .A(bundle_i[59]), .Y(_2505_) );
NAND2X1 NAND2X1_374 ( .A(_3645__27_), .B(_1039__bF_buf20), .Y(_2506_) );
OAI21X1 OAI21X1_880 ( .A(_2505_), .B(_1039__bF_buf20), .C(_2506_), .Y(_650_) );
INVX1 INVX1_82 ( .A(bundle_i[58]), .Y(_2507_) );
NAND2X1 NAND2X1_375 ( .A(_3645__26_), .B(_1039__bF_buf31), .Y(_2508_) );
OAI21X1 OAI21X1_881 ( .A(_2507_), .B(_1039__bF_buf31), .C(_2508_), .Y(_651_) );
INVX1 INVX1_83 ( .A(bundle_i[57]), .Y(_2509_) );
NAND2X1 NAND2X1_376 ( .A(_3645__25_), .B(_1039__bF_buf32), .Y(_2510_) );
OAI21X1 OAI21X1_882 ( .A(_2509_), .B(_1039__bF_buf32), .C(_2510_), .Y(_652_) );
INVX1 INVX1_84 ( .A(bundle_i[56]), .Y(_2511_) );
NAND2X1 NAND2X1_377 ( .A(_3645__24_), .B(_1039__bF_buf53), .Y(_2512_) );
OAI21X1 OAI21X1_883 ( .A(_2511_), .B(_1039__bF_buf53), .C(_2512_), .Y(_653_) );
INVX1 INVX1_85 ( .A(bundle_i[55]), .Y(_2513_) );
NAND2X1 NAND2X1_378 ( .A(_3645__23_), .B(_1039__bF_buf29), .Y(_2514_) );
OAI21X1 OAI21X1_884 ( .A(_2513_), .B(_1039__bF_buf29), .C(_2514_), .Y(_654_) );
INVX1 INVX1_86 ( .A(bundle_i[54]), .Y(_2515_) );
NAND2X1 NAND2X1_379 ( .A(_3645__22_), .B(_1039__bF_buf5), .Y(_2516_) );
OAI21X1 OAI21X1_885 ( .A(_2515_), .B(_1039__bF_buf5), .C(_2516_), .Y(_655_) );
INVX1 INVX1_87 ( .A(bundle_i[53]), .Y(_2517_) );
NAND2X1 NAND2X1_380 ( .A(_3645__21_), .B(_1039__bF_buf51), .Y(_2518_) );
OAI21X1 OAI21X1_886 ( .A(_2517_), .B(_1039__bF_buf51), .C(_2518_), .Y(_656_) );
INVX1 INVX1_88 ( .A(bundle_i[52]), .Y(_2519_) );
NAND2X1 NAND2X1_381 ( .A(_3645__20_), .B(_1039__bF_buf5), .Y(_2520_) );
OAI21X1 OAI21X1_887 ( .A(_2519_), .B(_1039__bF_buf5), .C(_2520_), .Y(_657_) );
INVX1 INVX1_89 ( .A(bundle_i[51]), .Y(_2521_) );
NAND2X1 NAND2X1_382 ( .A(_3645__19_), .B(_1039__bF_buf44), .Y(_2522_) );
OAI21X1 OAI21X1_888 ( .A(_2521_), .B(_1039__bF_buf44), .C(_2522_), .Y(_658_) );
INVX1 INVX1_90 ( .A(bundle_i[50]), .Y(_2523_) );
NAND2X1 NAND2X1_383 ( .A(_3645__18_), .B(_1039__bF_buf32), .Y(_2524_) );
OAI21X1 OAI21X1_889 ( .A(_2523_), .B(_1039__bF_buf32), .C(_2524_), .Y(_659_) );
INVX1 INVX1_91 ( .A(bundle_i[49]), .Y(_2525_) );
NAND2X1 NAND2X1_384 ( .A(_3645__17_), .B(_1039__bF_buf40), .Y(_2526_) );
OAI21X1 OAI21X1_890 ( .A(_2525_), .B(_1039__bF_buf29), .C(_2526_), .Y(_660_) );
INVX1 INVX1_92 ( .A(bundle_i[48]), .Y(_2527_) );
NAND2X1 NAND2X1_385 ( .A(_3645__16_), .B(_1039__bF_buf31), .Y(_2528_) );
OAI21X1 OAI21X1_891 ( .A(_2527_), .B(_1039__bF_buf31), .C(_2528_), .Y(_661_) );
INVX1 INVX1_93 ( .A(bundle_i[47]), .Y(_2529_) );
NAND2X1 NAND2X1_386 ( .A(_3645__15_), .B(_1039__bF_buf53), .Y(_2530_) );
OAI21X1 OAI21X1_892 ( .A(_2529_), .B(_1039__bF_buf53), .C(_2530_), .Y(_662_) );
INVX1 INVX1_94 ( .A(bundle_i[46]), .Y(_2531_) );
NAND2X1 NAND2X1_387 ( .A(_3645__14_), .B(_1039__bF_buf38), .Y(_2532_) );
OAI21X1 OAI21X1_893 ( .A(_2531_), .B(_1039__bF_buf38), .C(_2532_), .Y(_663_) );
INVX1 INVX1_95 ( .A(bundle_i[45]), .Y(_2533_) );
NAND2X1 NAND2X1_388 ( .A(_3645__13_), .B(_1039__bF_buf31), .Y(_2534_) );
OAI21X1 OAI21X1_894 ( .A(_2533_), .B(_1039__bF_buf31), .C(_2534_), .Y(_664_) );
INVX1 INVX1_96 ( .A(bundle_i[44]), .Y(_2535_) );
NAND2X1 NAND2X1_389 ( .A(_3645__12_), .B(_1039__bF_buf9), .Y(_2536_) );
OAI21X1 OAI21X1_895 ( .A(_2535_), .B(_1039__bF_buf9), .C(_2536_), .Y(_665_) );
INVX1 INVX1_97 ( .A(bundle_i[43]), .Y(_2537_) );
NAND2X1 NAND2X1_390 ( .A(_3645__11_), .B(_1039__bF_buf53), .Y(_2538_) );
OAI21X1 OAI21X1_896 ( .A(_2537_), .B(_1039__bF_buf53), .C(_2538_), .Y(_666_) );
INVX1 INVX1_98 ( .A(bundle_i[42]), .Y(_2539_) );
NAND2X1 NAND2X1_391 ( .A(_3645__10_), .B(_1039__bF_buf48), .Y(_2540_) );
OAI21X1 OAI21X1_897 ( .A(_2539_), .B(_1039__bF_buf48), .C(_2540_), .Y(_667_) );
INVX1 INVX1_99 ( .A(bundle_i[41]), .Y(_2541_) );
NAND2X1 NAND2X1_392 ( .A(_3645__9_), .B(_1039__bF_buf17), .Y(_2542_) );
OAI21X1 OAI21X1_898 ( .A(_2541_), .B(_1039__bF_buf17), .C(_2542_), .Y(_668_) );
INVX1 INVX1_100 ( .A(bundle_i[40]), .Y(_2543_) );
NAND2X1 NAND2X1_393 ( .A(_3645__8_), .B(_1039__bF_buf0), .Y(_2544_) );
OAI21X1 OAI21X1_899 ( .A(_2543_), .B(_1039__bF_buf5), .C(_2544_), .Y(_669_) );
INVX1 INVX1_101 ( .A(bundle_i[39]), .Y(_2545_) );
NAND2X1 NAND2X1_394 ( .A(_3645__7_), .B(_1039__bF_buf40), .Y(_2546_) );
OAI21X1 OAI21X1_900 ( .A(_2545_), .B(_1039__bF_buf40), .C(_2546_), .Y(_670_) );
INVX1 INVX1_102 ( .A(bundle_i[38]), .Y(_2547_) );
NAND2X1 NAND2X1_395 ( .A(_3645__6_), .B(_1039__bF_buf41), .Y(_2548_) );
OAI21X1 OAI21X1_901 ( .A(_2547_), .B(_1039__bF_buf41), .C(_2548_), .Y(_671_) );
INVX1 INVX1_103 ( .A(bundle_i[37]), .Y(_2549_) );
NAND2X1 NAND2X1_396 ( .A(_3645__5_), .B(_1039__bF_buf5), .Y(_2550_) );
OAI21X1 OAI21X1_902 ( .A(_2549_), .B(_1039__bF_buf5), .C(_2550_), .Y(_672_) );
INVX1 INVX1_104 ( .A(bundle_i[36]), .Y(_2551_) );
NAND2X1 NAND2X1_397 ( .A(_3645__4_), .B(_1039__bF_buf56), .Y(_2552_) );
OAI21X1 OAI21X1_903 ( .A(_2551_), .B(_1039__bF_buf56), .C(_2552_), .Y(_673_) );
INVX1 INVX1_105 ( .A(bundle_i[35]), .Y(_2553_) );
NAND2X1 NAND2X1_398 ( .A(_3645__3_), .B(_1039__bF_buf48), .Y(_2554_) );
OAI21X1 OAI21X1_904 ( .A(_2553_), .B(_1039__bF_buf48), .C(_2554_), .Y(_674_) );
INVX1 INVX1_106 ( .A(bundle_i[34]), .Y(_2555_) );
NAND2X1 NAND2X1_399 ( .A(_3645__2_), .B(_1039__bF_buf48), .Y(_2556_) );
OAI21X1 OAI21X1_905 ( .A(_2555_), .B(_1039__bF_buf48), .C(_2556_), .Y(_675_) );
INVX1 INVX1_107 ( .A(bundle_i[33]), .Y(_2557_) );
NAND2X1 NAND2X1_400 ( .A(_3645__1_), .B(_1039__bF_buf9), .Y(_2558_) );
OAI21X1 OAI21X1_906 ( .A(_2557_), .B(_1039__bF_buf9), .C(_2558_), .Y(_676_) );
INVX1 INVX1_108 ( .A(bundle_i[32]), .Y(_2559_) );
NAND2X1 NAND2X1_401 ( .A(_3645__0_), .B(_1039__bF_buf53), .Y(_2560_) );
OAI21X1 OAI21X1_907 ( .A(_2559_), .B(_1039__bF_buf53), .C(_2560_), .Y(_677_) );
INVX1 INVX1_109 ( .A(bundle_i[95]), .Y(_2561_) );
OAI21X1 OAI21X1_908 ( .A(_1100__bF_buf14_bF_buf0), .B(_1031__bF_buf6), .C(_3646__31_), .Y(_2562_) );
OAI21X1 OAI21X1_909 ( .A(_1101__bF_buf53), .B(_2561_), .C(_2562_), .Y(_678_) );
INVX1 INVX1_110 ( .A(bundle_i[94]), .Y(_2563_) );
OAI21X1 OAI21X1_910 ( .A(_1100__bF_buf13_bF_buf3), .B(_1031__bF_buf13), .C(_3646__30_), .Y(_2564_) );
OAI21X1 OAI21X1_911 ( .A(_1101__bF_buf39), .B(_2563_), .C(_2564_), .Y(_679_) );
INVX1 INVX1_111 ( .A(bundle_i[93]), .Y(_2565_) );
OAI21X1 OAI21X1_912 ( .A(_1100__bF_buf12_bF_buf2), .B(_1031__bF_buf73), .C(_3646__29_), .Y(_2566_) );
OAI21X1 OAI21X1_913 ( .A(_1101__bF_buf26), .B(_2565_), .C(_2566_), .Y(_680_) );
INVX1 INVX1_112 ( .A(bundle_i[92]), .Y(_2567_) );
OAI21X1 OAI21X1_914 ( .A(_1100__bF_buf11_bF_buf0), .B(_1031__bF_buf59), .C(_3646__28_), .Y(_2568_) );
OAI21X1 OAI21X1_915 ( .A(_1101__bF_buf36), .B(_2567_), .C(_2568_), .Y(_681_) );
INVX1 INVX1_113 ( .A(bundle_i[91]), .Y(_2569_) );
OAI21X1 OAI21X1_916 ( .A(_1100__bF_buf10_bF_buf0), .B(_1031__bF_buf50), .C(_3646__27_), .Y(_2570_) );
OAI21X1 OAI21X1_917 ( .A(_1101__bF_buf25), .B(_2569_), .C(_2570_), .Y(_682_) );
INVX1 INVX1_114 ( .A(bundle_i[90]), .Y(_2571_) );
OAI21X1 OAI21X1_918 ( .A(_1100__bF_buf9_bF_buf0), .B(_1031__bF_buf14), .C(_3646__26_), .Y(_2572_) );
OAI21X1 OAI21X1_919 ( .A(_1101__bF_buf40), .B(_2571_), .C(_2572_), .Y(_683_) );
INVX1 INVX1_115 ( .A(bundle_i[89]), .Y(_2573_) );
OAI21X1 OAI21X1_920 ( .A(_1100__bF_buf8_bF_buf2), .B(_1031__bF_buf50), .C(_3646__25_), .Y(_2574_) );
OAI21X1 OAI21X1_921 ( .A(_1101__bF_buf25), .B(_2573_), .C(_2574_), .Y(_684_) );
INVX1 INVX1_116 ( .A(bundle_i[88]), .Y(_2575_) );
OAI21X1 OAI21X1_922 ( .A(_1100__bF_buf7_bF_buf3), .B(_1031__bF_buf58), .C(_3646__24_), .Y(_2576_) );
OAI21X1 OAI21X1_923 ( .A(_1101__bF_buf38), .B(_2575_), .C(_2576_), .Y(_685_) );
INVX1 INVX1_117 ( .A(bundle_i[87]), .Y(_2577_) );
OAI21X1 OAI21X1_924 ( .A(_1100__bF_buf4), .B(_1031__bF_buf36), .C(_3646__23_), .Y(_2578_) );
OAI21X1 OAI21X1_925 ( .A(_1101__bF_buf36), .B(_2577_), .C(_2578_), .Y(_686_) );
INVX1 INVX1_118 ( .A(bundle_i[86]), .Y(_2579_) );
OAI21X1 OAI21X1_926 ( .A(_1100__bF_buf5), .B(_1031__bF_buf19), .C(_3646__22_), .Y(_2580_) );
OAI21X1 OAI21X1_927 ( .A(_1101__bF_buf55), .B(_2579_), .C(_2580_), .Y(_687_) );
INVX1 INVX1_119 ( .A(bundle_i[85]), .Y(_2581_) );
OAI21X1 OAI21X1_928 ( .A(_1100__bF_buf13), .B(_1031__bF_buf59), .C(_3646__21_), .Y(_2582_) );
OAI21X1 OAI21X1_929 ( .A(_1101__bF_buf36), .B(_2581_), .C(_2582_), .Y(_688_) );
INVX1 INVX1_120 ( .A(bundle_i[84]), .Y(_2583_) );
OAI21X1 OAI21X1_930 ( .A(_1100__bF_buf3), .B(_1031__bF_buf56), .C(_3646__20_), .Y(_2584_) );
OAI21X1 OAI21X1_931 ( .A(_1101__bF_buf56), .B(_2583_), .C(_2584_), .Y(_689_) );
INVX1 INVX1_121 ( .A(bundle_i[83]), .Y(_2585_) );
OAI21X1 OAI21X1_932 ( .A(_1100__bF_buf4), .B(_1031__bF_buf36), .C(_3646__19_), .Y(_2586_) );
OAI21X1 OAI21X1_933 ( .A(_1101__bF_buf43), .B(_2585_), .C(_2586_), .Y(_690_) );
INVX1 INVX1_122 ( .A(bundle_i[82]), .Y(_2587_) );
OAI21X1 OAI21X1_934 ( .A(_1100__bF_buf6), .B(_1031__bF_buf73), .C(_3646__18_), .Y(_2588_) );
OAI21X1 OAI21X1_935 ( .A(_1101__bF_buf26), .B(_2587_), .C(_2588_), .Y(_691_) );
INVX1 INVX1_123 ( .A(bundle_i[81]), .Y(_2589_) );
OAI21X1 OAI21X1_936 ( .A(_1100__bF_buf13), .B(_1031__bF_buf59), .C(_3646__17_), .Y(_2590_) );
OAI21X1 OAI21X1_937 ( .A(_1101__bF_buf36), .B(_2589_), .C(_2590_), .Y(_692_) );
INVX1 INVX1_124 ( .A(bundle_i[80]), .Y(_2591_) );
OAI21X1 OAI21X1_938 ( .A(_1100__bF_buf14_bF_buf1), .B(_1031__bF_buf58), .C(_3646__16_), .Y(_2592_) );
OAI21X1 OAI21X1_939 ( .A(_1101__bF_buf38), .B(_2591_), .C(_2592_), .Y(_693_) );
INVX1 INVX1_125 ( .A(bundle_i[79]), .Y(_2593_) );
OAI21X1 OAI21X1_940 ( .A(_1100__bF_buf13_bF_buf3), .B(_1031__bF_buf57), .C(_3646__15_), .Y(_2594_) );
OAI21X1 OAI21X1_941 ( .A(_1101__bF_buf35), .B(_2593_), .C(_2594_), .Y(_694_) );
INVX1 INVX1_126 ( .A(bundle_i[78]), .Y(_2595_) );
OAI21X1 OAI21X1_942 ( .A(_1100__bF_buf12_bF_buf0), .B(_1031__bF_buf62), .C(_3646__14_), .Y(_2596_) );
OAI21X1 OAI21X1_943 ( .A(_1101__bF_buf55), .B(_2595_), .C(_2596_), .Y(_695_) );
INVX1 INVX1_127 ( .A(bundle_i[77]), .Y(_2597_) );
OAI21X1 OAI21X1_944 ( .A(_1100__bF_buf11_bF_buf0), .B(_1031__bF_buf36), .C(_3646__13_), .Y(_2598_) );
OAI21X1 OAI21X1_945 ( .A(_1101__bF_buf36), .B(_2597_), .C(_2598_), .Y(_696_) );
INVX1 INVX1_128 ( .A(bundle_i[76]), .Y(_2599_) );
OAI21X1 OAI21X1_946 ( .A(_1100__bF_buf10_bF_buf0), .B(_1031__bF_buf50), .C(_3646__12_), .Y(_2600_) );
OAI21X1 OAI21X1_947 ( .A(_1101__bF_buf25), .B(_2599_), .C(_2600_), .Y(_697_) );
INVX1 INVX1_129 ( .A(bundle_i[75]), .Y(_2601_) );
OAI21X1 OAI21X1_948 ( .A(_1100__bF_buf9_bF_buf1), .B(_1031__bF_buf47), .C(_3646__11_), .Y(_2602_) );
OAI21X1 OAI21X1_949 ( .A(_1101__bF_buf14), .B(_2601_), .C(_2602_), .Y(_698_) );
INVX1 INVX1_130 ( .A(bundle_i[74]), .Y(_2603_) );
OAI21X1 OAI21X1_950 ( .A(_1100__bF_buf8_bF_buf0), .B(_1031__bF_buf20), .C(_3646__10_), .Y(_2604_) );
OAI21X1 OAI21X1_951 ( .A(_1101__bF_buf43), .B(_2603_), .C(_2604_), .Y(_699_) );
INVX1 INVX1_131 ( .A(bundle_i[73]), .Y(_2605_) );
OAI21X1 OAI21X1_952 ( .A(_1100__bF_buf7_bF_buf3), .B(_1031__bF_buf58), .C(_3646__9_), .Y(_2606_) );
OAI21X1 OAI21X1_953 ( .A(_1101__bF_buf38), .B(_2605_), .C(_2606_), .Y(_700_) );
INVX1 INVX1_132 ( .A(bundle_i[72]), .Y(_2607_) );
OAI21X1 OAI21X1_954 ( .A(_1100__bF_buf5), .B(_1031__bF_buf62), .C(_3646__8_), .Y(_2608_) );
OAI21X1 OAI21X1_955 ( .A(_1101__bF_buf55), .B(_2607_), .C(_2608_), .Y(_701_) );
INVX1 INVX1_133 ( .A(bundle_i[71]), .Y(_2609_) );
OAI21X1 OAI21X1_956 ( .A(_1100__bF_buf13), .B(_1031__bF_buf59), .C(_3646__7_), .Y(_2610_) );
OAI21X1 OAI21X1_957 ( .A(_1101__bF_buf36), .B(_2609_), .C(_2610_), .Y(_702_) );
INVX1 INVX1_134 ( .A(bundle_i[70]), .Y(_2611_) );
OAI21X1 OAI21X1_958 ( .A(_1100__bF_buf2), .B(_1031__bF_buf50), .C(_3646__6_), .Y(_2612_) );
OAI21X1 OAI21X1_959 ( .A(_1101__bF_buf25), .B(_2611_), .C(_2612_), .Y(_703_) );
INVX1 INVX1_135 ( .A(bundle_i[69]), .Y(_2613_) );
OAI21X1 OAI21X1_960 ( .A(_1100__bF_buf6), .B(_1031__bF_buf73), .C(_3646__5_), .Y(_2614_) );
OAI21X1 OAI21X1_961 ( .A(_1101__bF_buf26), .B(_2613_), .C(_2614_), .Y(_704_) );
INVX1 INVX1_136 ( .A(bundle_i[68]), .Y(_2615_) );
OAI21X1 OAI21X1_962 ( .A(_1100__bF_buf6), .B(_1031__bF_buf73), .C(_3646__4_), .Y(_2616_) );
OAI21X1 OAI21X1_963 ( .A(_1101__bF_buf26), .B(_2615_), .C(_2616_), .Y(_705_) );
INVX1 INVX1_137 ( .A(bundle_i[67]), .Y(_2617_) );
OAI21X1 OAI21X1_964 ( .A(_1100__bF_buf0), .B(_1031__bF_buf53), .C(_3646__3_), .Y(_2618_) );
OAI21X1 OAI21X1_965 ( .A(_1101__bF_buf48), .B(_2617_), .C(_2618_), .Y(_706_) );
INVX1 INVX1_138 ( .A(bundle_i[66]), .Y(_2619_) );
OAI21X1 OAI21X1_966 ( .A(_1100__bF_buf6), .B(_1031__bF_buf73), .C(_3646__2_), .Y(_2620_) );
OAI21X1 OAI21X1_967 ( .A(_1101__bF_buf26), .B(_2619_), .C(_2620_), .Y(_707_) );
INVX1 INVX1_139 ( .A(bundle_i[65]), .Y(_2621_) );
OAI21X1 OAI21X1_968 ( .A(_1100__bF_buf14_bF_buf1), .B(_1031__bF_buf56), .C(_3646__1_), .Y(_2622_) );
OAI21X1 OAI21X1_969 ( .A(_1101__bF_buf56), .B(_2621_), .C(_2622_), .Y(_708_) );
INVX1 INVX1_140 ( .A(bundle_i[64]), .Y(_2623_) );
OAI21X1 OAI21X1_970 ( .A(_1100__bF_buf13_bF_buf2), .B(_1031__bF_buf70), .C(_3646__0_), .Y(_2624_) );
OAI21X1 OAI21X1_971 ( .A(_1101__bF_buf1), .B(_2623_), .C(_2624_), .Y(_709_) );
INVX1 INVX1_141 ( .A(bundle_i[127]), .Y(_2625_) );
OAI21X1 OAI21X1_972 ( .A(_1101__bF_buf46), .B(_1135__bF_buf8_bF_buf2), .C(_3647__31_), .Y(_2626_) );
OAI21X1 OAI21X1_973 ( .A(_1134__bF_buf8), .B(_2625_), .C(_2626_), .Y(_710_) );
INVX1 INVX1_142 ( .A(bundle_i[126]), .Y(_2627_) );
OAI21X1 OAI21X1_974 ( .A(_1101__bF_buf42), .B(_1135__bF_buf7_bF_buf1), .C(_3647__30_), .Y(_2628_) );
OAI21X1 OAI21X1_975 ( .A(_1134__bF_buf10), .B(_2627_), .C(_2628_), .Y(_711_) );
INVX1 INVX1_143 ( .A(bundle_i[125]), .Y(_2629_) );
OAI21X1 OAI21X1_976 ( .A(_1101__bF_buf17), .B(_1135__bF_buf6_bF_buf3), .C(_3647__29_), .Y(_2630_) );
OAI21X1 OAI21X1_977 ( .A(_1134__bF_buf6), .B(_2629_), .C(_2630_), .Y(_712_) );
INVX1 INVX1_144 ( .A(bundle_i[124]), .Y(_2631_) );
OAI21X1 OAI21X1_978 ( .A(_1101__bF_buf15), .B(_1135__bF_buf5_bF_buf2), .C(_3647__28_), .Y(_2632_) );
OAI21X1 OAI21X1_979 ( .A(_1134__bF_buf12), .B(_2631_), .C(_2632_), .Y(_713_) );
INVX1 INVX1_145 ( .A(bundle_i[123]), .Y(_2633_) );
OAI21X1 OAI21X1_980 ( .A(_1101__bF_buf39), .B(_1135__bF_buf4_bF_buf3), .C(_3647__27_), .Y(_2634_) );
OAI21X1 OAI21X1_981 ( .A(_1134__bF_buf10), .B(_2633_), .C(_2634_), .Y(_714_) );
INVX1 INVX1_146 ( .A(bundle_i[122]), .Y(_2635_) );
OAI21X1 OAI21X1_982 ( .A(_1101__bF_buf27), .B(_1135__bF_buf3_bF_buf3), .C(_3647__26_), .Y(_2636_) );
OAI21X1 OAI21X1_983 ( .A(_1134__bF_buf9), .B(_2635_), .C(_2636_), .Y(_715_) );
INVX1 INVX1_147 ( .A(bundle_i[121]), .Y(_2637_) );
OAI21X1 OAI21X1_984 ( .A(_1101__bF_buf42), .B(_1135__bF_buf2_bF_buf0), .C(_3647__25_), .Y(_2638_) );
OAI21X1 OAI21X1_985 ( .A(_1134__bF_buf10), .B(_2637_), .C(_2638_), .Y(_716_) );
INVX1 INVX1_148 ( .A(bundle_i[120]), .Y(_2639_) );
OAI21X1 OAI21X1_986 ( .A(_1101__bF_buf21), .B(_1135__bF_buf1_bF_buf2), .C(_3647__24_), .Y(_2640_) );
OAI21X1 OAI21X1_987 ( .A(_1134__bF_buf0), .B(_2639_), .C(_2640_), .Y(_717_) );
INVX1 INVX1_149 ( .A(bundle_i[119]), .Y(_2641_) );
OAI21X1 OAI21X1_988 ( .A(_1101__bF_buf49), .B(_1135__bF_buf0), .C(_3647__23_), .Y(_2642_) );
OAI21X1 OAI21X1_989 ( .A(_1134__bF_buf8), .B(_2641_), .C(_2642_), .Y(_718_) );
INVX1 INVX1_150 ( .A(bundle_i[118]), .Y(_2643_) );
OAI21X1 OAI21X1_990 ( .A(_1101__bF_buf43), .B(_1135__bF_buf14_bF_buf1), .C(_3647__22_), .Y(_2644_) );
OAI21X1 OAI21X1_991 ( .A(_1134__bF_buf7), .B(_2643_), .C(_2644_), .Y(_719_) );
INVX1 INVX1_151 ( .A(bundle_i[117]), .Y(_2645_) );
OAI21X1 OAI21X1_992 ( .A(_1101__bF_buf43), .B(_1135__bF_buf13_bF_buf3), .C(_3647__21_), .Y(_2646_) );
OAI21X1 OAI21X1_993 ( .A(_1134__bF_buf7), .B(_2645_), .C(_2646_), .Y(_720_) );
INVX1 INVX1_152 ( .A(bundle_i[116]), .Y(_2647_) );
OAI21X1 OAI21X1_994 ( .A(_1101__bF_buf2), .B(_1135__bF_buf12_bF_buf0), .C(_3647__20_), .Y(_2648_) );
OAI21X1 OAI21X1_995 ( .A(_1134__bF_buf3), .B(_2647_), .C(_2648_), .Y(_721_) );
INVX1 INVX1_153 ( .A(bundle_i[115]), .Y(_2649_) );
OAI21X1 OAI21X1_996 ( .A(_1101__bF_buf40), .B(_1135__bF_buf11_bF_buf2), .C(_3647__19_), .Y(_2650_) );
OAI21X1 OAI21X1_997 ( .A(_1134__bF_buf0), .B(_2649_), .C(_2650_), .Y(_722_) );
INVX1 INVX1_154 ( .A(bundle_i[114]), .Y(_2651_) );
OAI21X1 OAI21X1_998 ( .A(_1101__bF_buf30), .B(_1135__bF_buf10_bF_buf1), .C(_3647__18_), .Y(_2652_) );
OAI21X1 OAI21X1_999 ( .A(_1134__bF_buf12), .B(_2651_), .C(_2652_), .Y(_723_) );
INVX1 INVX1_155 ( .A(bundle_i[113]), .Y(_2653_) );
OAI21X1 OAI21X1_1000 ( .A(_1101__bF_buf21), .B(_1135__bF_buf9_bF_buf3), .C(_3647__17_), .Y(_2654_) );
OAI21X1 OAI21X1_1001 ( .A(_1134__bF_buf0), .B(_2653_), .C(_2654_), .Y(_724_) );
INVX1 INVX1_156 ( .A(bundle_i[112]), .Y(_2655_) );
OAI21X1 OAI21X1_1002 ( .A(_1101__bF_buf35), .B(_1135__bF_buf8_bF_buf0), .C(_3647__16_), .Y(_2656_) );
OAI21X1 OAI21X1_1003 ( .A(_1134__bF_buf0), .B(_2655_), .C(_2656_), .Y(_725_) );
INVX1 INVX1_157 ( .A(bundle_i[111]), .Y(_2657_) );
OAI21X1 OAI21X1_1004 ( .A(_1101__bF_buf25), .B(_1135__bF_buf7_bF_buf3), .C(_3647__15_), .Y(_2658_) );
OAI21X1 OAI21X1_1005 ( .A(_1134__bF_buf0), .B(_2657_), .C(_2658_), .Y(_726_) );
INVX1 INVX1_158 ( .A(bundle_i[110]), .Y(_2659_) );
OAI21X1 OAI21X1_1006 ( .A(_1101__bF_buf28), .B(_1135__bF_buf6_bF_buf1), .C(_3647__14_), .Y(_2660_) );
OAI21X1 OAI21X1_1007 ( .A(_1134__bF_buf7), .B(_2659_), .C(_2660_), .Y(_727_) );
INVX1 INVX1_159 ( .A(bundle_i[109]), .Y(_2661_) );
OAI21X1 OAI21X1_1008 ( .A(_1101__bF_buf6), .B(_1135__bF_buf5_bF_buf0), .C(_3647__13_), .Y(_2662_) );
OAI21X1 OAI21X1_1009 ( .A(_1134__bF_buf1), .B(_2661_), .C(_2662_), .Y(_728_) );
INVX1 INVX1_160 ( .A(bundle_i[108]), .Y(_2663_) );
OAI21X1 OAI21X1_1010 ( .A(_1101__bF_buf21), .B(_1135__bF_buf4_bF_buf3), .C(_3647__12_), .Y(_2664_) );
OAI21X1 OAI21X1_1011 ( .A(_1134__bF_buf0), .B(_2663_), .C(_2664_), .Y(_729_) );
INVX1 INVX1_161 ( .A(bundle_i[107]), .Y(_2665_) );
OAI21X1 OAI21X1_1012 ( .A(_1101__bF_buf21), .B(_1135__bF_buf3_bF_buf3), .C(_3647__11_), .Y(_2666_) );
OAI21X1 OAI21X1_1013 ( .A(_1134__bF_buf0), .B(_2665_), .C(_2666_), .Y(_730_) );
INVX1 INVX1_162 ( .A(bundle_i[106]), .Y(_2667_) );
OAI21X1 OAI21X1_1014 ( .A(_1101__bF_buf22), .B(_1135__bF_buf2_bF_buf2), .C(_3647__10_), .Y(_2668_) );
OAI21X1 OAI21X1_1015 ( .A(_1134__bF_buf9), .B(_2667_), .C(_2668_), .Y(_731_) );
INVX1 INVX1_163 ( .A(bundle_i[105]), .Y(_2669_) );
OAI21X1 OAI21X1_1016 ( .A(_1101__bF_buf46), .B(_1135__bF_buf1_bF_buf3), .C(_3647__9_), .Y(_2670_) );
OAI21X1 OAI21X1_1017 ( .A(_1134__bF_buf8), .B(_2669_), .C(_2670_), .Y(_732_) );
INVX1 INVX1_164 ( .A(bundle_i[104]), .Y(_2671_) );
OAI21X1 OAI21X1_1018 ( .A(_1101__bF_buf54), .B(_1135__bF_buf1), .C(_3647__8_), .Y(_2672_) );
OAI21X1 OAI21X1_1019 ( .A(_1134__bF_buf7), .B(_2671_), .C(_2672_), .Y(_733_) );
INVX1 INVX1_165 ( .A(bundle_i[103]), .Y(_2673_) );
OAI21X1 OAI21X1_1020 ( .A(_1101__bF_buf43), .B(_1135__bF_buf14_bF_buf1), .C(_3647__7_), .Y(_2674_) );
OAI21X1 OAI21X1_1021 ( .A(_1134__bF_buf7), .B(_2673_), .C(_2674_), .Y(_734_) );
INVX1 INVX1_166 ( .A(bundle_i[102]), .Y(_2675_) );
OAI21X1 OAI21X1_1022 ( .A(_1101__bF_buf43), .B(_1135__bF_buf13_bF_buf3), .C(_3647__6_), .Y(_2676_) );
OAI21X1 OAI21X1_1023 ( .A(_1134__bF_buf7), .B(_2675_), .C(_2676_), .Y(_735_) );
INVX1 INVX1_167 ( .A(bundle_i[101]), .Y(_2677_) );
OAI21X1 OAI21X1_1024 ( .A(_1101__bF_buf25), .B(_1135__bF_buf12_bF_buf1), .C(_3647__5_), .Y(_2678_) );
OAI21X1 OAI21X1_1025 ( .A(_1134__bF_buf0), .B(_2677_), .C(_2678_), .Y(_736_) );
INVX1 INVX1_168 ( .A(bundle_i[100]), .Y(_2679_) );
OAI21X1 OAI21X1_1026 ( .A(_1101__bF_buf26), .B(_1135__bF_buf11_bF_buf1), .C(_3647__4_), .Y(_2680_) );
OAI21X1 OAI21X1_1027 ( .A(_1134__bF_buf1), .B(_2679_), .C(_2680_), .Y(_737_) );
INVX1 INVX1_169 ( .A(bundle_i[99]), .Y(_2681_) );
OAI21X1 OAI21X1_1028 ( .A(_1101__bF_buf15), .B(_1135__bF_buf10_bF_buf2), .C(_3647__3_), .Y(_2682_) );
OAI21X1 OAI21X1_1029 ( .A(_1134__bF_buf12), .B(_2681_), .C(_2682_), .Y(_738_) );
INVX1 INVX1_170 ( .A(bundle_i[98]), .Y(_2683_) );
OAI21X1 OAI21X1_1030 ( .A(_1101__bF_buf42), .B(_1135__bF_buf9_bF_buf2), .C(_3647__2_), .Y(_2684_) );
OAI21X1 OAI21X1_1031 ( .A(_1134__bF_buf10), .B(_2683_), .C(_2684_), .Y(_739_) );
INVX1 INVX1_171 ( .A(bundle_i[97]), .Y(_2685_) );
OAI21X1 OAI21X1_1032 ( .A(_1101__bF_buf7), .B(_1135__bF_buf8_bF_buf3), .C(_3647__1_), .Y(_2686_) );
OAI21X1 OAI21X1_1033 ( .A(_1134__bF_buf2), .B(_2685_), .C(_2686_), .Y(_740_) );
INVX1 INVX1_172 ( .A(bundle_i[96]), .Y(_2687_) );
OAI21X1 OAI21X1_1034 ( .A(_1101__bF_buf25), .B(_1135__bF_buf7_bF_buf3), .C(_3647__0_), .Y(_2688_) );
OAI21X1 OAI21X1_1035 ( .A(_1134__bF_buf0), .B(_2687_), .C(_2688_), .Y(_741_) );
INVX2 INVX2_54 ( .A(bundleAddress_i[63]), .Y(_2689_) );
NAND2X1 NAND2X1_402 ( .A(_3636__63_), .B(_1031__bF_buf66), .Y(_2690_) );
OAI21X1 OAI21X1_1036 ( .A(_1031__bF_buf66), .B(_2689_), .C(_2690_), .Y(_742_) );
INVX2 INVX2_55 ( .A(bundleAddress_i[62]), .Y(_2691_) );
NAND2X1 NAND2X1_403 ( .A(_3636__62_), .B(_1031__bF_buf12), .Y(_2692_) );
OAI21X1 OAI21X1_1037 ( .A(_1031__bF_buf12), .B(_2691_), .C(_2692_), .Y(_743_) );
INVX4 INVX4_32 ( .A(bundleAddress_i[61]), .Y(_2693_) );
NAND2X1 NAND2X1_404 ( .A(_3636__61_), .B(_1031__bF_buf35), .Y(_2694_) );
OAI21X1 OAI21X1_1038 ( .A(_2693_), .B(_1031__bF_buf35), .C(_2694_), .Y(_744_) );
INVX2 INVX2_56 ( .A(bundleAddress_i[60]), .Y(_2695_) );
NAND2X1 NAND2X1_405 ( .A(_3636__60_), .B(_1031__bF_buf76), .Y(_2696_) );
OAI21X1 OAI21X1_1039 ( .A(_1031__bF_buf76), .B(_2695_), .C(_2696_), .Y(_745_) );
INVX2 INVX2_57 ( .A(bundleAddress_i[59]), .Y(_2697_) );
NAND2X1 NAND2X1_406 ( .A(_3636__59_), .B(_1031__bF_buf41), .Y(_2698_) );
OAI21X1 OAI21X1_1040 ( .A(_1031__bF_buf41), .B(_2697_), .C(_2698_), .Y(_746_) );
INVX2 INVX2_58 ( .A(bundleAddress_i[58]), .Y(_2699_) );
NAND2X1 NAND2X1_407 ( .A(_3636__58_), .B(_1031__bF_buf41), .Y(_2700_) );
OAI21X1 OAI21X1_1041 ( .A(_1031__bF_buf41), .B(_2699_), .C(_2700_), .Y(_747_) );
INVX2 INVX2_59 ( .A(bundleAddress_i[57]), .Y(_2701_) );
NAND2X1 NAND2X1_408 ( .A(_3636__57_), .B(_1031__bF_buf41), .Y(_2702_) );
OAI21X1 OAI21X1_1042 ( .A(_1031__bF_buf41), .B(_2701_), .C(_2702_), .Y(_748_) );
INVX2 INVX2_60 ( .A(bundleAddress_i[56]), .Y(_2703_) );
NAND2X1 NAND2X1_409 ( .A(_3636__56_), .B(_1031__bF_buf35), .Y(_2704_) );
OAI21X1 OAI21X1_1043 ( .A(_1031__bF_buf35), .B(_2703_), .C(_2704_), .Y(_749_) );
INVX2 INVX2_61 ( .A(bundleAddress_i[55]), .Y(_2705_) );
NAND2X1 NAND2X1_410 ( .A(_3636__55_), .B(_1031__bF_buf6), .Y(_2706_) );
OAI21X1 OAI21X1_1044 ( .A(_1031__bF_buf35), .B(_2705_), .C(_2706_), .Y(_750_) );
INVX2 INVX2_62 ( .A(bundleAddress_i[54]), .Y(_2707_) );
NAND2X1 NAND2X1_411 ( .A(_3636__54_), .B(_1031__bF_buf6), .Y(_2708_) );
OAI21X1 OAI21X1_1045 ( .A(_1031__bF_buf6), .B(_2707_), .C(_2708_), .Y(_751_) );
INVX2 INVX2_63 ( .A(bundleAddress_i[53]), .Y(_2709_) );
NAND2X1 NAND2X1_412 ( .A(_3636__53_), .B(_1031__bF_buf60), .Y(_2710_) );
OAI21X1 OAI21X1_1046 ( .A(_1031__bF_buf60), .B(_2709_), .C(_2710_), .Y(_752_) );
INVX4 INVX4_33 ( .A(bundleAddress_i[52]), .Y(_2711_) );
NAND2X1 NAND2X1_413 ( .A(_3636__52_), .B(_1031__bF_buf2), .Y(_2712_) );
OAI21X1 OAI21X1_1047 ( .A(_1031__bF_buf2), .B(_2711_), .C(_2712_), .Y(_753_) );
INVX2 INVX2_64 ( .A(bundleAddress_i[51]), .Y(_2713_) );
NAND2X1 NAND2X1_414 ( .A(_3636__51_), .B(_1031__bF_buf2), .Y(_2714_) );
OAI21X1 OAI21X1_1048 ( .A(_1031__bF_buf2), .B(_2713_), .C(_2714_), .Y(_754_) );
INVX2 INVX2_65 ( .A(bundleAddress_i[50]), .Y(_2715_) );
NAND2X1 NAND2X1_415 ( .A(_3636__50_), .B(_1031__bF_buf48), .Y(_2716_) );
OAI21X1 OAI21X1_1049 ( .A(_1031__bF_buf48), .B(_2715_), .C(_2716_), .Y(_755_) );
INVX2 INVX2_66 ( .A(bundleAddress_i[49]), .Y(_2717_) );
NAND2X1 NAND2X1_416 ( .A(_3636__49_), .B(_1031__bF_buf48), .Y(_2718_) );
OAI21X1 OAI21X1_1050 ( .A(_1031__bF_buf48), .B(_2717_), .C(_2718_), .Y(_756_) );
INVX2 INVX2_67 ( .A(bundleAddress_i[48]), .Y(_2719_) );
NAND2X1 NAND2X1_417 ( .A(_3636__48_), .B(_1031__bF_buf3), .Y(_2720_) );
OAI21X1 OAI21X1_1051 ( .A(_1031__bF_buf3), .B(_2719_), .C(_2720_), .Y(_757_) );
INVX4 INVX4_34 ( .A(bundleAddress_i[47]), .Y(_2721_) );
NAND2X1 NAND2X1_418 ( .A(_3636__47_), .B(_1031__bF_buf32), .Y(_2722_) );
OAI21X1 OAI21X1_1052 ( .A(_1031__bF_buf32), .B(_2721_), .C(_2722_), .Y(_758_) );
INVX2 INVX2_68 ( .A(bundleAddress_i[46]), .Y(_2723_) );
NAND2X1 NAND2X1_419 ( .A(_3636__46_), .B(_1031__bF_buf29), .Y(_2724_) );
OAI21X1 OAI21X1_1053 ( .A(_1031__bF_buf3), .B(_2723_), .C(_2724_), .Y(_759_) );
INVX2 INVX2_69 ( .A(bundleAddress_i[45]), .Y(_2725_) );
NAND2X1 NAND2X1_420 ( .A(_3636__45_), .B(_1031__bF_buf77), .Y(_2726_) );
OAI21X1 OAI21X1_1054 ( .A(_1031__bF_buf77), .B(_2725_), .C(_2726_), .Y(_760_) );
INVX4 INVX4_35 ( .A(bundleAddress_i[44]), .Y(_2727_) );
NAND2X1 NAND2X1_421 ( .A(_3636__44_), .B(_1031__bF_buf17), .Y(_2728_) );
OAI21X1 OAI21X1_1055 ( .A(_1031__bF_buf17), .B(_2727_), .C(_2728_), .Y(_761_) );
INVX1 INVX1_173 ( .A(bundleAddress_i[43]), .Y(_2729_) );
NAND2X1 NAND2X1_422 ( .A(_3636__43_), .B(_1031__bF_buf34), .Y(_2730_) );
OAI21X1 OAI21X1_1056 ( .A(_1031__bF_buf34), .B(_2729_), .C(_2730_), .Y(_762_) );
INVX4 INVX4_36 ( .A(bundleAddress_i[42]), .Y(_2731_) );
NAND2X1 NAND2X1_423 ( .A(_3636__42_), .B(_1031__bF_buf34), .Y(_2732_) );
OAI21X1 OAI21X1_1057 ( .A(_1031__bF_buf34), .B(_2731_), .C(_2732_), .Y(_763_) );
INVX2 INVX2_70 ( .A(bundleAddress_i[41]), .Y(_2733_) );
NAND2X1 NAND2X1_424 ( .A(_3636__41_), .B(_1031__bF_buf19), .Y(_2734_) );
OAI21X1 OAI21X1_1058 ( .A(_1031__bF_buf19), .B(_2733_), .C(_2734_), .Y(_764_) );
INVX1 INVX1_174 ( .A(bundleAddress_i[40]), .Y(_2735_) );
NAND2X1 NAND2X1_425 ( .A(_3636__40_), .B(_1031__bF_buf62), .Y(_2736_) );
OAI21X1 OAI21X1_1059 ( .A(_1031__bF_buf62), .B(_2735_), .C(_2736_), .Y(_765_) );
INVX1 INVX1_175 ( .A(bundleAddress_i[39]), .Y(_2737_) );
NAND2X1 NAND2X1_426 ( .A(_3636__39_), .B(_1031__bF_buf34), .Y(_2738_) );
OAI21X1 OAI21X1_1060 ( .A(_1031__bF_buf34), .B(_2737_), .C(_2738_), .Y(_766_) );
INVX4 INVX4_37 ( .A(bundleAddress_i[38]), .Y(_2739_) );
NAND2X1 NAND2X1_427 ( .A(_3636__38_), .B(_1031__bF_buf17), .Y(_2740_) );
OAI21X1 OAI21X1_1061 ( .A(_1031__bF_buf17), .B(_2739_), .C(_2740_), .Y(_767_) );
INVX2 INVX2_71 ( .A(bundleAddress_i[37]), .Y(_2741_) );
NAND2X1 NAND2X1_428 ( .A(_3636__37_), .B(_1031__bF_buf71), .Y(_2742_) );
OAI21X1 OAI21X1_1062 ( .A(_1031__bF_buf71), .B(_2741_), .C(_2742_), .Y(_768_) );
INVX2 INVX2_72 ( .A(bundleAddress_i[36]), .Y(_2743_) );
NAND2X1 NAND2X1_429 ( .A(_3636__36_), .B(_1031__bF_buf71), .Y(_2744_) );
OAI21X1 OAI21X1_1063 ( .A(_1031__bF_buf71), .B(_2743_), .C(_2744_), .Y(_769_) );
INVX1 INVX1_176 ( .A(bundleAddress_i[35]), .Y(_2745_) );
NAND2X1 NAND2X1_430 ( .A(_3636__35_), .B(_1031__bF_buf77), .Y(_2746_) );
OAI21X1 OAI21X1_1064 ( .A(_1031__bF_buf71), .B(_2745_), .C(_2746_), .Y(_770_) );
INVX4 INVX4_38 ( .A(bundleAddress_i[34]), .Y(_2747_) );
NAND2X1 NAND2X1_431 ( .A(_3636__34_), .B(_1031__bF_buf11), .Y(_2748_) );
OAI21X1 OAI21X1_1065 ( .A(_1031__bF_buf11), .B(_2747_), .C(_2748_), .Y(_771_) );
INVX2 INVX2_73 ( .A(bundleAddress_i[33]), .Y(_2749_) );
NAND2X1 NAND2X1_432 ( .A(_3636__33_), .B(_1031__bF_buf11), .Y(_2750_) );
OAI21X1 OAI21X1_1066 ( .A(_1031__bF_buf11), .B(_2749_), .C(_2750_), .Y(_772_) );
INVX4 INVX4_39 ( .A(bundleAddress_i[32]), .Y(_2751_) );
NAND2X1 NAND2X1_433 ( .A(_3636__32_), .B(_1031__bF_buf47), .Y(_2752_) );
OAI21X1 OAI21X1_1067 ( .A(_1031__bF_buf47), .B(_2751_), .C(_2752_), .Y(_773_) );
INVX2 INVX2_74 ( .A(bundleAddress_i[31]), .Y(_2753_) );
NAND2X1 NAND2X1_434 ( .A(_3636__31_), .B(_1031__bF_buf7), .Y(_2754_) );
OAI21X1 OAI21X1_1068 ( .A(_1031__bF_buf7), .B(_2753_), .C(_2754_), .Y(_774_) );
INVX2 INVX2_75 ( .A(bundleAddress_i[30]), .Y(_2755_) );
NAND2X1 NAND2X1_435 ( .A(_3636__30_), .B(_1031__bF_buf7), .Y(_2756_) );
OAI21X1 OAI21X1_1069 ( .A(_1031__bF_buf7), .B(_2755_), .C(_2756_), .Y(_775_) );
INVX4 INVX4_40 ( .A(bundleAddress_i[29]), .Y(_2757_) );
NAND2X1 NAND2X1_436 ( .A(_3636__29_), .B(_1031__bF_buf64), .Y(_2758_) );
OAI21X1 OAI21X1_1070 ( .A(_1031__bF_buf64), .B(_2757_), .C(_2758_), .Y(_776_) );
INVX2 INVX2_76 ( .A(bundleAddress_i[28]), .Y(_2759_) );
NAND2X1 NAND2X1_437 ( .A(_3636__28_), .B(_1031__bF_buf4), .Y(_2760_) );
OAI21X1 OAI21X1_1071 ( .A(_1031__bF_buf4), .B(_2759_), .C(_2760_), .Y(_777_) );
INVX2 INVX2_77 ( .A(bundleAddress_i[27]), .Y(_2761_) );
NAND2X1 NAND2X1_438 ( .A(_3636__27_), .B(_1031__bF_buf38), .Y(_2762_) );
OAI21X1 OAI21X1_1072 ( .A(_1031__bF_buf18), .B(_2761_), .C(_2762_), .Y(_778_) );
INVX4 INVX4_41 ( .A(bundleAddress_i[26]), .Y(_2763_) );
NAND2X1 NAND2X1_439 ( .A(_3636__26_), .B(_1031__bF_buf18), .Y(_2764_) );
OAI21X1 OAI21X1_1073 ( .A(_1031__bF_buf18), .B(_2763_), .C(_2764_), .Y(_779_) );
INVX2 INVX2_78 ( .A(bundleAddress_i[25]), .Y(_2765_) );
NAND2X1 NAND2X1_440 ( .A(_3636__25_), .B(_1031__bF_buf4), .Y(_2766_) );
OAI21X1 OAI21X1_1074 ( .A(_1031__bF_buf4), .B(_2765_), .C(_2766_), .Y(_780_) );
INVX8 INVX8_3 ( .A(bundleAddress_i[24]), .Y(_2767_) );
NAND2X1 NAND2X1_441 ( .A(_3636__24_), .B(_1031__bF_buf38), .Y(_2768_) );
OAI21X1 OAI21X1_1075 ( .A(_1031__bF_buf38), .B(_2767_), .C(_2768_), .Y(_781_) );
INVX2 INVX2_79 ( .A(bundleAddress_i[23]), .Y(_2769_) );
NAND2X1 NAND2X1_442 ( .A(_3636__23_), .B(_1031__bF_buf38), .Y(_2770_) );
OAI21X1 OAI21X1_1076 ( .A(_1031__bF_buf38), .B(_2769_), .C(_2770_), .Y(_782_) );
INVX4 INVX4_42 ( .A(bundleAddress_i[22]), .Y(_2771_) );
NAND2X1 NAND2X1_443 ( .A(_3636__22_), .B(_1031__bF_buf4), .Y(_2772_) );
OAI21X1 OAI21X1_1077 ( .A(_1031__bF_buf38), .B(_2771_), .C(_2772_), .Y(_783_) );
INVX2 INVX2_80 ( .A(bundleAddress_i[21]), .Y(_2773_) );
NAND2X1 NAND2X1_444 ( .A(_3636__21_), .B(_1031__bF_buf46), .Y(_2774_) );
OAI21X1 OAI21X1_1078 ( .A(_1031__bF_buf46), .B(_2773_), .C(_2774_), .Y(_784_) );
INVX4 INVX4_43 ( .A(bundleAddress_i[20]), .Y(_2775_) );
NAND2X1 NAND2X1_445 ( .A(_3636__20_), .B(_1031__bF_buf44), .Y(_2776_) );
OAI21X1 OAI21X1_1079 ( .A(_1031__bF_buf44), .B(_2775_), .C(_2776_), .Y(_785_) );
INVX1 INVX1_177 ( .A(bundleAddress_i[19]), .Y(_2777_) );
NAND2X1 NAND2X1_446 ( .A(_3636__19_), .B(_1031__bF_buf7), .Y(_2778_) );
OAI21X1 OAI21X1_1080 ( .A(_1031__bF_buf7), .B(_2777_), .C(_2778_), .Y(_786_) );
INVX2 INVX2_81 ( .A(bundleAddress_i[18]), .Y(_2779_) );
NAND2X1 NAND2X1_447 ( .A(_3636__18_), .B(_1031__bF_buf7), .Y(_2780_) );
OAI21X1 OAI21X1_1081 ( .A(_1031__bF_buf46), .B(_2779_), .C(_2780_), .Y(_787_) );
INVX1 INVX1_178 ( .A(bundleAddress_i[17]), .Y(_2781_) );
NAND2X1 NAND2X1_448 ( .A(_3636__17_), .B(_1031__bF_buf28), .Y(_2782_) );
OAI21X1 OAI21X1_1082 ( .A(_1031__bF_buf28), .B(_2781_), .C(_2782_), .Y(_788_) );
INVX2 INVX2_82 ( .A(bundleAddress_i[16]), .Y(_2783_) );
NAND2X1 NAND2X1_449 ( .A(_3636__16_), .B(_1031__bF_buf49), .Y(_2784_) );
OAI21X1 OAI21X1_1083 ( .A(_1031__bF_buf49), .B(_2783_), .C(_2784_), .Y(_789_) );
INVX1 INVX1_179 ( .A(bundleAddress_i[15]), .Y(_2785_) );
NAND2X1 NAND2X1_450 ( .A(_3636__15_), .B(_1031__bF_buf40), .Y(_2786_) );
OAI21X1 OAI21X1_1084 ( .A(_1031__bF_buf13), .B(_2785_), .C(_2786_), .Y(_790_) );
INVX2 INVX2_83 ( .A(bundleAddress_i[14]), .Y(_2787_) );
NAND2X1 NAND2X1_451 ( .A(_3636__14_), .B(_1031__bF_buf46), .Y(_2788_) );
OAI21X1 OAI21X1_1085 ( .A(_1031__bF_buf46), .B(_2787_), .C(_2788_), .Y(_791_) );
INVX4 INVX4_44 ( .A(bundleAddress_i[13]), .Y(_2789_) );
NAND2X1 NAND2X1_452 ( .A(_3636__13_), .B(_1031__bF_buf24), .Y(_2790_) );
OAI21X1 OAI21X1_1086 ( .A(_1031__bF_buf24), .B(_2789_), .C(_2790_), .Y(_792_) );
INVX2 INVX2_84 ( .A(bundleAddress_i[12]), .Y(_2791_) );
NAND2X1 NAND2X1_453 ( .A(_3636__12_), .B(_1031__bF_buf24), .Y(_2792_) );
OAI21X1 OAI21X1_1087 ( .A(_1031__bF_buf24), .B(_2791_), .C(_2792_), .Y(_793_) );
INVX2 INVX2_85 ( .A(bundleAddress_i[11]), .Y(_2793_) );
NAND2X1 NAND2X1_454 ( .A(_3636__11_), .B(_1031__bF_buf24), .Y(_2794_) );
OAI21X1 OAI21X1_1088 ( .A(_1031__bF_buf24), .B(_2793_), .C(_2794_), .Y(_794_) );
INVX2 INVX2_86 ( .A(bundleAddress_i[10]), .Y(_2795_) );
NAND2X1 NAND2X1_455 ( .A(_3636__10_), .B(_1031__bF_buf57), .Y(_2796_) );
OAI21X1 OAI21X1_1089 ( .A(_1031__bF_buf57), .B(_2795_), .C(_2796_), .Y(_795_) );
INVX2 INVX2_87 ( .A(bundleAddress_i[9]), .Y(_2797_) );
NAND2X1 NAND2X1_456 ( .A(_3636__9_), .B(_1031__bF_buf14), .Y(_2798_) );
OAI21X1 OAI21X1_1090 ( .A(_1031__bF_buf14), .B(_2797_), .C(_2798_), .Y(_796_) );
INVX4 INVX4_45 ( .A(bundleAddress_i[8]), .Y(_2799_) );
NAND2X1 NAND2X1_457 ( .A(_3636__8_), .B(_1031__bF_buf31), .Y(_2800_) );
OAI21X1 OAI21X1_1091 ( .A(_1031__bF_buf31), .B(_2799_), .C(_2800_), .Y(_797_) );
INVX2 INVX2_88 ( .A(bundleAddress_i[7]), .Y(_2801_) );
NAND2X1 NAND2X1_458 ( .A(_3636__7_), .B(_1031__bF_buf45), .Y(_2802_) );
OAI21X1 OAI21X1_1092 ( .A(_1031__bF_buf45), .B(_2801_), .C(_2802_), .Y(_798_) );
INVX1 INVX1_180 ( .A(bundleAddress_i[6]), .Y(_2803_) );
NAND2X1 NAND2X1_459 ( .A(_3636__6_), .B(_1031__bF_buf14), .Y(_2804_) );
OAI21X1 OAI21X1_1093 ( .A(_1031__bF_buf45), .B(_2803_), .C(_2804_), .Y(_799_) );
INVX2 INVX2_89 ( .A(bundleAddress_i[5]), .Y(_2805_) );
NAND2X1 NAND2X1_460 ( .A(_3636__5_), .B(_1031__bF_buf58), .Y(_2806_) );
OAI21X1 OAI21X1_1094 ( .A(_1031__bF_buf58), .B(_2805_), .C(_2806_), .Y(_800_) );
INVX2 INVX2_90 ( .A(bundleAddress_i[4]), .Y(_2807_) );
NAND2X1 NAND2X1_461 ( .A(_3636__4_), .B(_1031__bF_buf40), .Y(_2808_) );
OAI21X1 OAI21X1_1095 ( .A(_1031__bF_buf28), .B(_2807_), .C(_2808_), .Y(_801_) );
INVX1 INVX1_181 ( .A(bundleAddress_i[3]), .Y(_2809_) );
NAND2X1 NAND2X1_462 ( .A(_3636__3_), .B(_1031__bF_buf58), .Y(_2810_) );
OAI21X1 OAI21X1_1096 ( .A(_1031__bF_buf31), .B(_2809_), .C(_2810_), .Y(_802_) );
INVX2 INVX2_91 ( .A(bundleAddress_i[2]), .Y(_2811_) );
NAND2X1 NAND2X1_463 ( .A(_3636__2_), .B(_1031__bF_buf31), .Y(_2812_) );
OAI21X1 OAI21X1_1097 ( .A(_1031__bF_buf31), .B(_2811_), .C(_2812_), .Y(_803_) );
INVX2 INVX2_92 ( .A(bundleAddress_i[1]), .Y(_2813_) );
NAND2X1 NAND2X1_464 ( .A(_3636__1_), .B(_1031__bF_buf49), .Y(_2814_) );
OAI21X1 OAI21X1_1098 ( .A(_1031__bF_buf28), .B(_2813_), .C(_2814_), .Y(_804_) );
INVX4 INVX4_46 ( .A(bundleAddress_i[0]), .Y(_2815_) );
NAND2X1 NAND2X1_465 ( .A(_3636__0_), .B(_1031__bF_buf28), .Y(_2816_) );
OAI21X1 OAI21X1_1099 ( .A(_1031__bF_buf28), .B(_2815_), .C(_2816_), .Y(_805_) );
NAND2X1 NAND2X1_466 ( .A(_3637__63_), .B(_1039__bF_buf3), .Y(_2817_) );
OAI21X1 OAI21X1_1100 ( .A(_2689_), .B(_1039__bF_buf3), .C(_2817_), .Y(_806_) );
NAND2X1 NAND2X1_467 ( .A(_3637__62_), .B(_1039__bF_buf7), .Y(_2818_) );
OAI21X1 OAI21X1_1101 ( .A(_2691_), .B(_1039__bF_buf7), .C(_2818_), .Y(_807_) );
NAND2X1 NAND2X1_468 ( .A(_3637__61_), .B(_1039__bF_buf40), .Y(_2819_) );
OAI21X1 OAI21X1_1102 ( .A(bundleAddress_i[61]), .B(_1039__bF_buf21), .C(_2819_), .Y(_808_) );
INVX1 INVX1_182 ( .A(_3637__60_), .Y(_2820_) );
NOR2X1 NOR2X1_121 ( .A(_2693_), .B(_2695_), .Y(_2821_) );
NOR2X1 NOR2X1_122 ( .A(bundleAddress_i[61]), .B(bundleAddress_i[60]), .Y(_2822_) );
NOR2X1 NOR2X1_123 ( .A(_2822_), .B(_2821_), .Y(_2823_) );
NAND2X1 NAND2X1_469 ( .A(_611__bF_buf7), .B(_2823_), .Y(_2824_) );
OAI21X1 OAI21X1_1103 ( .A(_2820_), .B(_611__bF_buf7), .C(_2824_), .Y(_809_) );
NAND2X1 NAND2X1_470 ( .A(bundleAddress_i[60]), .B(bundleAddress_i[59]), .Y(_2825_) );
OAI21X1 OAI21X1_1104 ( .A(_2693_), .B(_2695_), .C(_2697_), .Y(_2826_) );
OAI21X1 OAI21X1_1105 ( .A(_2693_), .B(_2825_), .C(_2826_), .Y(_2827_) );
NAND2X1 NAND2X1_471 ( .A(_3637__59_), .B(_1039__bF_buf21), .Y(_2828_) );
OAI21X1 OAI21X1_1106 ( .A(_2827_), .B(_1039__bF_buf21), .C(_2828_), .Y(_810_) );
INVX1 INVX1_183 ( .A(_2825_), .Y(_2829_) );
AOI21X1 AOI21X1_36 ( .A(bundleAddress_i[61]), .B(_2829_), .C(bundleAddress_i[58]), .Y(_2830_) );
INVX1 INVX1_184 ( .A(_2821_), .Y(_2831_) );
NAND2X1 NAND2X1_472 ( .A(bundleAddress_i[59]), .B(bundleAddress_i[58]), .Y(_2832_) );
OAI21X1 OAI21X1_1107 ( .A(_2831_), .B(_2832_), .C(_611__bF_buf4), .Y(_2833_) );
NAND2X1 NAND2X1_473 ( .A(_3637__58_), .B(_1039__bF_buf39), .Y(_2834_) );
OAI21X1 OAI21X1_1108 ( .A(_2833_), .B(_2830_), .C(_2834_), .Y(_811_) );
NAND2X1 NAND2X1_474 ( .A(bundleAddress_i[58]), .B(bundleAddress_i[57]), .Y(_2835_) );
NOR2X1 NOR2X1_124 ( .A(_2825_), .B(_2835_), .Y(_2836_) );
INVX4 INVX4_47 ( .A(_2836_), .Y(_2837_) );
OAI21X1 OAI21X1_1109 ( .A(_2831_), .B(_2832_), .C(_2701_), .Y(_2838_) );
OAI21X1 OAI21X1_1110 ( .A(_2837_), .B(_2693_), .C(_2838_), .Y(_2839_) );
NAND2X1 NAND2X1_475 ( .A(_3637__57_), .B(_1039__bF_buf39), .Y(_2840_) );
OAI21X1 OAI21X1_1111 ( .A(_2839_), .B(_1039__bF_buf39), .C(_2840_), .Y(_812_) );
INVX1 INVX1_185 ( .A(_2832_), .Y(_2841_) );
NAND2X1 NAND2X1_476 ( .A(_2841_), .B(_2821_), .Y(_2842_) );
OAI21X1 OAI21X1_1112 ( .A(_2842_), .B(_2701_), .C(_2703_), .Y(_2843_) );
NAND2X1 NAND2X1_477 ( .A(bundleAddress_i[57]), .B(bundleAddress_i[56]), .Y(_2844_) );
OAI21X1 OAI21X1_1113 ( .A(_2842_), .B(_2844_), .C(_2843_), .Y(_2845_) );
NAND2X1 NAND2X1_478 ( .A(_3637__56_), .B(_1039__bF_buf21), .Y(_2846_) );
OAI21X1 OAI21X1_1114 ( .A(_2845_), .B(_1039__bF_buf21), .C(_2846_), .Y(_813_) );
NAND2X1 NAND2X1_479 ( .A(_3637__55_), .B(_1039__bF_buf39), .Y(_2847_) );
NAND2X1 NAND2X1_480 ( .A(bundleAddress_i[56]), .B(bundleAddress_i[55]), .Y(_2848_) );
NOR2X1 NOR2X1_125 ( .A(_2848_), .B(_2837_), .Y(_2849_) );
INVX2 INVX2_93 ( .A(_2849_), .Y(_2850_) );
NOR2X1 NOR2X1_126 ( .A(_2693_), .B(_2850_), .Y(_2851_) );
OAI21X1 OAI21X1_1115 ( .A(_2842_), .B(_2844_), .C(_2705_), .Y(_2852_) );
NAND2X1 NAND2X1_481 ( .A(_611__bF_buf4), .B(_2852_), .Y(_2853_) );
OAI21X1 OAI21X1_1116 ( .A(_2851_), .B(_2853_), .C(_2847_), .Y(_814_) );
OAI21X1 OAI21X1_1117 ( .A(_2850_), .B(_2693_), .C(_2707_), .Y(_2854_) );
NAND2X1 NAND2X1_482 ( .A(bundleAddress_i[55]), .B(bundleAddress_i[54]), .Y(_2855_) );
NOR2X1 NOR2X1_127 ( .A(_2844_), .B(_2855_), .Y(_2856_) );
INVX2 INVX2_94 ( .A(_2856_), .Y(_2857_) );
OAI21X1 OAI21X1_1118 ( .A(_2842_), .B(_2857_), .C(_2854_), .Y(_2858_) );
NAND2X1 NAND2X1_483 ( .A(_3637__54_), .B(_1039__bF_buf33), .Y(_2859_) );
OAI21X1 OAI21X1_1119 ( .A(_2858_), .B(_1039__bF_buf33), .C(_2859_), .Y(_815_) );
NAND3X1 NAND3X1_38 ( .A(_2821_), .B(_2841_), .C(_2856_), .Y(_2860_) );
NOR2X1 NOR2X1_128 ( .A(_2709_), .B(_2860_), .Y(_2861_) );
INVX1 INVX1_186 ( .A(_2860_), .Y(_2862_) );
OAI21X1 OAI21X1_1120 ( .A(_2862_), .B(bundleAddress_i[53]), .C(_611__bF_buf4), .Y(_2863_) );
NAND2X1 NAND2X1_484 ( .A(_3637__53_), .B(_1039__bF_buf6), .Y(_2864_) );
OAI21X1 OAI21X1_1121 ( .A(_2863_), .B(_2861_), .C(_2864_), .Y(_816_) );
XNOR2X1 XNOR2X1_56 ( .A(_2861_), .B(bundleAddress_i[52]), .Y(_2865_) );
NAND2X1 NAND2X1_485 ( .A(_3637__52_), .B(_1039__bF_buf6), .Y(_2866_) );
OAI21X1 OAI21X1_1122 ( .A(_2865_), .B(_1039__bF_buf6), .C(_2866_), .Y(_817_) );
NAND2X1 NAND2X1_486 ( .A(_3637__51_), .B(_1039__bF_buf6), .Y(_2867_) );
INVX2 INVX2_95 ( .A(_2861_), .Y(_2868_) );
NAND2X1 NAND2X1_487 ( .A(bundleAddress_i[52]), .B(bundleAddress_i[51]), .Y(_2869_) );
NOR2X1 NOR2X1_129 ( .A(_2869_), .B(_2868_), .Y(_2870_) );
OAI21X1 OAI21X1_1123 ( .A(_2868_), .B(_2711_), .C(_2713_), .Y(_2871_) );
NAND2X1 NAND2X1_488 ( .A(_611__bF_buf4), .B(_2871_), .Y(_2872_) );
OAI21X1 OAI21X1_1124 ( .A(_2872_), .B(_2870_), .C(_2867_), .Y(_818_) );
OAI21X1 OAI21X1_1125 ( .A(_2868_), .B(_2869_), .C(_2715_), .Y(_2873_) );
NAND2X1 NAND2X1_489 ( .A(bundleAddress_i[50]), .B(_2870_), .Y(_2874_) );
NAND2X1 NAND2X1_490 ( .A(_2873_), .B(_2874_), .Y(_2875_) );
NAND2X1 NAND2X1_491 ( .A(_3637__50_), .B(_1039__bF_buf2), .Y(_2876_) );
OAI21X1 OAI21X1_1126 ( .A(_2875_), .B(_1039__bF_buf2), .C(_2876_), .Y(_819_) );
NAND2X1 NAND2X1_492 ( .A(_2717_), .B(_2874_), .Y(_2877_) );
INVX2 INVX2_96 ( .A(_2869_), .Y(_2878_) );
NAND3X1 NAND3X1_39 ( .A(bundleAddress_i[50]), .B(bundleAddress_i[49]), .C(_2878_), .Y(_2879_) );
OAI21X1 OAI21X1_1127 ( .A(_2868_), .B(_2879_), .C(_2877_), .Y(_2880_) );
NAND2X1 NAND2X1_493 ( .A(_3637__49_), .B(_1039__bF_buf2), .Y(_2881_) );
OAI21X1 OAI21X1_1128 ( .A(_2880_), .B(_1039__bF_buf2), .C(_2881_), .Y(_820_) );
NAND2X1 NAND2X1_494 ( .A(bundleAddress_i[53]), .B(bundleAddress_i[50]), .Y(_2882_) );
NOR2X1 NOR2X1_130 ( .A(_2869_), .B(_2882_), .Y(_2883_) );
NAND2X1 NAND2X1_495 ( .A(_2883_), .B(_2862_), .Y(_2884_) );
NOR2X1 NOR2X1_131 ( .A(_2717_), .B(_2884_), .Y(_2885_) );
XNOR2X1 XNOR2X1_57 ( .A(_2885_), .B(bundleAddress_i[48]), .Y(_2886_) );
NAND2X1 NAND2X1_496 ( .A(_3637__48_), .B(_1039__bF_buf27), .Y(_2887_) );
OAI21X1 OAI21X1_1129 ( .A(_2886_), .B(_1039__bF_buf13), .C(_2887_), .Y(_821_) );
NAND2X1 NAND2X1_497 ( .A(bundleAddress_i[49]), .B(bundleAddress_i[48]), .Y(_2888_) );
OR2X2 OR2X2_16 ( .A(_2884_), .B(_2888_), .Y(_2889_) );
XNOR2X1 XNOR2X1_58 ( .A(_2889_), .B(_2721_), .Y(_2890_) );
NAND2X1 NAND2X1_498 ( .A(_3637__47_), .B(_1039__bF_buf14), .Y(_2891_) );
OAI21X1 OAI21X1_1130 ( .A(_2890_), .B(_1039__bF_buf27), .C(_2891_), .Y(_822_) );
NAND2X1 NAND2X1_499 ( .A(_3637__46_), .B(_1039__bF_buf27), .Y(_2892_) );
NOR2X1 NOR2X1_132 ( .A(_2721_), .B(_2889_), .Y(_2893_) );
XNOR2X1 XNOR2X1_59 ( .A(_2893_), .B(bundleAddress_i[46]), .Y(_2894_) );
OAI21X1 OAI21X1_1131 ( .A(_2894_), .B(_1039__bF_buf27), .C(_2892_), .Y(_823_) );
NAND2X1 NAND2X1_500 ( .A(bundleAddress_i[47]), .B(bundleAddress_i[46]), .Y(_2895_) );
NOR2X1 NOR2X1_133 ( .A(_2888_), .B(_2895_), .Y(_2896_) );
NAND2X1 NAND2X1_501 ( .A(_2883_), .B(_2896_), .Y(_2897_) );
NOR2X1 NOR2X1_134 ( .A(_2897_), .B(_2860_), .Y(_2898_) );
NAND2X1 NAND2X1_502 ( .A(bundleAddress_i[45]), .B(_2898_), .Y(_2899_) );
INVX1 INVX1_187 ( .A(_2899_), .Y(_2900_) );
OAI21X1 OAI21X1_1132 ( .A(_2898_), .B(bundleAddress_i[45]), .C(_611__bF_buf6), .Y(_2901_) );
NAND2X1 NAND2X1_503 ( .A(_3637__45_), .B(_1039__bF_buf9), .Y(_2902_) );
OAI21X1 OAI21X1_1133 ( .A(_2900_), .B(_2901_), .C(_2902_), .Y(_824_) );
XNOR2X1 XNOR2X1_60 ( .A(_2899_), .B(_2727_), .Y(_2903_) );
NAND2X1 NAND2X1_504 ( .A(_3637__44_), .B(_1039__bF_buf51), .Y(_2904_) );
OAI21X1 OAI21X1_1134 ( .A(_2903_), .B(_1039__bF_buf51), .C(_2904_), .Y(_825_) );
NAND2X1 NAND2X1_505 ( .A(bundleAddress_i[44]), .B(bundleAddress_i[43]), .Y(_2905_) );
NOR2X1 NOR2X1_135 ( .A(_2905_), .B(_2899_), .Y(_2906_) );
INVX1 INVX1_188 ( .A(_2898_), .Y(_2907_) );
NOR2X1 NOR2X1_136 ( .A(_2725_), .B(_2727_), .Y(_2908_) );
INVX2 INVX2_97 ( .A(_2908_), .Y(_2909_) );
NOR2X1 NOR2X1_137 ( .A(_2909_), .B(_2907_), .Y(_2910_) );
OAI21X1 OAI21X1_1135 ( .A(_2910_), .B(bundleAddress_i[43]), .C(_611__bF_buf6), .Y(_2911_) );
NAND2X1 NAND2X1_506 ( .A(_3637__43_), .B(_1039__bF_buf45), .Y(_2912_) );
OAI21X1 OAI21X1_1136 ( .A(_2911_), .B(_2906_), .C(_2912_), .Y(_826_) );
NOR2X1 NOR2X1_138 ( .A(bundleAddress_i[42]), .B(_2906_), .Y(_2913_) );
NAND2X1 NAND2X1_507 ( .A(bundleAddress_i[43]), .B(_2910_), .Y(_2914_) );
OAI21X1 OAI21X1_1137 ( .A(_2914_), .B(_2731_), .C(_611__bF_buf6), .Y(_2915_) );
NAND2X1 NAND2X1_508 ( .A(_3637__42_), .B(_1039__bF_buf45), .Y(_2916_) );
OAI21X1 OAI21X1_1138 ( .A(_2915_), .B(_2913_), .C(_2916_), .Y(_827_) );
OAI21X1 OAI21X1_1139 ( .A(_2914_), .B(_2731_), .C(_2733_), .Y(_2917_) );
NAND2X1 NAND2X1_509 ( .A(bundleAddress_i[42]), .B(bundleAddress_i[41]), .Y(_2918_) );
OR2X2 OR2X2_17 ( .A(_2905_), .B(_2918_), .Y(_2919_) );
OAI21X1 OAI21X1_1140 ( .A(_2899_), .B(_2919_), .C(_2917_), .Y(_2920_) );
NAND2X1 NAND2X1_510 ( .A(_3637__41_), .B(_1039__bF_buf51), .Y(_2921_) );
OAI21X1 OAI21X1_1141 ( .A(_2920_), .B(_1039__bF_buf51), .C(_2921_), .Y(_828_) );
NOR2X1 NOR2X1_139 ( .A(_2919_), .B(_2899_), .Y(_2922_) );
XNOR2X1 XNOR2X1_61 ( .A(_2922_), .B(bundleAddress_i[40]), .Y(_2923_) );
NAND2X1 NAND2X1_511 ( .A(_3637__40_), .B(_1039__bF_buf45), .Y(_2924_) );
OAI21X1 OAI21X1_1142 ( .A(_2923_), .B(_1039__bF_buf45), .C(_2924_), .Y(_829_) );
NAND2X1 NAND2X1_512 ( .A(bundleAddress_i[45]), .B(bundleAddress_i[42]), .Y(_2925_) );
NOR2X1 NOR2X1_140 ( .A(_2905_), .B(_2925_), .Y(_2926_) );
NAND2X1 NAND2X1_513 ( .A(_2926_), .B(_2898_), .Y(_2927_) );
NAND2X1 NAND2X1_514 ( .A(bundleAddress_i[41]), .B(bundleAddress_i[40]), .Y(_2928_) );
NOR2X1 NOR2X1_141 ( .A(_2928_), .B(_2927_), .Y(_2929_) );
XNOR2X1 XNOR2X1_62 ( .A(_2929_), .B(bundleAddress_i[39]), .Y(_2930_) );
NAND2X1 NAND2X1_515 ( .A(_3637__39_), .B(_1039__bF_buf17), .Y(_2931_) );
OAI21X1 OAI21X1_1143 ( .A(_2930_), .B(_1039__bF_buf35), .C(_2931_), .Y(_830_) );
NAND2X1 NAND2X1_516 ( .A(_3637__38_), .B(_1039__bF_buf8), .Y(_2932_) );
NAND2X1 NAND2X1_517 ( .A(bundleAddress_i[39]), .B(_2929_), .Y(_2933_) );
XNOR2X1 XNOR2X1_63 ( .A(_2933_), .B(_2739_), .Y(_2934_) );
OAI21X1 OAI21X1_1144 ( .A(_2934_), .B(_1039__bF_buf8), .C(_2932_), .Y(_831_) );
NAND2X1 NAND2X1_518 ( .A(bundleAddress_i[39]), .B(bundleAddress_i[38]), .Y(_2935_) );
NOR2X1 NOR2X1_142 ( .A(_2928_), .B(_2935_), .Y(_2936_) );
NAND2X1 NAND2X1_519 ( .A(_2926_), .B(_2936_), .Y(_2937_) );
INVX1 INVX1_189 ( .A(_2937_), .Y(_2938_) );
NAND2X1 NAND2X1_520 ( .A(_2938_), .B(_2898_), .Y(_2939_) );
NOR2X1 NOR2X1_143 ( .A(_2741_), .B(_2939_), .Y(_2940_) );
INVX1 INVX1_190 ( .A(_2939_), .Y(_2941_) );
OAI21X1 OAI21X1_1145 ( .A(_2941_), .B(bundleAddress_i[37]), .C(_611__bF_buf7), .Y(_2942_) );
NAND2X1 NAND2X1_521 ( .A(_3637__37_), .B(_1039__bF_buf8), .Y(_2943_) );
OAI21X1 OAI21X1_1146 ( .A(_2942_), .B(_2940_), .C(_2943_), .Y(_832_) );
XNOR2X1 XNOR2X1_64 ( .A(_2940_), .B(bundleAddress_i[36]), .Y(_2944_) );
NAND2X1 NAND2X1_522 ( .A(_3637__36_), .B(_1039__bF_buf8), .Y(_2945_) );
OAI21X1 OAI21X1_1147 ( .A(_2944_), .B(_1039__bF_buf8), .C(_2945_), .Y(_833_) );
NAND2X1 NAND2X1_523 ( .A(bundleAddress_i[37]), .B(bundleAddress_i[36]), .Y(_2946_) );
NOR2X1 NOR2X1_144 ( .A(_2946_), .B(_2939_), .Y(_2947_) );
XNOR2X1 XNOR2X1_65 ( .A(_2947_), .B(bundleAddress_i[35]), .Y(_2948_) );
NAND2X1 NAND2X1_524 ( .A(_3637__35_), .B(_1039__bF_buf28), .Y(_2949_) );
OAI21X1 OAI21X1_1148 ( .A(_2948_), .B(_1039__bF_buf28), .C(_2949_), .Y(_834_) );
NAND2X1 NAND2X1_525 ( .A(_3637__34_), .B(_1039__bF_buf35), .Y(_2950_) );
NAND2X1 NAND2X1_526 ( .A(bundleAddress_i[35]), .B(_2947_), .Y(_2951_) );
XNOR2X1 XNOR2X1_66 ( .A(_2951_), .B(_2747_), .Y(_2952_) );
OAI21X1 OAI21X1_1149 ( .A(_2952_), .B(_1039__bF_buf35), .C(_2950_), .Y(_835_) );
NAND3X1 NAND3X1_40 ( .A(bundleAddress_i[37]), .B(bundleAddress_i[36]), .C(bundleAddress_i[35]), .Y(_2953_) );
INVX2 INVX2_98 ( .A(_2953_), .Y(_2954_) );
NAND2X1 NAND2X1_527 ( .A(bundleAddress_i[34]), .B(_2954_), .Y(_2955_) );
NOR2X1 NOR2X1_145 ( .A(_2955_), .B(_2939_), .Y(_2956_) );
NOR2X1 NOR2X1_146 ( .A(bundleAddress_i[33]), .B(_2956_), .Y(_2957_) );
NAND2X1 NAND2X1_528 ( .A(bundleAddress_i[33]), .B(_2956_), .Y(_2958_) );
NAND2X1 NAND2X1_529 ( .A(_611__bF_buf7), .B(_2958_), .Y(_2959_) );
NAND2X1 NAND2X1_530 ( .A(_3637__33_), .B(_1039__bF_buf35), .Y(_2960_) );
OAI21X1 OAI21X1_1150 ( .A(_2959_), .B(_2957_), .C(_2960_), .Y(_836_) );
INVX1 INVX1_191 ( .A(_3637__32_), .Y(_2961_) );
NOR2X1 NOR2X1_147 ( .A(bundleAddress_i[32]), .B(_2958_), .Y(_2962_) );
AOI21X1 AOI21X1_37 ( .A(bundleAddress_i[33]), .B(_2956_), .C(_2751_), .Y(_2963_) );
OAI21X1 OAI21X1_1151 ( .A(_2962_), .B(_2963_), .C(_611__bF_buf7), .Y(_2964_) );
OAI21X1 OAI21X1_1152 ( .A(_2961_), .B(_611__bF_buf7), .C(_2964_), .Y(_837_) );
NAND2X1 NAND2X1_531 ( .A(_3637__31_), .B(_1039__bF_buf35), .Y(_2965_) );
NOR2X1 NOR2X1_148 ( .A(_2751_), .B(_2958_), .Y(_2966_) );
NOR2X1 NOR2X1_149 ( .A(bundleAddress_i[31]), .B(_2966_), .Y(_2967_) );
NOR2X1 NOR2X1_150 ( .A(_2751_), .B(_2753_), .Y(_2968_) );
INVX2 INVX2_99 ( .A(_2968_), .Y(_2969_) );
OAI21X1 OAI21X1_1153 ( .A(_2958_), .B(_2969_), .C(_611__bF_buf7), .Y(_2970_) );
OAI21X1 OAI21X1_1154 ( .A(_2967_), .B(_2970_), .C(_2965_), .Y(_838_) );
NAND2X1 NAND2X1_532 ( .A(_3637__30_), .B(_1039__bF_buf35), .Y(_2971_) );
AOI21X1 AOI21X1_38 ( .A(bundleAddress_i[31]), .B(_2966_), .C(bundleAddress_i[30]), .Y(_2972_) );
NAND3X1 NAND3X1_41 ( .A(bundleAddress_i[32]), .B(bundleAddress_i[31]), .C(bundleAddress_i[30]), .Y(_2973_) );
OAI21X1 OAI21X1_1155 ( .A(_2958_), .B(_2973_), .C(_611__bF_buf7), .Y(_2974_) );
OAI21X1 OAI21X1_1156 ( .A(_2972_), .B(_2974_), .C(_2971_), .Y(_839_) );
INVX1 INVX1_192 ( .A(_2973_), .Y(_2975_) );
NOR2X1 NOR2X1_151 ( .A(_2747_), .B(_2749_), .Y(_2976_) );
NAND3X1 NAND3X1_42 ( .A(_2976_), .B(_2954_), .C(_2975_), .Y(_2977_) );
NOR2X1 NOR2X1_152 ( .A(_2937_), .B(_2977_), .Y(_2978_) );
NAND2X1 NAND2X1_533 ( .A(_2978_), .B(_2898_), .Y(_2979_) );
NOR2X1 NOR2X1_153 ( .A(_2757_), .B(_2979_), .Y(_2980_) );
AND2X2 AND2X2_23 ( .A(_2898_), .B(_2978_), .Y(_2981_) );
OAI21X1 OAI21X1_1157 ( .A(_2981_), .B(bundleAddress_i[29]), .C(_611__bF_buf6), .Y(_2982_) );
NAND2X1 NAND2X1_534 ( .A(_3637__29_), .B(_1039__bF_buf25), .Y(_2983_) );
OAI21X1 OAI21X1_1158 ( .A(_2982_), .B(_2980_), .C(_2983_), .Y(_840_) );
XNOR2X1 XNOR2X1_67 ( .A(_2980_), .B(bundleAddress_i[28]), .Y(_2984_) );
NAND2X1 NAND2X1_535 ( .A(_3637__28_), .B(_1039__bF_buf11), .Y(_2985_) );
OAI21X1 OAI21X1_1159 ( .A(_2984_), .B(_1039__bF_buf11), .C(_2985_), .Y(_841_) );
NAND2X1 NAND2X1_536 ( .A(bundleAddress_i[29]), .B(bundleAddress_i[28]), .Y(_2986_) );
NOR2X1 NOR2X1_154 ( .A(_2986_), .B(_2979_), .Y(_2987_) );
XNOR2X1 XNOR2X1_68 ( .A(_2987_), .B(bundleAddress_i[27]), .Y(_2988_) );
NAND2X1 NAND2X1_537 ( .A(_3637__27_), .B(_1039__bF_buf52), .Y(_2989_) );
OAI21X1 OAI21X1_1160 ( .A(_2988_), .B(_1039__bF_buf52), .C(_2989_), .Y(_842_) );
NAND2X1 NAND2X1_538 ( .A(_3637__26_), .B(_1039__bF_buf25), .Y(_2990_) );
NAND2X1 NAND2X1_539 ( .A(bundleAddress_i[27]), .B(_2987_), .Y(_2991_) );
XNOR2X1 XNOR2X1_69 ( .A(_2991_), .B(_2763_), .Y(_2992_) );
OAI21X1 OAI21X1_1161 ( .A(_2992_), .B(_1039__bF_buf25), .C(_2990_), .Y(_843_) );
NAND2X1 NAND2X1_540 ( .A(bundleAddress_i[28]), .B(bundleAddress_i[27]), .Y(_2993_) );
NAND2X1 NAND2X1_541 ( .A(bundleAddress_i[29]), .B(bundleAddress_i[26]), .Y(_2994_) );
NOR2X1 NOR2X1_155 ( .A(_2993_), .B(_2994_), .Y(_2995_) );
INVX2 INVX2_100 ( .A(_2995_), .Y(_2996_) );
NOR2X1 NOR2X1_156 ( .A(_2996_), .B(_2979_), .Y(_2997_) );
NAND2X1 NAND2X1_542 ( .A(bundleAddress_i[25]), .B(_2997_), .Y(_2998_) );
INVX1 INVX1_193 ( .A(_2998_), .Y(_2999_) );
OAI21X1 OAI21X1_1162 ( .A(_2997_), .B(bundleAddress_i[25]), .C(_611__bF_buf6), .Y(_3000_) );
NAND2X1 NAND2X1_543 ( .A(_3637__25_), .B(_1039__bF_buf11), .Y(_3001_) );
OAI21X1 OAI21X1_1163 ( .A(_2999_), .B(_3000_), .C(_3001_), .Y(_844_) );
XNOR2X1 XNOR2X1_70 ( .A(_2998_), .B(_2767_), .Y(_3002_) );
NAND2X1 NAND2X1_544 ( .A(_3637__24_), .B(_1039__bF_buf48), .Y(_3003_) );
OAI21X1 OAI21X1_1164 ( .A(_3002_), .B(_1039__bF_buf11), .C(_3003_), .Y(_845_) );
NAND2X1 NAND2X1_545 ( .A(_3637__23_), .B(_1039__bF_buf11), .Y(_3004_) );
NAND2X1 NAND2X1_546 ( .A(bundleAddress_i[24]), .B(bundleAddress_i[23]), .Y(_3005_) );
NOR2X1 NOR2X1_157 ( .A(_3005_), .B(_2998_), .Y(_3006_) );
OAI21X1 OAI21X1_1165 ( .A(_2998_), .B(_2767_), .C(_2769_), .Y(_3007_) );
NAND2X1 NAND2X1_547 ( .A(_611__bF_buf6), .B(_3007_), .Y(_3008_) );
OAI21X1 OAI21X1_1166 ( .A(_3008_), .B(_3006_), .C(_3004_), .Y(_846_) );
NAND2X1 NAND2X1_548 ( .A(_3637__22_), .B(_1039__bF_buf11), .Y(_3009_) );
NOR2X1 NOR2X1_158 ( .A(_2765_), .B(_2767_), .Y(_3010_) );
NAND3X1 NAND3X1_43 ( .A(bundleAddress_i[23]), .B(_3010_), .C(_2997_), .Y(_3011_) );
XNOR2X1 XNOR2X1_71 ( .A(_3011_), .B(_2771_), .Y(_3012_) );
OAI21X1 OAI21X1_1167 ( .A(_3012_), .B(_1039__bF_buf11), .C(_3009_), .Y(_847_) );
INVX2 INVX2_101 ( .A(_3005_), .Y(_3013_) );
NOR2X1 NOR2X1_159 ( .A(_2765_), .B(_2771_), .Y(_3014_) );
NAND3X1 NAND3X1_44 ( .A(_3013_), .B(_3014_), .C(_2995_), .Y(_3015_) );
NOR2X1 NOR2X1_160 ( .A(_3015_), .B(_2979_), .Y(_3016_) );
NAND2X1 NAND2X1_549 ( .A(bundleAddress_i[21]), .B(_3016_), .Y(_3017_) );
INVX1 INVX1_194 ( .A(_3017_), .Y(_3018_) );
OAI21X1 OAI21X1_1168 ( .A(_3016_), .B(bundleAddress_i[21]), .C(_611__bF_buf6), .Y(_3019_) );
NAND2X1 NAND2X1_550 ( .A(_3637__21_), .B(_1039__bF_buf25), .Y(_3020_) );
OAI21X1 OAI21X1_1169 ( .A(_3018_), .B(_3019_), .C(_3020_), .Y(_848_) );
XNOR2X1 XNOR2X1_72 ( .A(_3017_), .B(_2775_), .Y(_3021_) );
NAND2X1 NAND2X1_551 ( .A(_3637__20_), .B(_1039__bF_buf35), .Y(_3022_) );
OAI21X1 OAI21X1_1170 ( .A(_3021_), .B(_1039__bF_buf35), .C(_3022_), .Y(_849_) );
NAND2X1 NAND2X1_552 ( .A(_3637__19_), .B(_1039__bF_buf34), .Y(_3023_) );
NAND2X1 NAND2X1_553 ( .A(bundleAddress_i[20]), .B(bundleAddress_i[19]), .Y(_3024_) );
NOR2X1 NOR2X1_161 ( .A(_3024_), .B(_3017_), .Y(_3025_) );
OAI21X1 OAI21X1_1171 ( .A(_3017_), .B(_2775_), .C(_2777_), .Y(_3026_) );
NAND2X1 NAND2X1_554 ( .A(_611__bF_buf7), .B(_3026_), .Y(_3027_) );
OAI21X1 OAI21X1_1172 ( .A(_3027_), .B(_3025_), .C(_3023_), .Y(_850_) );
NAND2X1 NAND2X1_555 ( .A(_3637__18_), .B(_1039__bF_buf34), .Y(_3028_) );
NOR2X1 NOR2X1_162 ( .A(_2773_), .B(_2775_), .Y(_3029_) );
NAND3X1 NAND3X1_45 ( .A(bundleAddress_i[19]), .B(_3029_), .C(_3016_), .Y(_3030_) );
XNOR2X1 XNOR2X1_73 ( .A(_3030_), .B(_2779_), .Y(_3031_) );
OAI21X1 OAI21X1_1173 ( .A(_3031_), .B(_1039__bF_buf34), .C(_3028_), .Y(_851_) );
NAND2X1 NAND2X1_556 ( .A(bundleAddress_i[21]), .B(bundleAddress_i[18]), .Y(_3032_) );
NOR2X1 NOR2X1_163 ( .A(_3024_), .B(_3032_), .Y(_3033_) );
AOI21X1 AOI21X1_39 ( .A(_3033_), .B(_3016_), .C(bundleAddress_i[17]), .Y(_3034_) );
NAND3X1 NAND3X1_46 ( .A(bundleAddress_i[17]), .B(_3033_), .C(_3016_), .Y(_3035_) );
NAND2X1 NAND2X1_557 ( .A(_611__bF_buf2), .B(_3035_), .Y(_3036_) );
NAND2X1 NAND2X1_558 ( .A(_3637__17_), .B(_1039__bF_buf50), .Y(_3037_) );
OAI21X1 OAI21X1_1174 ( .A(_3036_), .B(_3034_), .C(_3037_), .Y(_852_) );
NAND2X1 NAND2X1_559 ( .A(_3637__16_), .B(_1039__bF_buf34), .Y(_3038_) );
INVX2 INVX2_102 ( .A(_3035_), .Y(_3039_) );
NOR2X1 NOR2X1_164 ( .A(bundleAddress_i[16]), .B(_3039_), .Y(_3040_) );
OAI21X1 OAI21X1_1175 ( .A(_3035_), .B(_2783_), .C(_611__bF_buf2), .Y(_3041_) );
OAI21X1 OAI21X1_1176 ( .A(_3040_), .B(_3041_), .C(_3038_), .Y(_853_) );
NAND2X1 NAND2X1_560 ( .A(_3637__15_), .B(_1039__bF_buf34), .Y(_3042_) );
AOI21X1 AOI21X1_40 ( .A(bundleAddress_i[16]), .B(_3039_), .C(bundleAddress_i[15]), .Y(_3043_) );
NAND2X1 NAND2X1_561 ( .A(bundleAddress_i[16]), .B(bundleAddress_i[15]), .Y(_3044_) );
OAI21X1 OAI21X1_1177 ( .A(_3035_), .B(_3044_), .C(_611__bF_buf2), .Y(_3045_) );
OAI21X1 OAI21X1_1178 ( .A(_3043_), .B(_3045_), .C(_3042_), .Y(_854_) );
NAND2X1 NAND2X1_562 ( .A(_3637__14_), .B(_1039__bF_buf50), .Y(_3046_) );
INVX1 INVX1_195 ( .A(_3044_), .Y(_3047_) );
AOI21X1 AOI21X1_41 ( .A(_3047_), .B(_3039_), .C(bundleAddress_i[14]), .Y(_3048_) );
NAND2X1 NAND2X1_563 ( .A(bundleAddress_i[17]), .B(bundleAddress_i[14]), .Y(_3049_) );
NOR2X1 NOR2X1_165 ( .A(_3044_), .B(_3049_), .Y(_3050_) );
NAND2X1 NAND2X1_564 ( .A(_3033_), .B(_3050_), .Y(_3051_) );
NOR2X1 NOR2X1_166 ( .A(_3051_), .B(_3015_), .Y(_3052_) );
NAND2X1 NAND2X1_565 ( .A(_3052_), .B(_2981_), .Y(_3053_) );
NAND2X1 NAND2X1_566 ( .A(_611__bF_buf3), .B(_3053_), .Y(_3054_) );
OAI21X1 OAI21X1_1179 ( .A(_3048_), .B(_3054_), .C(_3046_), .Y(_855_) );
AND2X2 AND2X2_24 ( .A(_2981_), .B(_3052_), .Y(_3055_) );
NOR2X1 NOR2X1_167 ( .A(bundleAddress_i[13]), .B(_3055_), .Y(_3056_) );
OAI21X1 OAI21X1_1180 ( .A(_3053_), .B(_2789_), .C(_611__bF_buf6), .Y(_3057_) );
NAND2X1 NAND2X1_567 ( .A(_3637__13_), .B(_1039__bF_buf25), .Y(_3058_) );
OAI21X1 OAI21X1_1181 ( .A(_3056_), .B(_3057_), .C(_3058_), .Y(_856_) );
NAND3X1 NAND3X1_47 ( .A(bundleAddress_i[13]), .B(bundleAddress_i[12]), .C(_3055_), .Y(_3059_) );
OAI21X1 OAI21X1_1182 ( .A(_3053_), .B(_2789_), .C(_2791_), .Y(_3060_) );
NAND2X1 NAND2X1_568 ( .A(_3060_), .B(_3059_), .Y(_3061_) );
NAND2X1 NAND2X1_569 ( .A(_3637__12_), .B(_1039__bF_buf36), .Y(_3062_) );
OAI21X1 OAI21X1_1183 ( .A(_3061_), .B(_1039__bF_buf36), .C(_3062_), .Y(_857_) );
NAND2X1 NAND2X1_570 ( .A(_3637__11_), .B(_1039__bF_buf36), .Y(_3063_) );
NOR2X1 NOR2X1_168 ( .A(_2791_), .B(_2793_), .Y(_3064_) );
INVX2 INVX2_103 ( .A(_3064_), .Y(_3065_) );
NOR3X1 NOR3X1_12 ( .A(_2789_), .B(_3065_), .C(_3053_), .Y(_3066_) );
NAND2X1 NAND2X1_571 ( .A(bundleAddress_i[13]), .B(bundleAddress_i[12]), .Y(_3067_) );
OAI21X1 OAI21X1_1184 ( .A(_3053_), .B(_3067_), .C(_2793_), .Y(_3068_) );
NAND2X1 NAND2X1_572 ( .A(_611__bF_buf6), .B(_3068_), .Y(_3069_) );
OAI21X1 OAI21X1_1185 ( .A(_3069_), .B(_3066_), .C(_3063_), .Y(_858_) );
NAND2X1 NAND2X1_573 ( .A(_3637__10_), .B(_1039__bF_buf36), .Y(_3070_) );
NOR3X1 NOR3X1_13 ( .A(_2793_), .B(_2795_), .C(_3059_), .Y(_3071_) );
OAI21X1 OAI21X1_1186 ( .A(_3066_), .B(bundleAddress_i[10]), .C(_611__bF_buf3), .Y(_3072_) );
OAI21X1 OAI21X1_1187 ( .A(_3071_), .B(_3072_), .C(_3070_), .Y(_859_) );
NAND2X1 NAND2X1_574 ( .A(bundleAddress_i[13]), .B(_3064_), .Y(_3073_) );
NOR2X1 NOR2X1_169 ( .A(_2795_), .B(_3073_), .Y(_3074_) );
INVX4 INVX4_48 ( .A(_3074_), .Y(_3075_) );
NOR3X1 NOR3X1_14 ( .A(_2797_), .B(_3075_), .C(_3053_), .Y(_3076_) );
OAI21X1 OAI21X1_1188 ( .A(_3053_), .B(_3075_), .C(_2797_), .Y(_3077_) );
NAND2X1 NAND2X1_575 ( .A(_611__bF_buf3), .B(_3077_), .Y(_3078_) );
NAND2X1 NAND2X1_576 ( .A(_3637__9_), .B(_1039__bF_buf36), .Y(_3079_) );
OAI21X1 OAI21X1_1189 ( .A(_3078_), .B(_3076_), .C(_3079_), .Y(_860_) );
NAND2X1 NAND2X1_577 ( .A(_3637__8_), .B(_1039__bF_buf36), .Y(_3080_) );
NOR2X1 NOR2X1_170 ( .A(bundleAddress_i[8]), .B(_3076_), .Y(_3081_) );
NAND3X1 NAND3X1_48 ( .A(bundleAddress_i[9]), .B(_3074_), .C(_3055_), .Y(_3082_) );
OAI21X1 OAI21X1_1190 ( .A(_3082_), .B(_2799_), .C(_611__bF_buf3), .Y(_3083_) );
OAI21X1 OAI21X1_1191 ( .A(_3083_), .B(_3081_), .C(_3080_), .Y(_861_) );
NAND2X1 NAND2X1_578 ( .A(_3637__7_), .B(_1039__bF_buf49), .Y(_3084_) );
AOI21X1 AOI21X1_42 ( .A(bundleAddress_i[8]), .B(_3076_), .C(bundleAddress_i[7]), .Y(_3085_) );
NOR2X1 NOR2X1_171 ( .A(_2799_), .B(_2801_), .Y(_3086_) );
INVX2 INVX2_104 ( .A(_3086_), .Y(_3087_) );
OAI21X1 OAI21X1_1192 ( .A(_3082_), .B(_3087_), .C(_611__bF_buf3), .Y(_3088_) );
OAI21X1 OAI21X1_1193 ( .A(_3088_), .B(_3085_), .C(_3084_), .Y(_862_) );
NAND2X1 NAND2X1_579 ( .A(_3637__6_), .B(_1039__bF_buf36), .Y(_3089_) );
AOI21X1 AOI21X1_43 ( .A(_3086_), .B(_3076_), .C(bundleAddress_i[6]), .Y(_3090_) );
INVX1 INVX1_196 ( .A(_3073_), .Y(_3091_) );
NAND2X1 NAND2X1_580 ( .A(bundleAddress_i[6]), .B(_3086_), .Y(_3092_) );
INVX1 INVX1_197 ( .A(_3092_), .Y(_3093_) );
NOR2X1 NOR2X1_172 ( .A(_2795_), .B(_2797_), .Y(_3094_) );
NAND3X1 NAND3X1_49 ( .A(_3094_), .B(_3091_), .C(_3093_), .Y(_3095_) );
OAI21X1 OAI21X1_1194 ( .A(_3053_), .B(_3095_), .C(_611__bF_buf3), .Y(_3096_) );
OAI21X1 OAI21X1_1195 ( .A(_3090_), .B(_3096_), .C(_3089_), .Y(_863_) );
INVX1 INVX1_198 ( .A(_3095_), .Y(_3097_) );
NAND3X1 NAND3X1_50 ( .A(_3052_), .B(_3097_), .C(_2981_), .Y(_3098_) );
NOR2X1 NOR2X1_173 ( .A(_2805_), .B(_3098_), .Y(_3099_) );
OAI21X1 OAI21X1_1196 ( .A(_3053_), .B(_3095_), .C(_2805_), .Y(_3100_) );
NAND2X1 NAND2X1_581 ( .A(_611__bF_buf3), .B(_3100_), .Y(_3101_) );
NAND2X1 NAND2X1_582 ( .A(_3637__5_), .B(_1039__bF_buf50), .Y(_3102_) );
OAI21X1 OAI21X1_1197 ( .A(_3101_), .B(_3099_), .C(_3102_), .Y(_864_) );
NAND2X1 NAND2X1_583 ( .A(_3637__4_), .B(_1039__bF_buf49), .Y(_3103_) );
NOR2X1 NOR2X1_174 ( .A(bundleAddress_i[4]), .B(_3099_), .Y(_3104_) );
NAND3X1 NAND3X1_51 ( .A(bundleAddress_i[5]), .B(_3097_), .C(_3055_), .Y(_3105_) );
OAI21X1 OAI21X1_1198 ( .A(_3105_), .B(_2807_), .C(_611__bF_buf2), .Y(_3106_) );
OAI21X1 OAI21X1_1199 ( .A(_3106_), .B(_3104_), .C(_3103_), .Y(_865_) );
NAND2X1 NAND2X1_584 ( .A(_3637__3_), .B(_1039__bF_buf50), .Y(_3107_) );
AOI21X1 AOI21X1_44 ( .A(bundleAddress_i[4]), .B(_3099_), .C(bundleAddress_i[3]), .Y(_3108_) );
NOR2X1 NOR2X1_175 ( .A(_2807_), .B(_2809_), .Y(_3109_) );
INVX1 INVX1_199 ( .A(_3109_), .Y(_3110_) );
OAI21X1 OAI21X1_1200 ( .A(_3105_), .B(_3110_), .C(_611__bF_buf3), .Y(_3111_) );
OAI21X1 OAI21X1_1201 ( .A(_3111_), .B(_3108_), .C(_3107_), .Y(_866_) );
NAND2X1 NAND2X1_585 ( .A(_3637__2_), .B(_1039__bF_buf50), .Y(_3112_) );
AOI21X1 AOI21X1_45 ( .A(_3109_), .B(_3099_), .C(bundleAddress_i[2]), .Y(_3113_) );
NAND2X1 NAND2X1_586 ( .A(bundleAddress_i[5]), .B(_3109_), .Y(_3114_) );
NOR2X1 NOR2X1_176 ( .A(_2811_), .B(_3114_), .Y(_3115_) );
INVX4 INVX4_49 ( .A(_3115_), .Y(_3116_) );
OAI21X1 OAI21X1_1202 ( .A(_3098_), .B(_3116_), .C(_611__bF_buf2), .Y(_3117_) );
OAI21X1 OAI21X1_1203 ( .A(_3113_), .B(_3117_), .C(_3112_), .Y(_867_) );
NAND2X1 NAND2X1_587 ( .A(_3637__1_), .B(_1039__bF_buf50), .Y(_3118_) );
NOR3X1 NOR3X1_15 ( .A(_2813_), .B(_3116_), .C(_3098_), .Y(_3119_) );
OAI21X1 OAI21X1_1204 ( .A(_3098_), .B(_3116_), .C(_2813_), .Y(_3120_) );
NAND2X1 NAND2X1_588 ( .A(_611__bF_buf2), .B(_3120_), .Y(_3121_) );
OAI21X1 OAI21X1_1205 ( .A(_3121_), .B(_3119_), .C(_3118_), .Y(_868_) );
NAND2X1 NAND2X1_589 ( .A(_3637__0_), .B(_1039__bF_buf50), .Y(_3122_) );
AND2X2 AND2X2_25 ( .A(_3119_), .B(bundleAddress_i[0]), .Y(_3123_) );
OAI21X1 OAI21X1_1206 ( .A(_3119_), .B(bundleAddress_i[0]), .C(_611__bF_buf2), .Y(_3124_) );
OAI21X1 OAI21X1_1207 ( .A(_3123_), .B(_3124_), .C(_3122_), .Y(_869_) );
OAI21X1 OAI21X1_1208 ( .A(_1100__bF_buf12_bF_buf0), .B(_1031__bF_buf52), .C(_3638__63_), .Y(_3125_) );
OAI21X1 OAI21X1_1209 ( .A(_1101__bF_buf31), .B(_2689_), .C(_3125_), .Y(_870_) );
OAI21X1 OAI21X1_1210 ( .A(_1100__bF_buf11_bF_buf2), .B(_1031__bF_buf22), .C(_3638__62_), .Y(_3126_) );
OAI21X1 OAI21X1_1211 ( .A(_1101__bF_buf54), .B(_2691_), .C(_3126_), .Y(_871_) );
OAI21X1 OAI21X1_1212 ( .A(_1100__bF_buf10_bF_buf2), .B(_1031__bF_buf76), .C(_3638__61_), .Y(_3127_) );
OAI21X1 OAI21X1_1213 ( .A(_1101__bF_buf47), .B(_2693_), .C(_3127_), .Y(_872_) );
OAI21X1 OAI21X1_1214 ( .A(_1100__bF_buf9_bF_buf2), .B(_1031__bF_buf35), .C(_3638__60_), .Y(_3128_) );
OAI21X1 OAI21X1_1215 ( .A(_1101__bF_buf53), .B(bundleAddress_i[60]), .C(_3128_), .Y(_873_) );
NAND2X1 NAND2X1_590 ( .A(_2695_), .B(_2697_), .Y(_3129_) );
NAND2X1 NAND2X1_591 ( .A(_2825_), .B(_3129_), .Y(_3130_) );
OAI21X1 OAI21X1_1216 ( .A(_1100__bF_buf8_bF_buf0), .B(_1031__bF_buf20), .C(_3638__59_), .Y(_3131_) );
OAI21X1 OAI21X1_1217 ( .A(_3130_), .B(_1101__bF_buf53), .C(_3131_), .Y(_874_) );
NOR2X1 NOR2X1_177 ( .A(bundleAddress_i[58]), .B(_2829_), .Y(_3132_) );
OAI21X1 OAI21X1_1218 ( .A(_2699_), .B(_2825_), .C(_612__bF_buf5), .Y(_3133_) );
OAI21X1 OAI21X1_1219 ( .A(_1100__bF_buf7_bF_buf2), .B(_1031__bF_buf6), .C(_3638__58_), .Y(_3134_) );
OAI21X1 OAI21X1_1220 ( .A(_3133_), .B(_3132_), .C(_3134_), .Y(_875_) );
OAI21X1 OAI21X1_1221 ( .A(_2825_), .B(_2699_), .C(_2701_), .Y(_3135_) );
OAI21X1 OAI21X1_1222 ( .A(_2825_), .B(_2835_), .C(_3135_), .Y(_3136_) );
OAI21X1 OAI21X1_1223 ( .A(_1100__bF_buf11), .B(_1031__bF_buf6), .C(_3638__57_), .Y(_3137_) );
OAI21X1 OAI21X1_1224 ( .A(_3136_), .B(_1101__bF_buf53), .C(_3137_), .Y(_876_) );
NOR2X1 NOR2X1_178 ( .A(bundleAddress_i[56]), .B(_2836_), .Y(_3138_) );
OAI21X1 OAI21X1_1225 ( .A(_2837_), .B(_2703_), .C(_612__bF_buf5), .Y(_3139_) );
OAI21X1 OAI21X1_1226 ( .A(_1100__bF_buf11), .B(_1031__bF_buf6), .C(_3638__56_), .Y(_3140_) );
OAI21X1 OAI21X1_1227 ( .A(_3139_), .B(_3138_), .C(_3140_), .Y(_877_) );
OAI21X1 OAI21X1_1228 ( .A(_2837_), .B(_2703_), .C(_2705_), .Y(_3141_) );
OAI21X1 OAI21X1_1229 ( .A(_2837_), .B(_2848_), .C(_3141_), .Y(_3142_) );
OAI21X1 OAI21X1_1230 ( .A(_1100__bF_buf11), .B(_1031__bF_buf6), .C(_3638__55_), .Y(_3143_) );
OAI21X1 OAI21X1_1231 ( .A(_3142_), .B(_1101__bF_buf53), .C(_3143_), .Y(_878_) );
XNOR2X1 XNOR2X1_74 ( .A(_2849_), .B(bundleAddress_i[54]), .Y(_3144_) );
OAI21X1 OAI21X1_1232 ( .A(_1100__bF_buf9), .B(_1031__bF_buf76), .C(_3638__54_), .Y(_3145_) );
OAI21X1 OAI21X1_1233 ( .A(_3144_), .B(_1101__bF_buf47), .C(_3145_), .Y(_879_) );
NOR2X1 NOR2X1_179 ( .A(_2707_), .B(_2850_), .Y(_3146_) );
XNOR2X1 XNOR2X1_75 ( .A(_3146_), .B(bundleAddress_i[53]), .Y(_3147_) );
OAI21X1 OAI21X1_1234 ( .A(_1100__bF_buf4), .B(_1031__bF_buf6), .C(_3638__53_), .Y(_3148_) );
OAI21X1 OAI21X1_1235 ( .A(_3147_), .B(_1101__bF_buf47), .C(_3148_), .Y(_880_) );
NAND2X1 NAND2X1_592 ( .A(bundleAddress_i[54]), .B(bundleAddress_i[53]), .Y(_3149_) );
NOR2X1 NOR2X1_180 ( .A(_2848_), .B(_3149_), .Y(_3150_) );
NAND2X1 NAND2X1_593 ( .A(_2836_), .B(_3150_), .Y(_3151_) );
XNOR2X1 XNOR2X1_76 ( .A(_3151_), .B(_2711_), .Y(_3152_) );
OAI21X1 OAI21X1_1236 ( .A(_1100__bF_buf9), .B(_1031__bF_buf76), .C(_3638__52_), .Y(_3153_) );
OAI21X1 OAI21X1_1237 ( .A(_3152_), .B(_1101__bF_buf33), .C(_3153_), .Y(_881_) );
OAI21X1 OAI21X1_1238 ( .A(_3151_), .B(_2711_), .C(_2713_), .Y(_3154_) );
OAI21X1 OAI21X1_1239 ( .A(_2869_), .B(_3151_), .C(_3154_), .Y(_3155_) );
OAI21X1 OAI21X1_1240 ( .A(_1100__bF_buf0), .B(_1031__bF_buf2), .C(_3638__51_), .Y(_3156_) );
OAI21X1 OAI21X1_1241 ( .A(_3155_), .B(_1101__bF_buf33), .C(_3156_), .Y(_882_) );
NAND2X1 NAND2X1_594 ( .A(bundleAddress_i[50]), .B(_2878_), .Y(_3157_) );
OAI21X1 OAI21X1_1242 ( .A(_3151_), .B(_2869_), .C(_2715_), .Y(_3158_) );
OAI21X1 OAI21X1_1243 ( .A(_3157_), .B(_3151_), .C(_3158_), .Y(_3159_) );
OAI21X1 OAI21X1_1244 ( .A(_1100__bF_buf14_bF_buf3), .B(_1031__bF_buf54), .C(_3638__50_), .Y(_3160_) );
OAI21X1 OAI21X1_1245 ( .A(_3159_), .B(_1101__bF_buf52), .C(_3160_), .Y(_883_) );
OAI21X1 OAI21X1_1246 ( .A(_3151_), .B(_3157_), .C(_2717_), .Y(_3161_) );
OAI21X1 OAI21X1_1247 ( .A(_2879_), .B(_3151_), .C(_3161_), .Y(_3162_) );
OAI21X1 OAI21X1_1248 ( .A(_1100__bF_buf13_bF_buf0), .B(_1031__bF_buf60), .C(_3638__49_), .Y(_3163_) );
OAI21X1 OAI21X1_1249 ( .A(_3162_), .B(_1101__bF_buf33), .C(_3163_), .Y(_884_) );
NOR2X1 NOR2X1_181 ( .A(_2879_), .B(_3151_), .Y(_3164_) );
XNOR2X1 XNOR2X1_77 ( .A(_3164_), .B(bundleAddress_i[48]), .Y(_3165_) );
OAI21X1 OAI21X1_1250 ( .A(_1100__bF_buf12_bF_buf3), .B(_1031__bF_buf48), .C(_3638__48_), .Y(_3166_) );
OAI21X1 OAI21X1_1251 ( .A(_3165_), .B(_1101__bF_buf29), .C(_3166_), .Y(_885_) );
NOR2X1 NOR2X1_182 ( .A(_2719_), .B(_2721_), .Y(_3167_) );
INVX2 INVX2_105 ( .A(_3167_), .Y(_3168_) );
NOR2X1 NOR2X1_183 ( .A(_3157_), .B(_3151_), .Y(_3169_) );
NAND2X1 NAND2X1_595 ( .A(bundleAddress_i[49]), .B(_3169_), .Y(_3170_) );
INVX1 INVX1_200 ( .A(_3164_), .Y(_3171_) );
OAI21X1 OAI21X1_1252 ( .A(_3171_), .B(_2719_), .C(_2721_), .Y(_3172_) );
OAI21X1 OAI21X1_1253 ( .A(_3168_), .B(_3170_), .C(_3172_), .Y(_3173_) );
OAI21X1 OAI21X1_1254 ( .A(_1100__bF_buf11_bF_buf3), .B(_1031__bF_buf29), .C(_3638__47_), .Y(_3174_) );
OAI21X1 OAI21X1_1255 ( .A(_3173_), .B(_1101__bF_buf52), .C(_3174_), .Y(_886_) );
OAI21X1 OAI21X1_1256 ( .A(_3170_), .B(_3168_), .C(_2723_), .Y(_3175_) );
NOR2X1 NOR2X1_184 ( .A(_3168_), .B(_3170_), .Y(_3176_) );
NAND2X1 NAND2X1_596 ( .A(bundleAddress_i[46]), .B(_3176_), .Y(_3177_) );
NAND2X1 NAND2X1_597 ( .A(_3175_), .B(_3177_), .Y(_3178_) );
OAI21X1 OAI21X1_1257 ( .A(_1100__bF_buf10_bF_buf2), .B(_1031__bF_buf48), .C(_3638__46_), .Y(_3179_) );
OAI21X1 OAI21X1_1258 ( .A(_3178_), .B(_1101__bF_buf29), .C(_3179_), .Y(_887_) );
OAI21X1 OAI21X1_1259 ( .A(_1100__bF_buf9_bF_buf2), .B(_1031__bF_buf32), .C(_3638__45_), .Y(_3180_) );
AOI21X1 AOI21X1_46 ( .A(bundleAddress_i[46]), .B(_3176_), .C(bundleAddress_i[45]), .Y(_3181_) );
NAND3X1 NAND3X1_52 ( .A(bundleAddress_i[46]), .B(bundleAddress_i[45]), .C(_3167_), .Y(_3182_) );
OAI21X1 OAI21X1_1260 ( .A(_3170_), .B(_3182_), .C(_612__bF_buf5), .Y(_3183_) );
OAI21X1 OAI21X1_1261 ( .A(_3181_), .B(_3183_), .C(_3180_), .Y(_888_) );
INVX1 INVX1_201 ( .A(_3151_), .Y(_3184_) );
NOR2X1 NOR2X1_185 ( .A(_2879_), .B(_3182_), .Y(_3185_) );
NAND2X1 NAND2X1_598 ( .A(_3184_), .B(_3185_), .Y(_3186_) );
XNOR2X1 XNOR2X1_78 ( .A(_3186_), .B(_2727_), .Y(_3187_) );
OAI21X1 OAI21X1_1262 ( .A(_1100__bF_buf8_bF_buf3), .B(_1031__bF_buf64), .C(_3638__44_), .Y(_3188_) );
OAI21X1 OAI21X1_1263 ( .A(_3187_), .B(_1101__bF_buf50), .C(_3188_), .Y(_889_) );
OAI21X1 OAI21X1_1264 ( .A(_3186_), .B(_2727_), .C(_2729_), .Y(_3189_) );
OAI21X1 OAI21X1_1265 ( .A(_2905_), .B(_3186_), .C(_3189_), .Y(_3190_) );
OAI21X1 OAI21X1_1266 ( .A(_1100__bF_buf7_bF_buf0), .B(_1031__bF_buf64), .C(_3638__43_), .Y(_3191_) );
OAI21X1 OAI21X1_1267 ( .A(_3190_), .B(_1101__bF_buf22), .C(_3191_), .Y(_890_) );
OR2X2 OR2X2_18 ( .A(_2905_), .B(_2731_), .Y(_3192_) );
OAI21X1 OAI21X1_1268 ( .A(_3186_), .B(_2905_), .C(_2731_), .Y(_3193_) );
OAI21X1 OAI21X1_1269 ( .A(_3192_), .B(_3186_), .C(_3193_), .Y(_3194_) );
OAI21X1 OAI21X1_1270 ( .A(_1100__bF_buf1), .B(_1031__bF_buf64), .C(_3638__42_), .Y(_3195_) );
OAI21X1 OAI21X1_1271 ( .A(_3194_), .B(_1101__bF_buf50), .C(_3195_), .Y(_891_) );
NOR2X1 NOR2X1_186 ( .A(_3192_), .B(_3186_), .Y(_3196_) );
NOR2X1 NOR2X1_187 ( .A(bundleAddress_i[41]), .B(_3196_), .Y(_3197_) );
OAI21X1 OAI21X1_1272 ( .A(_3186_), .B(_2919_), .C(_612__bF_buf3), .Y(_3198_) );
OAI21X1 OAI21X1_1273 ( .A(_1100__bF_buf5), .B(_1031__bF_buf17), .C(_3638__41_), .Y(_3199_) );
OAI21X1 OAI21X1_1274 ( .A(_3197_), .B(_3198_), .C(_3199_), .Y(_892_) );
NOR2X1 NOR2X1_188 ( .A(bundleAddress_i[40]), .B(_3198_), .Y(_3200_) );
INVX1 INVX1_202 ( .A(_2928_), .Y(_3201_) );
NAND2X1 NAND2X1_599 ( .A(_3201_), .B(_3196_), .Y(_3202_) );
MUX2X1 MUX2X1_2 ( .A(_3202_), .B(_3638__40_), .S(_612__bF_buf3), .Y(_3203_) );
NOR2X1 NOR2X1_189 ( .A(_3200_), .B(_3203_), .Y(_893_) );
INVX1 INVX1_203 ( .A(_2919_), .Y(_3204_) );
AND2X2 AND2X2_26 ( .A(_3185_), .B(_3184_), .Y(_3205_) );
NAND2X1 NAND2X1_600 ( .A(_3204_), .B(_3205_), .Y(_3206_) );
OAI21X1 OAI21X1_1275 ( .A(_3206_), .B(_2735_), .C(_2737_), .Y(_3207_) );
NAND3X1 NAND3X1_53 ( .A(bundleAddress_i[39]), .B(_3201_), .C(_3196_), .Y(_3208_) );
NAND2X1 NAND2X1_601 ( .A(_3208_), .B(_3207_), .Y(_3209_) );
OAI21X1 OAI21X1_1276 ( .A(_1100__bF_buf5), .B(_1031__bF_buf17), .C(_3638__39_), .Y(_3210_) );
OAI21X1 OAI21X1_1277 ( .A(_3209_), .B(_1101__bF_buf5), .C(_3210_), .Y(_894_) );
OAI21X1 OAI21X1_1278 ( .A(_1100__bF_buf5), .B(_1031__bF_buf17), .C(_3638__38_), .Y(_3211_) );
AND2X2 AND2X2_27 ( .A(_3208_), .B(_2739_), .Y(_3212_) );
OAI21X1 OAI21X1_1279 ( .A(_3208_), .B(_2739_), .C(_612__bF_buf3), .Y(_3213_) );
OAI21X1 OAI21X1_1280 ( .A(_3212_), .B(_3213_), .C(_3211_), .Y(_895_) );
NAND2X1 NAND2X1_602 ( .A(bundleAddress_i[40]), .B(bundleAddress_i[39]), .Y(_3214_) );
INVX1 INVX1_204 ( .A(_3214_), .Y(_3215_) );
NOR2X1 NOR2X1_190 ( .A(_2919_), .B(_3186_), .Y(_3216_) );
NAND3X1 NAND3X1_54 ( .A(bundleAddress_i[38]), .B(_3215_), .C(_3216_), .Y(_3217_) );
XNOR2X1 XNOR2X1_79 ( .A(_3217_), .B(_2741_), .Y(_3218_) );
OAI21X1 OAI21X1_1281 ( .A(_1100__bF_buf7), .B(_1031__bF_buf77), .C(_3638__37_), .Y(_3219_) );
OAI21X1 OAI21X1_1282 ( .A(_3218_), .B(_1101__bF_buf20), .C(_3219_), .Y(_896_) );
NAND2X1 NAND2X1_603 ( .A(bundleAddress_i[38]), .B(bundleAddress_i[37]), .Y(_3220_) );
OR2X2 OR2X2_19 ( .A(_3214_), .B(_3220_), .Y(_3221_) );
NOR2X1 NOR2X1_191 ( .A(_2919_), .B(_3221_), .Y(_3222_) );
INVX1 INVX1_205 ( .A(_3222_), .Y(_3223_) );
NOR2X1 NOR2X1_192 ( .A(_3223_), .B(_3186_), .Y(_3224_) );
XNOR2X1 XNOR2X1_80 ( .A(_3224_), .B(bundleAddress_i[36]), .Y(_3225_) );
OAI21X1 OAI21X1_1283 ( .A(_1100__bF_buf1), .B(_1031__bF_buf44), .C(_3638__36_), .Y(_3226_) );
OAI21X1 OAI21X1_1284 ( .A(_3225_), .B(_1101__bF_buf13), .C(_3226_), .Y(_897_) );
OAI21X1 OAI21X1_1285 ( .A(_1100__bF_buf5), .B(_1031__bF_buf71), .C(_3638__35_), .Y(_3227_) );
NOR2X1 NOR2X1_193 ( .A(_3221_), .B(_3206_), .Y(_3228_) );
AOI21X1 AOI21X1_47 ( .A(bundleAddress_i[36]), .B(_3228_), .C(bundleAddress_i[35]), .Y(_3229_) );
NAND2X1 NAND2X1_604 ( .A(bundleAddress_i[36]), .B(bundleAddress_i[35]), .Y(_3230_) );
INVX1 INVX1_206 ( .A(_3221_), .Y(_3231_) );
NAND2X1 NAND2X1_605 ( .A(_3231_), .B(_3216_), .Y(_3232_) );
OAI21X1 OAI21X1_1286 ( .A(_3232_), .B(_3230_), .C(_612__bF_buf3), .Y(_3233_) );
OAI21X1 OAI21X1_1287 ( .A(_3229_), .B(_3233_), .C(_3227_), .Y(_898_) );
OAI21X1 OAI21X1_1288 ( .A(_1100__bF_buf14_bF_buf3), .B(_1031__bF_buf71), .C(_3638__34_), .Y(_3234_) );
NOR2X1 NOR2X1_194 ( .A(_3230_), .B(_3232_), .Y(_3235_) );
NOR2X1 NOR2X1_195 ( .A(bundleAddress_i[34]), .B(_3235_), .Y(_3236_) );
INVX1 INVX1_207 ( .A(_3230_), .Y(_3237_) );
NAND2X1 NAND2X1_606 ( .A(_3237_), .B(_3228_), .Y(_3238_) );
OAI21X1 OAI21X1_1289 ( .A(_3238_), .B(_2747_), .C(_612__bF_buf3), .Y(_3239_) );
OAI21X1 OAI21X1_1290 ( .A(_3239_), .B(_3236_), .C(_3234_), .Y(_899_) );
OAI21X1 OAI21X1_1291 ( .A(_1100__bF_buf13_bF_buf2), .B(_1031__bF_buf70), .C(_3638__33_), .Y(_3240_) );
AOI21X1 AOI21X1_48 ( .A(bundleAddress_i[34]), .B(_3235_), .C(bundleAddress_i[33]), .Y(_3241_) );
AND2X2 AND2X2_28 ( .A(_2976_), .B(_3237_), .Y(_3242_) );
AND2X2 AND2X2_29 ( .A(_3224_), .B(_3242_), .Y(_3243_) );
OR2X2 OR2X2_20 ( .A(_3243_), .B(_1101__bF_buf13), .Y(_3244_) );
OAI21X1 OAI21X1_1292 ( .A(_3241_), .B(_3244_), .C(_3240_), .Y(_900_) );
XNOR2X1 XNOR2X1_81 ( .A(_3243_), .B(bundleAddress_i[32]), .Y(_3245_) );
OAI21X1 OAI21X1_1293 ( .A(_1100__bF_buf12_bF_buf1), .B(_1031__bF_buf49), .C(_3638__32_), .Y(_3246_) );
OAI21X1 OAI21X1_1294 ( .A(_3245_), .B(_1101__bF_buf51), .C(_3246_), .Y(_901_) );
OAI21X1 OAI21X1_1295 ( .A(_1100__bF_buf11_bF_buf1), .B(_1031__bF_buf7), .C(_3638__31_), .Y(_3247_) );
AOI21X1 AOI21X1_49 ( .A(bundleAddress_i[32]), .B(_3243_), .C(bundleAddress_i[31]), .Y(_3248_) );
NAND3X1 NAND3X1_55 ( .A(_2968_), .B(_3242_), .C(_3224_), .Y(_3249_) );
NAND2X1 NAND2X1_607 ( .A(_612__bF_buf0), .B(_3249_), .Y(_3250_) );
OAI21X1 OAI21X1_1296 ( .A(_3248_), .B(_3250_), .C(_3247_), .Y(_902_) );
AND2X2 AND2X2_30 ( .A(_3249_), .B(_2755_), .Y(_3251_) );
OAI21X1 OAI21X1_1297 ( .A(_1100__bF_buf10_bF_buf1), .B(_1031__bF_buf44), .C(_3638__30_), .Y(_3252_) );
OAI21X1 OAI21X1_1298 ( .A(_3249_), .B(_2755_), .C(_612__bF_buf3), .Y(_3253_) );
OAI21X1 OAI21X1_1299 ( .A(_3251_), .B(_3253_), .C(_3252_), .Y(_903_) );
NOR2X1 NOR2X1_196 ( .A(_2757_), .B(_2973_), .Y(_3254_) );
NAND3X1 NAND3X1_56 ( .A(_3242_), .B(_3254_), .C(_3222_), .Y(_3255_) );
OAI21X1 OAI21X1_1300 ( .A(_3249_), .B(_2755_), .C(_2757_), .Y(_3256_) );
OAI21X1 OAI21X1_1301 ( .A(_3186_), .B(_3255_), .C(_3256_), .Y(_3257_) );
OAI21X1 OAI21X1_1302 ( .A(_1100__bF_buf9_bF_buf1), .B(_1031__bF_buf7), .C(_3638__29_), .Y(_3258_) );
OAI21X1 OAI21X1_1303 ( .A(_3257_), .B(_1101__bF_buf9), .C(_3258_), .Y(_904_) );
NOR2X1 NOR2X1_197 ( .A(_3255_), .B(_3186_), .Y(_3259_) );
XNOR2X1 XNOR2X1_82 ( .A(_3259_), .B(bundleAddress_i[28]), .Y(_3260_) );
OAI21X1 OAI21X1_1304 ( .A(_1100__bF_buf8_bF_buf2), .B(_1031__bF_buf38), .C(_3638__28_), .Y(_3261_) );
OAI21X1 OAI21X1_1305 ( .A(_3260_), .B(_1101__bF_buf27), .C(_3261_), .Y(_905_) );
INVX2 INVX2_106 ( .A(_3259_), .Y(_3262_) );
OAI21X1 OAI21X1_1306 ( .A(_3262_), .B(_2759_), .C(_2761_), .Y(_3263_) );
OAI21X1 OAI21X1_1307 ( .A(_2993_), .B(_3262_), .C(_3263_), .Y(_3264_) );
OAI21X1 OAI21X1_1308 ( .A(_1100__bF_buf7_bF_buf0), .B(_1031__bF_buf18), .C(_3638__27_), .Y(_3265_) );
OAI21X1 OAI21X1_1309 ( .A(_3264_), .B(_1101__bF_buf10), .C(_3265_), .Y(_906_) );
INVX1 INVX1_208 ( .A(_2993_), .Y(_3266_) );
NAND2X1 NAND2X1_608 ( .A(_3266_), .B(_3259_), .Y(_3267_) );
XNOR2X1 XNOR2X1_83 ( .A(_3267_), .B(_2763_), .Y(_3268_) );
OAI21X1 OAI21X1_1310 ( .A(_1100__bF_buf1), .B(_1031__bF_buf18), .C(_3638__26_), .Y(_3269_) );
OAI21X1 OAI21X1_1311 ( .A(_3268_), .B(_1101__bF_buf22), .C(_3269_), .Y(_907_) );
OAI21X1 OAI21X1_1312 ( .A(_1100__bF_buf1), .B(_1031__bF_buf18), .C(_3638__25_), .Y(_3270_) );
NOR2X1 NOR2X1_198 ( .A(_2763_), .B(_3267_), .Y(_3271_) );
NOR2X1 NOR2X1_199 ( .A(bundleAddress_i[25]), .B(_3271_), .Y(_3272_) );
NAND2X1 NAND2X1_609 ( .A(bundleAddress_i[26]), .B(bundleAddress_i[25]), .Y(_3273_) );
NOR2X1 NOR2X1_200 ( .A(_2993_), .B(_3273_), .Y(_3274_) );
NAND2X1 NAND2X1_610 ( .A(_3274_), .B(_3259_), .Y(_3275_) );
NAND2X1 NAND2X1_611 ( .A(_612__bF_buf3), .B(_3275_), .Y(_3276_) );
OAI21X1 OAI21X1_1313 ( .A(_3272_), .B(_3276_), .C(_3270_), .Y(_908_) );
XNOR2X1 XNOR2X1_84 ( .A(_3275_), .B(_2767_), .Y(_3277_) );
OAI21X1 OAI21X1_1314 ( .A(_1100__bF_buf1), .B(_1031__bF_buf18), .C(_3638__24_), .Y(_3278_) );
OAI21X1 OAI21X1_1315 ( .A(_3277_), .B(_1101__bF_buf10), .C(_3278_), .Y(_909_) );
OAI21X1 OAI21X1_1316 ( .A(_1100__bF_buf1), .B(_1031__bF_buf38), .C(_3638__23_), .Y(_3279_) );
OAI21X1 OAI21X1_1317 ( .A(_3275_), .B(_2767_), .C(_2769_), .Y(_3280_) );
OAI21X1 OAI21X1_1318 ( .A(_3005_), .B(_3275_), .C(_3280_), .Y(_3281_) );
OAI21X1 OAI21X1_1319 ( .A(_3281_), .B(_1101__bF_buf27), .C(_3279_), .Y(_910_) );
OAI21X1 OAI21X1_1320 ( .A(_1100__bF_buf1), .B(_1031__bF_buf38), .C(_3638__22_), .Y(_3282_) );
AND2X2 AND2X2_31 ( .A(_3259_), .B(_3274_), .Y(_3283_) );
AOI21X1 AOI21X1_50 ( .A(_3013_), .B(_3283_), .C(bundleAddress_i[22]), .Y(_3284_) );
NAND2X1 NAND2X1_612 ( .A(_3013_), .B(_3283_), .Y(_3285_) );
OAI21X1 OAI21X1_1321 ( .A(_3285_), .B(_2771_), .C(_612__bF_buf2), .Y(_3286_) );
OAI21X1 OAI21X1_1322 ( .A(_3286_), .B(_3284_), .C(_3282_), .Y(_911_) );
INVX1 INVX1_209 ( .A(_3638__21_), .Y(_3287_) );
NOR3X1 NOR3X1_16 ( .A(_2771_), .B(_3005_), .C(_3275_), .Y(_3288_) );
NAND2X1 NAND2X1_613 ( .A(bundleAddress_i[22]), .B(bundleAddress_i[21]), .Y(_3289_) );
NOR2X1 NOR2X1_201 ( .A(_3005_), .B(_3289_), .Y(_3290_) );
NAND2X1 NAND2X1_614 ( .A(_3274_), .B(_3290_), .Y(_3291_) );
NOR3X1 NOR3X1_17 ( .A(_3255_), .B(_3291_), .C(_3186_), .Y(_3292_) );
NOR2X1 NOR2X1_202 ( .A(_1101__bF_buf19), .B(_3292_), .Y(_3293_) );
OAI21X1 OAI21X1_1323 ( .A(_3288_), .B(bundleAddress_i[21]), .C(_3293_), .Y(_3294_) );
OAI21X1 OAI21X1_1324 ( .A(_3287_), .B(_612__bF_buf2), .C(_3294_), .Y(_912_) );
NAND2X1 NAND2X1_615 ( .A(bundleAddress_i[20]), .B(_3292_), .Y(_3295_) );
OAI21X1 OAI21X1_1325 ( .A(_3262_), .B(_3291_), .C(_2775_), .Y(_3296_) );
NAND2X1 NAND2X1_616 ( .A(_3295_), .B(_3296_), .Y(_3297_) );
OAI21X1 OAI21X1_1326 ( .A(_1100__bF_buf1), .B(_1031__bF_buf44), .C(_3638__20_), .Y(_3298_) );
OAI21X1 OAI21X1_1327 ( .A(_3297_), .B(_1101__bF_buf19), .C(_3298_), .Y(_913_) );
OAI21X1 OAI21X1_1328 ( .A(_1100__bF_buf1), .B(_1031__bF_buf44), .C(_3638__19_), .Y(_3299_) );
AOI21X1 AOI21X1_51 ( .A(bundleAddress_i[20]), .B(_3292_), .C(bundleAddress_i[19]), .Y(_3300_) );
INVX1 INVX1_210 ( .A(_3255_), .Y(_3301_) );
INVX2 INVX2_107 ( .A(_3291_), .Y(_3302_) );
NAND3X1 NAND3X1_57 ( .A(_3302_), .B(_3205_), .C(_3301_), .Y(_3303_) );
OAI21X1 OAI21X1_1329 ( .A(_3303_), .B(_3024_), .C(_612__bF_buf0), .Y(_3304_) );
OAI21X1 OAI21X1_1330 ( .A(_3304_), .B(_3300_), .C(_3299_), .Y(_914_) );
OAI21X1 OAI21X1_1331 ( .A(_1100__bF_buf14_bF_buf3), .B(_1031__bF_buf64), .C(_3638__18_), .Y(_3305_) );
NOR2X1 NOR2X1_203 ( .A(_3024_), .B(_3303_), .Y(_3306_) );
XNOR2X1 XNOR2X1_85 ( .A(_3306_), .B(bundleAddress_i[18]), .Y(_3307_) );
OAI21X1 OAI21X1_1332 ( .A(_3307_), .B(_1101__bF_buf22), .C(_3305_), .Y(_915_) );
OAI21X1 OAI21X1_1333 ( .A(_1100__bF_buf13_bF_buf3), .B(_1031__bF_buf28), .C(_3638__17_), .Y(_3308_) );
AOI21X1 AOI21X1_52 ( .A(bundleAddress_i[18]), .B(_3306_), .C(bundleAddress_i[17]), .Y(_3309_) );
NAND2X1 NAND2X1_617 ( .A(bundleAddress_i[18]), .B(bundleAddress_i[17]), .Y(_3310_) );
NOR2X1 NOR2X1_204 ( .A(_3024_), .B(_3310_), .Y(_3311_) );
INVX1 INVX1_211 ( .A(_3311_), .Y(_3312_) );
OAI21X1 OAI21X1_1334 ( .A(_3303_), .B(_3312_), .C(_612__bF_buf0), .Y(_3313_) );
OAI21X1 OAI21X1_1335 ( .A(_3309_), .B(_3313_), .C(_3308_), .Y(_916_) );
OAI21X1 OAI21X1_1336 ( .A(_1100__bF_buf12_bF_buf1), .B(_1031__bF_buf49), .C(_3638__16_), .Y(_3314_) );
NAND2X1 NAND2X1_618 ( .A(_3311_), .B(_3292_), .Y(_3315_) );
INVX1 INVX1_212 ( .A(_3315_), .Y(_3316_) );
NOR2X1 NOR2X1_205 ( .A(bundleAddress_i[16]), .B(_3316_), .Y(_3317_) );
OAI21X1 OAI21X1_1337 ( .A(_3315_), .B(_2783_), .C(_612__bF_buf0), .Y(_3318_) );
OAI21X1 OAI21X1_1338 ( .A(_3317_), .B(_3318_), .C(_3314_), .Y(_917_) );
OAI21X1 OAI21X1_1339 ( .A(_1100__bF_buf11_bF_buf1), .B(_1031__bF_buf46), .C(_3638__15_), .Y(_3319_) );
AOI21X1 AOI21X1_53 ( .A(bundleAddress_i[16]), .B(_3316_), .C(bundleAddress_i[15]), .Y(_3320_) );
OAI21X1 OAI21X1_1340 ( .A(_3315_), .B(_3044_), .C(_612__bF_buf0), .Y(_3321_) );
OAI21X1 OAI21X1_1341 ( .A(_3320_), .B(_3321_), .C(_3319_), .Y(_918_) );
NAND3X1 NAND3X1_58 ( .A(_3047_), .B(_3311_), .C(_3292_), .Y(_3322_) );
INVX1 INVX1_213 ( .A(_3322_), .Y(_3323_) );
NOR2X1 NOR2X1_206 ( .A(bundleAddress_i[14]), .B(_3323_), .Y(_3324_) );
OAI21X1 OAI21X1_1342 ( .A(_1100__bF_buf10_bF_buf0), .B(_1031__bF_buf46), .C(_3638__14_), .Y(_3325_) );
OAI21X1 OAI21X1_1343 ( .A(_3322_), .B(_2787_), .C(_612__bF_buf0), .Y(_3326_) );
OAI21X1 OAI21X1_1344 ( .A(_3324_), .B(_3326_), .C(_3325_), .Y(_919_) );
OAI21X1 OAI21X1_1345 ( .A(_1100__bF_buf9_bF_buf0), .B(_1031__bF_buf46), .C(_3638__13_), .Y(_3327_) );
AOI21X1 AOI21X1_54 ( .A(bundleAddress_i[14]), .B(_3323_), .C(bundleAddress_i[13]), .Y(_3328_) );
NAND2X1 NAND2X1_619 ( .A(bundleAddress_i[14]), .B(bundleAddress_i[13]), .Y(_3329_) );
NOR2X1 NOR2X1_207 ( .A(_3044_), .B(_3329_), .Y(_3330_) );
AND2X2 AND2X2_32 ( .A(_3311_), .B(_3330_), .Y(_3331_) );
NAND2X1 NAND2X1_620 ( .A(_3331_), .B(_3302_), .Y(_3332_) );
OAI21X1 OAI21X1_1346 ( .A(_3262_), .B(_3332_), .C(_612__bF_buf3), .Y(_3333_) );
OAI21X1 OAI21X1_1347 ( .A(_3328_), .B(_3333_), .C(_3327_), .Y(_920_) );
NOR3X1 NOR3X1_18 ( .A(_3255_), .B(_3332_), .C(_3186_), .Y(_3334_) );
XNOR2X1 XNOR2X1_86 ( .A(_3334_), .B(bundleAddress_i[12]), .Y(_3335_) );
OAI21X1 OAI21X1_1348 ( .A(_1100__bF_buf8_bF_buf2), .B(_1031__bF_buf57), .C(_3638__12_), .Y(_3336_) );
OAI21X1 OAI21X1_1349 ( .A(_3335_), .B(_1101__bF_buf35), .C(_3336_), .Y(_921_) );
OAI21X1 OAI21X1_1350 ( .A(_1100__bF_buf7_bF_buf3), .B(_1031__bF_buf31), .C(_3638__11_), .Y(_3337_) );
AOI21X1 AOI21X1_55 ( .A(bundleAddress_i[12]), .B(_3334_), .C(bundleAddress_i[11]), .Y(_3338_) );
AND2X2 AND2X2_33 ( .A(_3302_), .B(_3331_), .Y(_3339_) );
NAND3X1 NAND3X1_59 ( .A(_3339_), .B(_3205_), .C(_3301_), .Y(_3340_) );
OAI21X1 OAI21X1_1351 ( .A(_3340_), .B(_3065_), .C(_612__bF_buf2), .Y(_3341_) );
OAI21X1 OAI21X1_1352 ( .A(_3341_), .B(_3338_), .C(_3337_), .Y(_922_) );
OAI21X1 OAI21X1_1353 ( .A(_1100__bF_buf2), .B(_1031__bF_buf46), .C(_3638__10_), .Y(_3342_) );
NOR2X1 NOR2X1_208 ( .A(_3065_), .B(_3340_), .Y(_3343_) );
XNOR2X1 XNOR2X1_87 ( .A(_3343_), .B(bundleAddress_i[10]), .Y(_3344_) );
OAI21X1 OAI21X1_1354 ( .A(_3344_), .B(_1101__bF_buf58), .C(_3342_), .Y(_923_) );
OAI21X1 OAI21X1_1355 ( .A(_1100__bF_buf2), .B(_1031__bF_buf24), .C(_3638__9_), .Y(_3345_) );
AOI21X1 AOI21X1_56 ( .A(bundleAddress_i[10]), .B(_3343_), .C(bundleAddress_i[9]), .Y(_3346_) );
NAND2X1 NAND2X1_621 ( .A(_3064_), .B(_3094_), .Y(_3347_) );
OAI21X1 OAI21X1_1356 ( .A(_3340_), .B(_3347_), .C(_612__bF_buf2), .Y(_3348_) );
OAI21X1 OAI21X1_1357 ( .A(_3346_), .B(_3348_), .C(_3345_), .Y(_924_) );
OAI21X1 OAI21X1_1358 ( .A(_1100__bF_buf2), .B(_1031__bF_buf31), .C(_3638__8_), .Y(_3349_) );
INVX1 INVX1_214 ( .A(_3347_), .Y(_3350_) );
NAND2X1 NAND2X1_622 ( .A(_3350_), .B(_3334_), .Y(_3351_) );
INVX1 INVX1_215 ( .A(_3351_), .Y(_3352_) );
NOR2X1 NOR2X1_209 ( .A(bundleAddress_i[8]), .B(_3352_), .Y(_3353_) );
OAI21X1 OAI21X1_1359 ( .A(_3351_), .B(_2799_), .C(_612__bF_buf2), .Y(_3354_) );
OAI21X1 OAI21X1_1360 ( .A(_3353_), .B(_3354_), .C(_3349_), .Y(_925_) );
OAI21X1 OAI21X1_1361 ( .A(_1100__bF_buf2), .B(_1031__bF_buf14), .C(_3638__7_), .Y(_3355_) );
OAI21X1 OAI21X1_1362 ( .A(_3351_), .B(_2799_), .C(_2801_), .Y(_3356_) );
OAI21X1 OAI21X1_1363 ( .A(_3087_), .B(_3351_), .C(_3356_), .Y(_3357_) );
OAI21X1 OAI21X1_1364 ( .A(_3357_), .B(_1101__bF_buf58), .C(_3355_), .Y(_926_) );
OAI21X1 OAI21X1_1365 ( .A(_1100__bF_buf2), .B(_1031__bF_buf31), .C(_3638__6_), .Y(_3358_) );
AOI21X1 AOI21X1_57 ( .A(_3086_), .B(_3352_), .C(bundleAddress_i[6]), .Y(_3359_) );
OAI21X1 OAI21X1_1366 ( .A(_3351_), .B(_3092_), .C(_612__bF_buf2), .Y(_3360_) );
OAI21X1 OAI21X1_1367 ( .A(_3359_), .B(_3360_), .C(_3358_), .Y(_927_) );
NAND3X1 NAND3X1_60 ( .A(bundleAddress_i[5]), .B(_3064_), .C(_3094_), .Y(_3361_) );
NOR2X1 NOR2X1_210 ( .A(_3092_), .B(_3361_), .Y(_3362_) );
INVX1 INVX1_216 ( .A(_3362_), .Y(_3363_) );
OAI21X1 OAI21X1_1368 ( .A(_3351_), .B(_3092_), .C(_2805_), .Y(_3364_) );
OAI21X1 OAI21X1_1369 ( .A(_3340_), .B(_3363_), .C(_3364_), .Y(_3365_) );
OAI21X1 OAI21X1_1370 ( .A(_1100__bF_buf1), .B(_1031__bF_buf24), .C(_3638__5_), .Y(_3366_) );
OAI21X1 OAI21X1_1371 ( .A(_3365_), .B(_1101__bF_buf19), .C(_3366_), .Y(_928_) );
OAI21X1 OAI21X1_1372 ( .A(_1100__bF_buf2), .B(_1031__bF_buf58), .C(_3638__4_), .Y(_3367_) );
NOR2X1 NOR2X1_211 ( .A(_3363_), .B(_3340_), .Y(_3368_) );
XNOR2X1 XNOR2X1_88 ( .A(_3368_), .B(bundleAddress_i[4]), .Y(_3369_) );
OAI21X1 OAI21X1_1373 ( .A(_3369_), .B(_1101__bF_buf38), .C(_3367_), .Y(_929_) );
OAI21X1 OAI21X1_1374 ( .A(_1100__bF_buf14_bF_buf1), .B(_1031__bF_buf40), .C(_3638__3_), .Y(_3370_) );
AOI21X1 AOI21X1_58 ( .A(bundleAddress_i[4]), .B(_3368_), .C(bundleAddress_i[3]), .Y(_3371_) );
NAND3X1 NAND3X1_61 ( .A(_3109_), .B(_3362_), .C(_3334_), .Y(_3372_) );
NAND2X1 NAND2X1_623 ( .A(_612__bF_buf0), .B(_3372_), .Y(_3373_) );
OAI21X1 OAI21X1_1375 ( .A(_3371_), .B(_3373_), .C(_3370_), .Y(_930_) );
INVX1 INVX1_217 ( .A(_3372_), .Y(_3374_) );
NOR2X1 NOR2X1_212 ( .A(bundleAddress_i[2]), .B(_3374_), .Y(_3375_) );
OAI21X1 OAI21X1_1376 ( .A(_1100__bF_buf13_bF_buf3), .B(_1031__bF_buf31), .C(_3638__2_), .Y(_3376_) );
OAI21X1 OAI21X1_1377 ( .A(_3372_), .B(_2811_), .C(_612__bF_buf2), .Y(_3377_) );
OAI21X1 OAI21X1_1378 ( .A(_3375_), .B(_3377_), .C(_3376_), .Y(_931_) );
OAI21X1 OAI21X1_1379 ( .A(_1100__bF_buf12_bF_buf1), .B(_1031__bF_buf28), .C(_3638__1_), .Y(_3378_) );
AOI21X1 AOI21X1_59 ( .A(bundleAddress_i[2]), .B(_3374_), .C(bundleAddress_i[1]), .Y(_3379_) );
NOR2X1 NOR2X1_213 ( .A(_2811_), .B(_2813_), .Y(_3380_) );
INVX1 INVX1_218 ( .A(_3380_), .Y(_3381_) );
OAI21X1 OAI21X1_1380 ( .A(_3372_), .B(_3381_), .C(_612__bF_buf0), .Y(_3382_) );
OAI21X1 OAI21X1_1381 ( .A(_3379_), .B(_3382_), .C(_3378_), .Y(_932_) );
NOR2X1 NOR2X1_214 ( .A(_3110_), .B(_3381_), .Y(_3383_) );
NAND3X1 NAND3X1_62 ( .A(_3362_), .B(_3383_), .C(_3334_), .Y(_3384_) );
XNOR2X1 XNOR2X1_89 ( .A(_3384_), .B(_2815_), .Y(_3385_) );
OAI21X1 OAI21X1_1382 ( .A(_1100__bF_buf11_bF_buf1), .B(_1031__bF_buf28), .C(_3638__0_), .Y(_3386_) );
OAI21X1 OAI21X1_1383 ( .A(_3385_), .B(_1101__bF_buf17), .C(_3386_), .Y(_933_) );
OAI21X1 OAI21X1_1384 ( .A(_1101__bF_buf1), .B(_1135__bF_buf6_bF_buf0), .C(_3639__63_), .Y(_3387_) );
OAI21X1 OAI21X1_1385 ( .A(_2689_), .B(_1134__bF_buf2), .C(_3387_), .Y(_934_) );
OAI21X1 OAI21X1_1386 ( .A(_1101__bF_buf54), .B(_1135__bF_buf5_bF_buf0), .C(_3639__62_), .Y(_3388_) );
OAI21X1 OAI21X1_1387 ( .A(_2691_), .B(_1134__bF_buf7), .C(_3388_), .Y(_935_) );
OAI21X1 OAI21X1_1388 ( .A(_1101__bF_buf0), .B(_1135__bF_buf4_bF_buf0), .C(_3639__61_), .Y(_3389_) );
OAI21X1 OAI21X1_1389 ( .A(bundleAddress_i[61]), .B(_1134__bF_buf13), .C(_3389_), .Y(_936_) );
OAI21X1 OAI21X1_1390 ( .A(_1101__bF_buf11), .B(_1135__bF_buf3_bF_buf2), .C(_3639__60_), .Y(_3390_) );
OAI21X1 OAI21X1_1391 ( .A(_2823_), .B(_1134__bF_buf12), .C(_3390_), .Y(_937_) );
OAI21X1 OAI21X1_1392 ( .A(bundleAddress_i[61]), .B(bundleAddress_i[60]), .C(bundleAddress_i[59]), .Y(_3391_) );
OAI21X1 OAI21X1_1393 ( .A(_3129_), .B(bundleAddress_i[61]), .C(_3391_), .Y(_3392_) );
OAI21X1 OAI21X1_1394 ( .A(_1101__bF_buf34), .B(_1135__bF_buf2_bF_buf1), .C(_3639__59_), .Y(_3393_) );
OAI21X1 OAI21X1_1395 ( .A(_3392_), .B(_1134__bF_buf4), .C(_3393_), .Y(_938_) );
OAI21X1 OAI21X1_1396 ( .A(_2822_), .B(_2697_), .C(_2699_), .Y(_3394_) );
OAI21X1 OAI21X1_1397 ( .A(_2822_), .B(_2832_), .C(_3394_), .Y(_3395_) );
OAI21X1 OAI21X1_1398 ( .A(_1101__bF_buf53), .B(_1135__bF_buf1_bF_buf1), .C(_3639__58_), .Y(_3396_) );
OAI21X1 OAI21X1_1399 ( .A(_3395_), .B(_1134__bF_buf13), .C(_3396_), .Y(_939_) );
NOR2X1 NOR2X1_215 ( .A(_2832_), .B(_2822_), .Y(_3397_) );
XNOR2X1 XNOR2X1_90 ( .A(_3397_), .B(bundleAddress_i[57]), .Y(_3398_) );
OAI21X1 OAI21X1_1400 ( .A(_1101__bF_buf28), .B(_1135__bF_buf14), .C(_3639__57_), .Y(_3399_) );
OAI21X1 OAI21X1_1401 ( .A(_3398_), .B(_1134__bF_buf13), .C(_3399_), .Y(_940_) );
INVX4 INVX4_50 ( .A(_3397_), .Y(_3400_) );
OAI21X1 OAI21X1_1402 ( .A(_3400_), .B(_2701_), .C(_2703_), .Y(_3401_) );
OAI21X1 OAI21X1_1403 ( .A(_2844_), .B(_3400_), .C(_3401_), .Y(_3402_) );
OAI21X1 OAI21X1_1404 ( .A(_1101__bF_buf33), .B(_1135__bF_buf14_bF_buf0), .C(_3639__56_), .Y(_3403_) );
OAI21X1 OAI21X1_1405 ( .A(_3402_), .B(_1134__bF_buf13), .C(_3403_), .Y(_941_) );
NOR2X1 NOR2X1_216 ( .A(_2844_), .B(_3400_), .Y(_3404_) );
INVX1 INVX1_219 ( .A(_3404_), .Y(_3405_) );
NOR2X1 NOR2X1_217 ( .A(_2705_), .B(_3405_), .Y(_3406_) );
OAI21X1 OAI21X1_1406 ( .A(_3404_), .B(bundleAddress_i[55]), .C(_613__bF_buf3), .Y(_3407_) );
OAI21X1 OAI21X1_1407 ( .A(_1101__bF_buf0), .B(_1135__bF_buf13_bF_buf3), .C(_3639__55_), .Y(_3408_) );
OAI21X1 OAI21X1_1408 ( .A(_3406_), .B(_3407_), .C(_3408_), .Y(_942_) );
OAI21X1 OAI21X1_1409 ( .A(_3405_), .B(_2705_), .C(_2707_), .Y(_3409_) );
OAI21X1 OAI21X1_1410 ( .A(_2857_), .B(_3400_), .C(_3409_), .Y(_3410_) );
OAI21X1 OAI21X1_1411 ( .A(_1101__bF_buf34), .B(_1135__bF_buf12_bF_buf2), .C(_3639__54_), .Y(_3411_) );
OAI21X1 OAI21X1_1412 ( .A(_3410_), .B(_1134__bF_buf13), .C(_3411_), .Y(_943_) );
NAND2X1 NAND2X1_624 ( .A(_2856_), .B(_3397_), .Y(_3412_) );
NOR2X1 NOR2X1_218 ( .A(_2709_), .B(_3412_), .Y(_3413_) );
INVX2 INVX2_108 ( .A(_3413_), .Y(_3414_) );
OAI21X1 OAI21X1_1413 ( .A(_3400_), .B(_2857_), .C(_2709_), .Y(_3415_) );
NAND2X1 NAND2X1_625 ( .A(_3415_), .B(_3414_), .Y(_3416_) );
OAI21X1 OAI21X1_1414 ( .A(_1101__bF_buf33), .B(_1135__bF_buf11_bF_buf0), .C(_3639__53_), .Y(_3417_) );
OAI21X1 OAI21X1_1415 ( .A(_3416_), .B(_1134__bF_buf14), .C(_3417_), .Y(_944_) );
XNOR2X1 XNOR2X1_91 ( .A(_3413_), .B(bundleAddress_i[52]), .Y(_3418_) );
OAI21X1 OAI21X1_1416 ( .A(_1101__bF_buf8), .B(_1135__bF_buf10_bF_buf2), .C(_3639__52_), .Y(_3419_) );
OAI21X1 OAI21X1_1417 ( .A(_3418_), .B(_1134__bF_buf14), .C(_3419_), .Y(_945_) );
AOI21X1 AOI21X1_60 ( .A(bundleAddress_i[52]), .B(_3413_), .C(bundleAddress_i[51]), .Y(_3420_) );
OAI21X1 OAI21X1_1418 ( .A(_3414_), .B(_2869_), .C(_613__bF_buf0), .Y(_3421_) );
OAI21X1 OAI21X1_1419 ( .A(_1101__bF_buf23), .B(_1135__bF_buf9_bF_buf0), .C(_3639__51_), .Y(_3422_) );
OAI21X1 OAI21X1_1420 ( .A(_3421_), .B(_3420_), .C(_3422_), .Y(_946_) );
OAI21X1 OAI21X1_1421 ( .A(_3414_), .B(_2869_), .C(_2715_), .Y(_3423_) );
OAI21X1 OAI21X1_1422 ( .A(_3157_), .B(_3414_), .C(_3423_), .Y(_3424_) );
OAI21X1 OAI21X1_1423 ( .A(_1101__bF_buf33), .B(_1135__bF_buf8_bF_buf1), .C(_3639__50_), .Y(_3425_) );
OAI21X1 OAI21X1_1424 ( .A(_3424_), .B(_1134__bF_buf14), .C(_3425_), .Y(_947_) );
NAND3X1 NAND3X1_63 ( .A(bundleAddress_i[50]), .B(_2878_), .C(_3413_), .Y(_3426_) );
NOR2X1 NOR2X1_219 ( .A(_2717_), .B(_3426_), .Y(_3427_) );
INVX1 INVX1_220 ( .A(_3426_), .Y(_3428_) );
OAI21X1 OAI21X1_1425 ( .A(_3428_), .B(bundleAddress_i[49]), .C(_613__bF_buf0), .Y(_3429_) );
OAI21X1 OAI21X1_1426 ( .A(_1101__bF_buf8), .B(_1135__bF_buf7_bF_buf2), .C(_3639__49_), .Y(_3430_) );
OAI21X1 OAI21X1_1427 ( .A(_3429_), .B(_3427_), .C(_3430_), .Y(_948_) );
XNOR2X1 XNOR2X1_92 ( .A(_3427_), .B(bundleAddress_i[48]), .Y(_3431_) );
OAI21X1 OAI21X1_1428 ( .A(_1101__bF_buf8), .B(_1135__bF_buf6_bF_buf2), .C(_3639__48_), .Y(_3432_) );
OAI21X1 OAI21X1_1429 ( .A(_3431_), .B(_1134__bF_buf12), .C(_3432_), .Y(_949_) );
INVX1 INVX1_221 ( .A(_3427_), .Y(_3433_) );
OAI21X1 OAI21X1_1430 ( .A(_3433_), .B(_2719_), .C(_2721_), .Y(_3434_) );
OAI21X1 OAI21X1_1431 ( .A(_3168_), .B(_3433_), .C(_3434_), .Y(_3435_) );
OAI21X1 OAI21X1_1432 ( .A(_1101__bF_buf52), .B(_1135__bF_buf5_bF_buf2), .C(_3639__47_), .Y(_3436_) );
OAI21X1 OAI21X1_1433 ( .A(_3435_), .B(_1134__bF_buf12), .C(_3436_), .Y(_950_) );
NAND2X1 NAND2X1_626 ( .A(_3167_), .B(_3427_), .Y(_3437_) );
XNOR2X1 XNOR2X1_93 ( .A(_3437_), .B(_2723_), .Y(_3438_) );
OAI21X1 OAI21X1_1434 ( .A(_1101__bF_buf52), .B(_1135__bF_buf4_bF_buf1), .C(_3639__46_), .Y(_3439_) );
OAI21X1 OAI21X1_1435 ( .A(_3438_), .B(_1134__bF_buf12), .C(_3439_), .Y(_951_) );
NOR2X1 NOR2X1_220 ( .A(_2897_), .B(_3412_), .Y(_3440_) );
NAND2X1 NAND2X1_627 ( .A(bundleAddress_i[45]), .B(_3440_), .Y(_3441_) );
OAI21X1 OAI21X1_1436 ( .A(_3412_), .B(_2897_), .C(_2725_), .Y(_3442_) );
NAND2X1 NAND2X1_628 ( .A(_3442_), .B(_3441_), .Y(_3443_) );
OAI21X1 OAI21X1_1437 ( .A(_1101__bF_buf11), .B(_1135__bF_buf3_bF_buf2), .C(_3639__45_), .Y(_3444_) );
OAI21X1 OAI21X1_1438 ( .A(_3443_), .B(_1134__bF_buf12), .C(_3444_), .Y(_952_) );
INVX4 INVX4_51 ( .A(_3440_), .Y(_3445_) );
OAI21X1 OAI21X1_1439 ( .A(_3445_), .B(_2725_), .C(_2727_), .Y(_3446_) );
OAI21X1 OAI21X1_1440 ( .A(_2909_), .B(_3445_), .C(_3446_), .Y(_3447_) );
OAI21X1 OAI21X1_1441 ( .A(_1101__bF_buf5), .B(_1135__bF_buf2_bF_buf3), .C(_3639__44_), .Y(_3448_) );
OAI21X1 OAI21X1_1442 ( .A(_3447_), .B(_1134__bF_buf5), .C(_3448_), .Y(_953_) );
NOR2X1 NOR2X1_221 ( .A(_2909_), .B(_3445_), .Y(_3449_) );
NAND2X1 NAND2X1_629 ( .A(bundleAddress_i[43]), .B(_3449_), .Y(_3450_) );
INVX1 INVX1_222 ( .A(_3450_), .Y(_3451_) );
OAI21X1 OAI21X1_1443 ( .A(_3449_), .B(bundleAddress_i[43]), .C(_613__bF_buf2), .Y(_3452_) );
OAI21X1 OAI21X1_1444 ( .A(_1101__bF_buf55), .B(_1135__bF_buf1_bF_buf3), .C(_3639__43_), .Y(_3453_) );
OAI21X1 OAI21X1_1445 ( .A(_3451_), .B(_3452_), .C(_3453_), .Y(_954_) );
XNOR2X1 XNOR2X1_94 ( .A(_3450_), .B(_2731_), .Y(_3454_) );
OAI21X1 OAI21X1_1446 ( .A(_1101__bF_buf10), .B(_1135__bF_buf3), .C(_3639__42_), .Y(_3455_) );
OAI21X1 OAI21X1_1447 ( .A(_3454_), .B(_1134__bF_buf5), .C(_3455_), .Y(_955_) );
OAI21X1 OAI21X1_1448 ( .A(_3450_), .B(_2731_), .C(_2733_), .Y(_3456_) );
OAI21X1 OAI21X1_1449 ( .A(_2919_), .B(_3441_), .C(_3456_), .Y(_3457_) );
OAI21X1 OAI21X1_1450 ( .A(_1101__bF_buf50), .B(_1135__bF_buf14_bF_buf2), .C(_3639__41_), .Y(_3458_) );
OAI21X1 OAI21X1_1451 ( .A(_3457_), .B(_1134__bF_buf5), .C(_3458_), .Y(_956_) );
NOR2X1 NOR2X1_222 ( .A(_2919_), .B(_3441_), .Y(_3459_) );
XNOR2X1 XNOR2X1_95 ( .A(_3459_), .B(bundleAddress_i[40]), .Y(_3460_) );
OAI21X1 OAI21X1_1452 ( .A(_1101__bF_buf10), .B(_1135__bF_buf13_bF_buf0), .C(_3639__40_), .Y(_3461_) );
OAI21X1 OAI21X1_1453 ( .A(_3460_), .B(_1134__bF_buf5), .C(_3461_), .Y(_957_) );
OAI21X1 OAI21X1_1454 ( .A(_1101__bF_buf5), .B(_1135__bF_buf12_bF_buf3), .C(_3639__39_), .Y(_3462_) );
NAND2X1 NAND2X1_630 ( .A(_2926_), .B(_3440_), .Y(_3463_) );
NOR2X1 NOR2X1_223 ( .A(_2928_), .B(_3463_), .Y(_3464_) );
XNOR2X1 XNOR2X1_96 ( .A(_3464_), .B(bundleAddress_i[39]), .Y(_3465_) );
OAI21X1 OAI21X1_1455 ( .A(_3465_), .B(_1134__bF_buf5), .C(_3462_), .Y(_958_) );
NAND2X1 NAND2X1_631 ( .A(bundleAddress_i[39]), .B(_3464_), .Y(_3466_) );
XNOR2X1 XNOR2X1_97 ( .A(_3466_), .B(_2739_), .Y(_3467_) );
OAI21X1 OAI21X1_1456 ( .A(_1101__bF_buf20), .B(_1135__bF_buf11_bF_buf3), .C(_3639__38_), .Y(_3468_) );
OAI21X1 OAI21X1_1457 ( .A(_3467_), .B(_1134__bF_buf11), .C(_3468_), .Y(_959_) );
NOR2X1 NOR2X1_224 ( .A(_2937_), .B(_3445_), .Y(_3469_) );
NAND2X1 NAND2X1_632 ( .A(bundleAddress_i[37]), .B(_3469_), .Y(_3470_) );
OAI21X1 OAI21X1_1458 ( .A(_3445_), .B(_2937_), .C(_2741_), .Y(_3471_) );
NAND2X1 NAND2X1_633 ( .A(_3471_), .B(_3470_), .Y(_3472_) );
OAI21X1 OAI21X1_1459 ( .A(_1101__bF_buf20), .B(_1135__bF_buf10_bF_buf1), .C(_3639__37_), .Y(_3473_) );
OAI21X1 OAI21X1_1460 ( .A(_3472_), .B(_1134__bF_buf11), .C(_3473_), .Y(_960_) );
XNOR2X1 XNOR2X1_98 ( .A(_3470_), .B(_2743_), .Y(_3474_) );
OAI21X1 OAI21X1_1461 ( .A(_1101__bF_buf13), .B(_1135__bF_buf9_bF_buf3), .C(_3639__36_), .Y(_3475_) );
OAI21X1 OAI21X1_1462 ( .A(_3474_), .B(_1134__bF_buf11), .C(_3475_), .Y(_961_) );
INVX2 INVX2_109 ( .A(_3469_), .Y(_3476_) );
OAI21X1 OAI21X1_1463 ( .A(_3470_), .B(_2743_), .C(_2745_), .Y(_3477_) );
OAI21X1 OAI21X1_1464 ( .A(_2953_), .B(_3476_), .C(_3477_), .Y(_3478_) );
OAI21X1 OAI21X1_1465 ( .A(_1101__bF_buf41), .B(_1135__bF_buf8_bF_buf3), .C(_3639__35_), .Y(_3479_) );
OAI21X1 OAI21X1_1466 ( .A(_3478_), .B(_1134__bF_buf11), .C(_3479_), .Y(_962_) );
OAI21X1 OAI21X1_1467 ( .A(_3476_), .B(_2953_), .C(_2747_), .Y(_3480_) );
OAI21X1 OAI21X1_1468 ( .A(_2955_), .B(_3476_), .C(_3480_), .Y(_3481_) );
OAI21X1 OAI21X1_1469 ( .A(_1101__bF_buf22), .B(_1135__bF_buf7_bF_buf1), .C(_3639__34_), .Y(_3482_) );
OAI21X1 OAI21X1_1470 ( .A(_3481_), .B(_1134__bF_buf9), .C(_3482_), .Y(_963_) );
OAI21X1 OAI21X1_1471 ( .A(_3476_), .B(_2955_), .C(_2749_), .Y(_3483_) );
NAND3X1 NAND3X1_64 ( .A(_2954_), .B(_2976_), .C(_3469_), .Y(_3484_) );
NAND2X1 NAND2X1_634 ( .A(_3484_), .B(_3483_), .Y(_3485_) );
OAI21X1 OAI21X1_1472 ( .A(_1101__bF_buf13), .B(_1135__bF_buf6_bF_buf0), .C(_3639__33_), .Y(_3486_) );
OAI21X1 OAI21X1_1473 ( .A(_3485_), .B(_1134__bF_buf11), .C(_3486_), .Y(_964_) );
XNOR2X1 XNOR2X1_99 ( .A(_3484_), .B(_2751_), .Y(_3487_) );
OAI21X1 OAI21X1_1474 ( .A(_1101__bF_buf51), .B(_1135__bF_buf5_bF_buf1), .C(_3639__32_), .Y(_3488_) );
OAI21X1 OAI21X1_1475 ( .A(_3487_), .B(_1134__bF_buf2), .C(_3488_), .Y(_965_) );
OAI21X1 OAI21X1_1476 ( .A(_3484_), .B(_2751_), .C(_2753_), .Y(_3489_) );
OAI21X1 OAI21X1_1477 ( .A(_2969_), .B(_3484_), .C(_3489_), .Y(_3490_) );
OAI21X1 OAI21X1_1478 ( .A(_1101__bF_buf9), .B(_1135__bF_buf4_bF_buf3), .C(_3639__31_), .Y(_3491_) );
OAI21X1 OAI21X1_1479 ( .A(_3490_), .B(_1134__bF_buf2), .C(_3491_), .Y(_966_) );
OAI21X1 OAI21X1_1480 ( .A(_1101__bF_buf9), .B(_1135__bF_buf3_bF_buf3), .C(_3639__30_), .Y(_3492_) );
NAND2X1 NAND2X1_635 ( .A(_3440_), .B(_2978_), .Y(_3493_) );
OAI21X1 OAI21X1_1481 ( .A(_3484_), .B(_2969_), .C(_2755_), .Y(_3494_) );
NAND2X1 NAND2X1_636 ( .A(_3493_), .B(_3494_), .Y(_3495_) );
OAI21X1 OAI21X1_1482 ( .A(_3495_), .B(_1134__bF_buf6), .C(_3492_), .Y(_967_) );
XNOR2X1 XNOR2X1_100 ( .A(_3493_), .B(_2757_), .Y(_3496_) );
OAI21X1 OAI21X1_1483 ( .A(_1101__bF_buf19), .B(_1135__bF_buf2_bF_buf2), .C(_3639__29_), .Y(_3497_) );
OAI21X1 OAI21X1_1484 ( .A(_3496_), .B(_1134__bF_buf9), .C(_3497_), .Y(_968_) );
OAI21X1 OAI21X1_1485 ( .A(_3493_), .B(_2757_), .C(_2759_), .Y(_3498_) );
OAI21X1 OAI21X1_1486 ( .A(_2986_), .B(_3493_), .C(_3498_), .Y(_3499_) );
OAI21X1 OAI21X1_1487 ( .A(_1101__bF_buf27), .B(_1135__bF_buf1_bF_buf2), .C(_3639__28_), .Y(_3500_) );
OAI21X1 OAI21X1_1488 ( .A(_3499_), .B(_1134__bF_buf9), .C(_3500_), .Y(_969_) );
NAND2X1 NAND2X1_637 ( .A(bundleAddress_i[29]), .B(_3266_), .Y(_3501_) );
OAI21X1 OAI21X1_1489 ( .A(_3493_), .B(_2986_), .C(_2761_), .Y(_3502_) );
OAI21X1 OAI21X1_1490 ( .A(_3501_), .B(_3493_), .C(_3502_), .Y(_3503_) );
OAI21X1 OAI21X1_1491 ( .A(_1101__bF_buf19), .B(_1135__bF_buf7), .C(_3639__27_), .Y(_3504_) );
OAI21X1 OAI21X1_1492 ( .A(_3503_), .B(_1134__bF_buf9), .C(_3504_), .Y(_970_) );
OAI21X1 OAI21X1_1493 ( .A(_3493_), .B(_3501_), .C(_2763_), .Y(_3505_) );
OAI21X1 OAI21X1_1494 ( .A(_2996_), .B(_3493_), .C(_3505_), .Y(_3506_) );
OAI21X1 OAI21X1_1495 ( .A(_1101__bF_buf22), .B(_1135__bF_buf14_bF_buf2), .C(_3639__26_), .Y(_3507_) );
OAI21X1 OAI21X1_1496 ( .A(_3506_), .B(_1134__bF_buf9), .C(_3507_), .Y(_971_) );
OAI21X1 OAI21X1_1497 ( .A(_3493_), .B(_2996_), .C(_2765_), .Y(_3508_) );
INVX1 INVX1_223 ( .A(_3493_), .Y(_3509_) );
NAND3X1 NAND3X1_65 ( .A(bundleAddress_i[29]), .B(_3274_), .C(_3509_), .Y(_3510_) );
NAND2X1 NAND2X1_638 ( .A(_3508_), .B(_3510_), .Y(_3511_) );
OAI21X1 OAI21X1_1498 ( .A(_1101__bF_buf27), .B(_1135__bF_buf13_bF_buf0), .C(_3639__25_), .Y(_3512_) );
OAI21X1 OAI21X1_1499 ( .A(_3511_), .B(_1134__bF_buf9), .C(_3512_), .Y(_972_) );
XNOR2X1 XNOR2X1_101 ( .A(_3510_), .B(_2767_), .Y(_3513_) );
OAI21X1 OAI21X1_1500 ( .A(_1101__bF_buf10), .B(_1135__bF_buf12_bF_buf3), .C(_3639__24_), .Y(_3514_) );
OAI21X1 OAI21X1_1501 ( .A(_3513_), .B(_1134__bF_buf5), .C(_3514_), .Y(_973_) );
OAI21X1 OAI21X1_1502 ( .A(_3510_), .B(_2767_), .C(_2769_), .Y(_3515_) );
OAI21X1 OAI21X1_1503 ( .A(_3005_), .B(_3510_), .C(_3515_), .Y(_3516_) );
OAI21X1 OAI21X1_1504 ( .A(_1101__bF_buf21), .B(_1135__bF_buf11_bF_buf2), .C(_3639__23_), .Y(_3517_) );
OAI21X1 OAI21X1_1505 ( .A(_3516_), .B(_1134__bF_buf9), .C(_3517_), .Y(_974_) );
OAI21X1 OAI21X1_1506 ( .A(_3510_), .B(_3005_), .C(_2771_), .Y(_3518_) );
OAI21X1 OAI21X1_1507 ( .A(_3015_), .B(_3493_), .C(_3518_), .Y(_3519_) );
OAI21X1 OAI21X1_1508 ( .A(_1101__bF_buf58), .B(_1135__bF_buf10_bF_buf0), .C(_3639__22_), .Y(_3520_) );
OAI21X1 OAI21X1_1509 ( .A(_3519_), .B(_1134__bF_buf6), .C(_3520_), .Y(_975_) );
INVX1 INVX1_224 ( .A(_3015_), .Y(_3521_) );
NAND3X1 NAND3X1_66 ( .A(_3521_), .B(_3440_), .C(_2978_), .Y(_3522_) );
NOR2X1 NOR2X1_225 ( .A(_2773_), .B(_3522_), .Y(_3523_) );
INVX2 INVX2_110 ( .A(_3523_), .Y(_3524_) );
OAI21X1 OAI21X1_1510 ( .A(_3493_), .B(_3015_), .C(_2773_), .Y(_3525_) );
NAND2X1 NAND2X1_639 ( .A(_3525_), .B(_3524_), .Y(_3526_) );
OAI21X1 OAI21X1_1511 ( .A(_1101__bF_buf19), .B(_1135__bF_buf9_bF_buf3), .C(_3639__21_), .Y(_3527_) );
OAI21X1 OAI21X1_1512 ( .A(_3526_), .B(_1134__bF_buf6), .C(_3527_), .Y(_976_) );
XNOR2X1 XNOR2X1_102 ( .A(_3523_), .B(bundleAddress_i[20]), .Y(_3528_) );
OAI21X1 OAI21X1_1513 ( .A(_1101__bF_buf58), .B(_1135__bF_buf8_bF_buf0), .C(_3639__20_), .Y(_3529_) );
OAI21X1 OAI21X1_1514 ( .A(_3528_), .B(_1134__bF_buf6), .C(_3529_), .Y(_977_) );
OAI21X1 OAI21X1_1515 ( .A(_1101__bF_buf9), .B(_1135__bF_buf7_bF_buf1), .C(_3639__19_), .Y(_3530_) );
AOI21X1 AOI21X1_61 ( .A(bundleAddress_i[20]), .B(_3523_), .C(bundleAddress_i[19]), .Y(_3531_) );
OAI21X1 OAI21X1_1516 ( .A(_3524_), .B(_3024_), .C(_613__bF_buf4), .Y(_3532_) );
OAI21X1 OAI21X1_1517 ( .A(_3532_), .B(_3531_), .C(_3530_), .Y(_978_) );
INVX2 INVX2_111 ( .A(_3033_), .Y(_3533_) );
OAI21X1 OAI21X1_1518 ( .A(_3524_), .B(_3024_), .C(_2779_), .Y(_3534_) );
OAI21X1 OAI21X1_1519 ( .A(_3533_), .B(_3522_), .C(_3534_), .Y(_3535_) );
OAI21X1 OAI21X1_1520 ( .A(_1101__bF_buf51), .B(_1135__bF_buf6_bF_buf3), .C(_3639__18_), .Y(_3536_) );
OAI21X1 OAI21X1_1521 ( .A(_3535_), .B(_1134__bF_buf6), .C(_3536_), .Y(_979_) );
NOR2X1 NOR2X1_226 ( .A(_3533_), .B(_3522_), .Y(_3537_) );
NAND2X1 NAND2X1_640 ( .A(bundleAddress_i[17]), .B(_3537_), .Y(_3538_) );
OAI21X1 OAI21X1_1522 ( .A(_3522_), .B(_3533_), .C(_2781_), .Y(_3539_) );
NAND2X1 NAND2X1_641 ( .A(_3539_), .B(_3538_), .Y(_3540_) );
OAI21X1 OAI21X1_1523 ( .A(_1101__bF_buf51), .B(_1135__bF_buf5_bF_buf1), .C(_3639__17_), .Y(_3541_) );
OAI21X1 OAI21X1_1524 ( .A(_3540_), .B(_1134__bF_buf6), .C(_3541_), .Y(_980_) );
OAI21X1 OAI21X1_1525 ( .A(_1101__bF_buf51), .B(_1135__bF_buf4_bF_buf3), .C(_3639__16_), .Y(_3542_) );
INVX1 INVX1_225 ( .A(_3538_), .Y(_3543_) );
NOR2X1 NOR2X1_227 ( .A(bundleAddress_i[16]), .B(_3543_), .Y(_3544_) );
OAI21X1 OAI21X1_1526 ( .A(_3538_), .B(_2783_), .C(_613__bF_buf4), .Y(_3545_) );
OAI21X1 OAI21X1_1527 ( .A(_3544_), .B(_3545_), .C(_3542_), .Y(_981_) );
OAI21X1 OAI21X1_1528 ( .A(_1101__bF_buf58), .B(_1135__bF_buf3_bF_buf0), .C(_3639__15_), .Y(_3546_) );
AOI21X1 AOI21X1_62 ( .A(bundleAddress_i[16]), .B(_3543_), .C(bundleAddress_i[15]), .Y(_3547_) );
OAI21X1 OAI21X1_1529 ( .A(_3538_), .B(_3044_), .C(_613__bF_buf4), .Y(_3548_) );
OAI21X1 OAI21X1_1530 ( .A(_3547_), .B(_3548_), .C(_3546_), .Y(_982_) );
OAI21X1 OAI21X1_1531 ( .A(_3538_), .B(_3044_), .C(_2787_), .Y(_3549_) );
NAND3X1 NAND3X1_67 ( .A(_3440_), .B(_2978_), .C(_3052_), .Y(_3550_) );
NAND2X1 NAND2X1_642 ( .A(_3550_), .B(_3549_), .Y(_3551_) );
OAI21X1 OAI21X1_1532 ( .A(_1101__bF_buf9), .B(_1135__bF_buf2_bF_buf2), .C(_3639__14_), .Y(_3552_) );
OAI21X1 OAI21X1_1533 ( .A(_3551_), .B(_1134__bF_buf2), .C(_3552_), .Y(_983_) );
XNOR2X1 XNOR2X1_103 ( .A(_3550_), .B(_2789_), .Y(_3553_) );
OAI21X1 OAI21X1_1534 ( .A(_1101__bF_buf27), .B(_1135__bF_buf1_bF_buf2), .C(_3639__13_), .Y(_3554_) );
OAI21X1 OAI21X1_1535 ( .A(_3553_), .B(_1134__bF_buf9), .C(_3554_), .Y(_984_) );
OAI21X1 OAI21X1_1536 ( .A(_3550_), .B(_2789_), .C(_2791_), .Y(_3555_) );
OAI21X1 OAI21X1_1537 ( .A(_3067_), .B(_3550_), .C(_3555_), .Y(_3556_) );
OAI21X1 OAI21X1_1538 ( .A(_1101__bF_buf19), .B(_1135__bF_buf7), .C(_3639__12_), .Y(_3557_) );
OAI21X1 OAI21X1_1539 ( .A(_3556_), .B(_1134__bF_buf9), .C(_3557_), .Y(_985_) );
OAI21X1 OAI21X1_1540 ( .A(_1101__bF_buf19), .B(_1135__bF_buf14_bF_buf2), .C(_3639__11_), .Y(_3558_) );
NOR2X1 NOR2X1_228 ( .A(_2789_), .B(_3550_), .Y(_3559_) );
AOI21X1 AOI21X1_63 ( .A(bundleAddress_i[12]), .B(_3559_), .C(bundleAddress_i[11]), .Y(_3560_) );
OAI21X1 OAI21X1_1541 ( .A(_3550_), .B(_3073_), .C(_613__bF_buf2), .Y(_3561_) );
OAI21X1 OAI21X1_1542 ( .A(_3560_), .B(_3561_), .C(_3558_), .Y(_986_) );
OAI21X1 OAI21X1_1543 ( .A(_3550_), .B(_3073_), .C(_2795_), .Y(_3562_) );
OAI21X1 OAI21X1_1544 ( .A(_3075_), .B(_3550_), .C(_3562_), .Y(_3563_) );
OAI21X1 OAI21X1_1545 ( .A(_1101__bF_buf27), .B(_1135__bF_buf13_bF_buf0), .C(_3639__10_), .Y(_3564_) );
OAI21X1 OAI21X1_1546 ( .A(_3563_), .B(_1134__bF_buf9), .C(_3564_), .Y(_987_) );
NOR2X1 NOR2X1_229 ( .A(_3075_), .B(_3550_), .Y(_3565_) );
NAND2X1 NAND2X1_643 ( .A(bundleAddress_i[9]), .B(_3565_), .Y(_3566_) );
OAI21X1 OAI21X1_1547 ( .A(_3550_), .B(_3075_), .C(_2797_), .Y(_3567_) );
NAND2X1 NAND2X1_644 ( .A(_3567_), .B(_3566_), .Y(_3568_) );
OAI21X1 OAI21X1_1548 ( .A(_1101__bF_buf40), .B(_1135__bF_buf12_bF_buf1), .C(_3639__9_), .Y(_3569_) );
OAI21X1 OAI21X1_1549 ( .A(_3568_), .B(_1134__bF_buf0), .C(_3569_), .Y(_988_) );
OAI21X1 OAI21X1_1550 ( .A(_1101__bF_buf40), .B(_1135__bF_buf11_bF_buf2), .C(_3639__8_), .Y(_3570_) );
INVX1 INVX1_226 ( .A(_3566_), .Y(_3571_) );
NOR2X1 NOR2X1_230 ( .A(bundleAddress_i[8]), .B(_3571_), .Y(_3572_) );
OAI21X1 OAI21X1_1551 ( .A(_3566_), .B(_2799_), .C(_613__bF_buf2), .Y(_3573_) );
OAI21X1 OAI21X1_1552 ( .A(_3572_), .B(_3573_), .C(_3570_), .Y(_989_) );
OAI21X1 OAI21X1_1553 ( .A(_1101__bF_buf58), .B(_1135__bF_buf10_bF_buf0), .C(_3639__7_), .Y(_3574_) );
AOI21X1 AOI21X1_64 ( .A(bundleAddress_i[8]), .B(_3571_), .C(bundleAddress_i[7]), .Y(_3575_) );
OAI21X1 OAI21X1_1554 ( .A(_3566_), .B(_3087_), .C(_613__bF_buf2), .Y(_3576_) );
OAI21X1 OAI21X1_1555 ( .A(_3575_), .B(_3576_), .C(_3574_), .Y(_990_) );
INVX1 INVX1_227 ( .A(_3639__6_), .Y(_3577_) );
OAI21X1 OAI21X1_1556 ( .A(_3566_), .B(_3087_), .C(_2803_), .Y(_3578_) );
OR2X2 OR2X2_21 ( .A(_3550_), .B(_3095_), .Y(_3579_) );
NAND3X1 NAND3X1_68 ( .A(_613__bF_buf2), .B(_3579_), .C(_3578_), .Y(_3580_) );
OAI21X1 OAI21X1_1557 ( .A(_3577_), .B(_613__bF_buf2), .C(_3580_), .Y(_991_) );
NOR2X1 NOR2X1_231 ( .A(_3095_), .B(_3550_), .Y(_3581_) );
NAND2X1 NAND2X1_645 ( .A(bundleAddress_i[5]), .B(_3581_), .Y(_3582_) );
OAI21X1 OAI21X1_1558 ( .A(_3550_), .B(_3095_), .C(_2805_), .Y(_3583_) );
NAND2X1 NAND2X1_646 ( .A(_3583_), .B(_3582_), .Y(_3584_) );
OAI21X1 OAI21X1_1559 ( .A(_1101__bF_buf58), .B(_1135__bF_buf9_bF_buf3), .C(_3639__5_), .Y(_3585_) );
OAI21X1 OAI21X1_1560 ( .A(_3584_), .B(_1134__bF_buf6), .C(_3585_), .Y(_992_) );
OAI21X1 OAI21X1_1561 ( .A(_1101__bF_buf38), .B(_1135__bF_buf8_bF_buf0), .C(_3639__4_), .Y(_3586_) );
INVX2 INVX2_112 ( .A(_3582_), .Y(_3587_) );
NOR2X1 NOR2X1_232 ( .A(bundleAddress_i[4]), .B(_3587_), .Y(_3588_) );
OAI21X1 OAI21X1_1562 ( .A(_3582_), .B(_2807_), .C(_613__bF_buf4), .Y(_3589_) );
OAI21X1 OAI21X1_1563 ( .A(_3588_), .B(_3589_), .C(_3586_), .Y(_993_) );
OAI21X1 OAI21X1_1564 ( .A(_1101__bF_buf38), .B(_1135__bF_buf7_bF_buf3), .C(_3639__3_), .Y(_3590_) );
AOI21X1 AOI21X1_65 ( .A(bundleAddress_i[4]), .B(_3587_), .C(bundleAddress_i[3]), .Y(_3591_) );
OAI21X1 OAI21X1_1565 ( .A(_3579_), .B(_3114_), .C(_613__bF_buf4), .Y(_3592_) );
OAI21X1 OAI21X1_1566 ( .A(_3591_), .B(_3592_), .C(_3590_), .Y(_994_) );
AOI21X1 AOI21X1_66 ( .A(_3109_), .B(_3587_), .C(bundleAddress_i[2]), .Y(_3593_) );
OAI21X1 OAI21X1_1567 ( .A(_3579_), .B(_3116_), .C(_613__bF_buf4), .Y(_3594_) );
OAI21X1 OAI21X1_1568 ( .A(_1101__bF_buf58), .B(_1135__bF_buf6_bF_buf3), .C(_3639__2_), .Y(_3595_) );
OAI21X1 OAI21X1_1569 ( .A(_3593_), .B(_3594_), .C(_3595_), .Y(_995_) );
NAND3X1 NAND3X1_69 ( .A(bundleAddress_i[1]), .B(_3115_), .C(_3581_), .Y(_3596_) );
OAI21X1 OAI21X1_1570 ( .A(_3579_), .B(_3116_), .C(_2813_), .Y(_3597_) );
NAND2X1 NAND2X1_647 ( .A(_3596_), .B(_3597_), .Y(_3598_) );
OAI21X1 OAI21X1_1571 ( .A(_1101__bF_buf51), .B(_1135__bF_buf5_bF_buf1), .C(_3639__1_), .Y(_3599_) );
OAI21X1 OAI21X1_1572 ( .A(_3598_), .B(_1134__bF_buf6), .C(_3599_), .Y(_996_) );
XNOR2X1 XNOR2X1_104 ( .A(_3596_), .B(_2815_), .Y(_3600_) );
OAI21X1 OAI21X1_1573 ( .A(_1101__bF_buf17), .B(_1135__bF_buf4_bF_buf3), .C(_3639__0_), .Y(_3601_) );
OAI21X1 OAI21X1_1574 ( .A(_3600_), .B(_1134__bF_buf6), .C(_3601_), .Y(_997_) );
INVX2 INVX2_113 ( .A(is64Bit_i), .Y(_3602_) );
NAND2X1 NAND2X1_648 ( .A(_3648_), .B(_1031__bF_buf60), .Y(_3603_) );
OAI21X1 OAI21X1_1575 ( .A(_1031__bF_buf60), .B(_3602_), .C(_3603_), .Y(_998_) );
NAND2X1 NAND2X1_649 ( .A(_3649_), .B(_1039__bF_buf24), .Y(_3604_) );
OAI21X1 OAI21X1_1576 ( .A(_3602_), .B(_1039__bF_buf24), .C(_3604_), .Y(_999_) );
OAI21X1 OAI21X1_1577 ( .A(_1100__bF_buf10_bF_buf1), .B(_1031__bF_buf64), .C(_3650_), .Y(_3605_) );
OAI21X1 OAI21X1_1578 ( .A(_1101__bF_buf50), .B(_3602_), .C(_3605_), .Y(_1000_) );
OAI21X1 OAI21X1_1579 ( .A(_1101__bF_buf50), .B(_1135__bF_buf3_bF_buf3), .C(_3651_), .Y(_3606_) );
OAI21X1 OAI21X1_1580 ( .A(_3602_), .B(_1134__bF_buf5), .C(_3606_), .Y(_1001_) );
NAND2X1 NAND2X1_650 ( .A(_3656__31_), .B(_1031__bF_buf75), .Y(_3607_) );
OAI21X1 OAI21X1_1581 ( .A(_1031__bF_buf66), .B(_1038_), .C(_3607_), .Y(_1002_) );
NAND2X1 NAND2X1_651 ( .A(_3656__30_), .B(_1031__bF_buf72), .Y(_3608_) );
OAI21X1 OAI21X1_1582 ( .A(_1031__bF_buf72), .B(_1041_), .C(_3608_), .Y(_1003_) );
NAND2X1 NAND2X1_652 ( .A(_3656__29_), .B(_1031__bF_buf39), .Y(_3609_) );
OAI21X1 OAI21X1_1583 ( .A(_1031__bF_buf39), .B(_1043_), .C(_3609_), .Y(_1004_) );
NAND2X1 NAND2X1_653 ( .A(_3656__28_), .B(_1031__bF_buf77), .Y(_3610_) );
OAI21X1 OAI21X1_1584 ( .A(_1031__bF_buf77), .B(_1045_), .C(_3610_), .Y(_1005_) );
NAND2X1 NAND2X1_654 ( .A(_3656__27_), .B(_1031__bF_buf21), .Y(_3611_) );
OAI21X1 OAI21X1_1585 ( .A(_1031__bF_buf21), .B(_1047_), .C(_3611_), .Y(_1006_) );
NAND2X1 NAND2X1_655 ( .A(_3656__26_), .B(_1031__bF_buf50), .Y(_3612_) );
OAI21X1 OAI21X1_1586 ( .A(_1031__bF_buf50), .B(_1049_), .C(_3612_), .Y(_1007_) );
NAND2X1 NAND2X1_656 ( .A(_3656__25_), .B(_1031__bF_buf61), .Y(_3613_) );
OAI21X1 OAI21X1_1587 ( .A(_1031__bF_buf61), .B(_1051_), .C(_3613_), .Y(_1008_) );
NAND2X1 NAND2X1_657 ( .A(_3656__24_), .B(_1031__bF_buf52), .Y(_3614_) );
OAI21X1 OAI21X1_1588 ( .A(_1031__bF_buf52), .B(_1053_), .C(_3614_), .Y(_1009_) );
NAND2X1 NAND2X1_658 ( .A(_3656__23_), .B(_1031__bF_buf39), .Y(_3615_) );
OAI21X1 OAI21X1_1589 ( .A(_1031__bF_buf39), .B(_1055_), .C(_3615_), .Y(_1010_) );
NAND2X1 NAND2X1_659 ( .A(_3656__22_), .B(_1031__bF_buf8), .Y(_3616_) );
OAI21X1 OAI21X1_1590 ( .A(_1031__bF_buf8), .B(_1057_), .C(_3616_), .Y(_1011_) );
NAND2X1 NAND2X1_660 ( .A(_3656__21_), .B(_1031__bF_buf39), .Y(_3617_) );
OAI21X1 OAI21X1_1591 ( .A(_1031__bF_buf39), .B(_1059_), .C(_3617_), .Y(_1012_) );
NAND2X1 NAND2X1_661 ( .A(_3656__20_), .B(_1031__bF_buf22), .Y(_3618_) );
OAI21X1 OAI21X1_1592 ( .A(_1031__bF_buf22), .B(_1061_), .C(_3618_), .Y(_1013_) );
NAND2X1 NAND2X1_662 ( .A(_3656__19_), .B(_1031__bF_buf12), .Y(_3619_) );
OAI21X1 OAI21X1_1593 ( .A(_1031__bF_buf12), .B(_1063_), .C(_3619_), .Y(_1014_) );
NAND2X1 NAND2X1_663 ( .A(_3656__18_), .B(_1031__bF_buf25), .Y(_3620_) );
OAI21X1 OAI21X1_1594 ( .A(_1031__bF_buf25), .B(_1065_), .C(_3620_), .Y(_1015_) );
NAND2X1 NAND2X1_664 ( .A(_3656__17_), .B(_1031__bF_buf75), .Y(_3621_) );
OAI21X1 OAI21X1_1595 ( .A(_1031__bF_buf75), .B(_1067_), .C(_3621_), .Y(_1016_) );
NAND2X1 NAND2X1_665 ( .A(_3656__16_), .B(_1031__bF_buf8), .Y(_3622_) );
OAI21X1 OAI21X1_1596 ( .A(_1031__bF_buf8), .B(_1069_), .C(_3622_), .Y(_1017_) );
NAND2X1 NAND2X1_666 ( .A(_3656__15_), .B(_1031__bF_buf76), .Y(_3623_) );
OAI21X1 OAI21X1_1597 ( .A(_1031__bF_buf76), .B(_1071_), .C(_3623_), .Y(_1018_) );
NAND2X1 NAND2X1_667 ( .A(_3656__14_), .B(_1031__bF_buf8), .Y(_3624_) );
OAI21X1 OAI21X1_1598 ( .A(_1031__bF_buf70), .B(_1073_), .C(_3624_), .Y(_1019_) );
NAND2X1 NAND2X1_668 ( .A(_3656__13_), .B(_1031__bF_buf22), .Y(_3625_) );
OAI21X1 OAI21X1_1599 ( .A(_1031__bF_buf12), .B(_1075_), .C(_3625_), .Y(_1020_) );
NAND2X1 NAND2X1_669 ( .A(_3656__12_), .B(_1031__bF_buf67), .Y(_3626_) );
OAI21X1 OAI21X1_1600 ( .A(_1031__bF_buf67), .B(_1077_), .C(_3626_), .Y(_1021_) );
NAND2X1 NAND2X1_670 ( .A(_3656__11_), .B(_1031__bF_buf49), .Y(_3627_) );
OAI21X1 OAI21X1_1601 ( .A(_1031__bF_buf49), .B(_1079_), .C(_3627_), .Y(_1022_) );
NAND2X1 NAND2X1_671 ( .A(_3656__10_), .B(_1031__bF_buf22), .Y(_3628_) );
OAI21X1 OAI21X1_1602 ( .A(_1031__bF_buf36), .B(_1081_), .C(_3628_), .Y(_1023_) );
NAND2X1 NAND2X1_672 ( .A(_3656__9_), .B(_1031__bF_buf9), .Y(_3629_) );
OAI21X1 OAI21X1_1603 ( .A(_1031__bF_buf29), .B(_1083_), .C(_3629_), .Y(_1024_) );
NAND2X1 NAND2X1_673 ( .A(_3656__8_), .B(_1031__bF_buf56), .Y(_3630_) );
OAI21X1 OAI21X1_1604 ( .A(_1031__bF_buf56), .B(_1085_), .C(_3630_), .Y(_1025_) );
NAND2X1 NAND2X1_674 ( .A(_3656__7_), .B(_1031__bF_buf19), .Y(_3631_) );
OAI21X1 OAI21X1_1605 ( .A(_1031__bF_buf19), .B(_1087_), .C(_3631_), .Y(_1026_) );
NAND2X1 NAND2X1_675 ( .A(_3656__6_), .B(_1031__bF_buf62), .Y(_3632_) );
OAI21X1 OAI21X1_1606 ( .A(_1031__bF_buf62), .B(_1089_), .C(_3632_), .Y(_1027_) );
NAND2X1 NAND2X1_676 ( .A(_3656__5_), .B(_1031__bF_buf39), .Y(_3633_) );
OAI21X1 OAI21X1_1607 ( .A(_1031__bF_buf39), .B(_1091_), .C(_3633_), .Y(_1028_) );
NAND2X1 NAND2X1_677 ( .A(_3656__4_), .B(_1031__bF_buf9), .Y(_3634_) );
OAI21X1 OAI21X1_1608 ( .A(_1031__bF_buf9), .B(_1093_), .C(_3634_), .Y(_1029_) );
NAND2X1 NAND2X1_678 ( .A(_3656__3_), .B(_1031__bF_buf20), .Y(_3635_) );
OAI21X1 OAI21X1_1609 ( .A(_1031__bF_buf20), .B(_1095_), .C(_3635_), .Y(_1030_) );
INVX8 INVX8_4 ( .A(enable_i_bF_buf2), .Y(_1031_) );
INVX2 INVX2_114 ( .A(bundlePid_i[2]), .Y(_1032_) );
NAND2X1 NAND2X1_679 ( .A(_3656__2_), .B(_1031__bF_buf57), .Y(_1033_) );
OAI21X1 OAI21X1_1610 ( .A(_1031__bF_buf50), .B(_1032_), .C(_1033_), .Y(_0_) );
INVX2 INVX2_115 ( .A(bundlePid_i[1]), .Y(_1034_) );
NAND2X1 NAND2X1_680 ( .A(_3656__1_), .B(_1031__bF_buf15), .Y(_1035_) );
OAI21X1 OAI21X1_1611 ( .A(_1031__bF_buf15), .B(_1034_), .C(_1035_), .Y(_1_) );
INVX2 INVX2_116 ( .A(bundlePid_i[0]), .Y(_1036_) );
NAND2X1 NAND2X1_681 ( .A(_3656__0_), .B(_1031__bF_buf68), .Y(_1037_) );
OAI21X1 OAI21X1_1612 ( .A(_1031__bF_buf68), .B(_1036_), .C(_1037_), .Y(_2_) );
INVX2 INVX2_117 ( .A(bundlePid_i[31]), .Y(_1038_) );
OAI21X1 OAI21X1_1613 ( .A(bundleLen_i[1]), .B(bundleLen_i[0]), .C(enable_i_bF_buf2), .Y(_1039_) );
NAND2X1 NAND2X1_682 ( .A(_3657__31_), .B(_1039__bF_buf3), .Y(_1040_) );
OAI21X1 OAI21X1_1614 ( .A(_1038_), .B(_1039__bF_buf34), .C(_1040_), .Y(_3_) );
INVX2 INVX2_118 ( .A(bundlePid_i[30]), .Y(_1041_) );
NAND2X1 NAND2X1_683 ( .A(_3657__30_), .B(_1039__bF_buf2), .Y(_1042_) );
OAI21X1 OAI21X1_1615 ( .A(_1041_), .B(_1039__bF_buf2), .C(_1042_), .Y(_4_) );
INVX2 INVX2_119 ( .A(bundlePid_i[29]), .Y(_1043_) );
NAND2X1 NAND2X1_684 ( .A(_3657__29_), .B(_1039__bF_buf10), .Y(_1044_) );
OAI21X1 OAI21X1_1616 ( .A(_1043_), .B(_1039__bF_buf10), .C(_1044_), .Y(_5_) );
INVX2 INVX2_120 ( .A(bundlePid_i[28]), .Y(_1045_) );
NAND2X1 NAND2X1_685 ( .A(_3657__28_), .B(_1039__bF_buf45), .Y(_1046_) );
OAI21X1 OAI21X1_1617 ( .A(_1045_), .B(_1039__bF_buf45), .C(_1046_), .Y(_6_) );
INVX2 INVX2_121 ( .A(bundlePid_i[27]), .Y(_1047_) );
NAND2X1 NAND2X1_686 ( .A(_3657__27_), .B(_1039__bF_buf57), .Y(_1048_) );
OAI21X1 OAI21X1_1618 ( .A(_1047_), .B(_1039__bF_buf57), .C(_1048_), .Y(_7_) );
INVX2 INVX2_122 ( .A(bundlePid_i[26]), .Y(_1049_) );
NAND2X1 NAND2X1_687 ( .A(_3657__26_), .B(_1039__bF_buf31), .Y(_1050_) );
OAI21X1 OAI21X1_1619 ( .A(_1049_), .B(_1039__bF_buf31), .C(_1050_), .Y(_8_) );
INVX2 INVX2_123 ( .A(bundlePid_i[25]), .Y(_1051_) );
NAND2X1 NAND2X1_688 ( .A(_3657__25_), .B(_1039__bF_buf20), .Y(_1052_) );
OAI21X1 OAI21X1_1620 ( .A(_1051_), .B(_1039__bF_buf20), .C(_1052_), .Y(_9_) );
INVX2 INVX2_124 ( .A(bundlePid_i[24]), .Y(_1053_) );
NAND2X1 NAND2X1_689 ( .A(_3657__24_), .B(_1039__bF_buf30), .Y(_1054_) );
OAI21X1 OAI21X1_1621 ( .A(_1053_), .B(_1039__bF_buf30), .C(_1054_), .Y(_10_) );
INVX2 INVX2_125 ( .A(bundlePid_i[23]), .Y(_1055_) );
NAND2X1 NAND2X1_690 ( .A(_3657__23_), .B(_1039__bF_buf44), .Y(_1056_) );
OAI21X1 OAI21X1_1622 ( .A(_1055_), .B(_1039__bF_buf44), .C(_1056_), .Y(_11_) );
INVX2 INVX2_126 ( .A(bundlePid_i[22]), .Y(_1057_) );
NAND2X1 NAND2X1_691 ( .A(_3657__22_), .B(_1039__bF_buf19), .Y(_1058_) );
OAI21X1 OAI21X1_1623 ( .A(_1057_), .B(_1039__bF_buf19), .C(_1058_), .Y(_12_) );
INVX2 INVX2_127 ( .A(bundlePid_i[21]), .Y(_1059_) );
NAND2X1 NAND2X1_692 ( .A(_3657__21_), .B(_1039__bF_buf44), .Y(_1060_) );
OAI21X1 OAI21X1_1624 ( .A(_1059_), .B(_1039__bF_buf42), .C(_1060_), .Y(_13_) );
INVX2 INVX2_128 ( .A(bundlePid_i[20]), .Y(_1061_) );
NAND2X1 NAND2X1_693 ( .A(_3657__20_), .B(_1039__bF_buf26), .Y(_1062_) );
OAI21X1 OAI21X1_1625 ( .A(_1061_), .B(_1039__bF_buf26), .C(_1062_), .Y(_14_) );
INVX2 INVX2_129 ( .A(bundlePid_i[19]), .Y(_1063_) );
NAND2X1 NAND2X1_694 ( .A(_3657__19_), .B(_1039__bF_buf54), .Y(_1064_) );
OAI21X1 OAI21X1_1626 ( .A(_1063_), .B(_1039__bF_buf54), .C(_1064_), .Y(_15_) );
INVX2 INVX2_130 ( .A(bundlePid_i[18]), .Y(_1065_) );
NAND2X1 NAND2X1_695 ( .A(_3657__18_), .B(_1039__bF_buf25), .Y(_1066_) );
OAI21X1 OAI21X1_1627 ( .A(_1065_), .B(_1039__bF_buf25), .C(_1066_), .Y(_16_) );
INVX2 INVX2_131 ( .A(bundlePid_i[17]), .Y(_1067_) );
NAND2X1 NAND2X1_696 ( .A(_3657__17_), .B(_1039__bF_buf34), .Y(_1068_) );
OAI21X1 OAI21X1_1628 ( .A(_1067_), .B(_1039__bF_buf34), .C(_1068_), .Y(_17_) );
INVX2 INVX2_132 ( .A(bundlePid_i[16]), .Y(_1069_) );
NAND2X1 NAND2X1_697 ( .A(_3657__16_), .B(_1039__bF_buf19), .Y(_1070_) );
OAI21X1 OAI21X1_1629 ( .A(_1069_), .B(_1039__bF_buf19), .C(_1070_), .Y(_18_) );
INVX2 INVX2_133 ( .A(bundlePid_i[15]), .Y(_1071_) );
NAND2X1 NAND2X1_698 ( .A(_3657__15_), .B(_1039__bF_buf6), .Y(_1072_) );
OAI21X1 OAI21X1_1630 ( .A(_1071_), .B(_1039__bF_buf39), .C(_1072_), .Y(_19_) );
INVX2 INVX2_134 ( .A(bundlePid_i[14]), .Y(_1073_) );
NAND2X1 NAND2X1_699 ( .A(_3657__14_), .B(_1039__bF_buf17), .Y(_1074_) );
OAI21X1 OAI21X1_1631 ( .A(_1073_), .B(_1039__bF_buf17), .C(_1074_), .Y(_20_) );
INVX2 INVX2_135 ( .A(bundlePid_i[13]), .Y(_1075_) );
NAND2X1 NAND2X1_700 ( .A(_3657__13_), .B(_1039__bF_buf7), .Y(_1076_) );
OAI21X1 OAI21X1_1632 ( .A(_1075_), .B(_1039__bF_buf54), .C(_1076_), .Y(_21_) );
INVX2 INVX2_136 ( .A(bundlePid_i[12]), .Y(_1077_) );
NAND2X1 NAND2X1_701 ( .A(_3657__12_), .B(_1039__bF_buf4), .Y(_1078_) );
OAI21X1 OAI21X1_1633 ( .A(_1077_), .B(_1039__bF_buf4), .C(_1078_), .Y(_22_) );
INVX2 INVX2_137 ( .A(bundlePid_i[11]), .Y(_1079_) );
NAND2X1 NAND2X1_702 ( .A(_3657__11_), .B(_1039__bF_buf42), .Y(_1080_) );
OAI21X1 OAI21X1_1634 ( .A(_1079_), .B(_1039__bF_buf18), .C(_1080_), .Y(_23_) );
INVX2 INVX2_138 ( .A(bundlePid_i[10]), .Y(_1081_) );
NAND2X1 NAND2X1_703 ( .A(_3657__10_), .B(_1039__bF_buf26), .Y(_1082_) );
OAI21X1 OAI21X1_1635 ( .A(_1081_), .B(_1039__bF_buf26), .C(_1082_), .Y(_24_) );
INVX2 INVX2_139 ( .A(bundlePid_i[9]), .Y(_1083_) );
NAND2X1 NAND2X1_704 ( .A(_3657__9_), .B(_1039__bF_buf14), .Y(_1084_) );
OAI21X1 OAI21X1_1636 ( .A(_1083_), .B(_1039__bF_buf14), .C(_1084_), .Y(_25_) );
INVX2 INVX2_140 ( .A(bundlePid_i[8]), .Y(_1085_) );
NAND2X1 NAND2X1_705 ( .A(_3657__8_), .B(_1039__bF_buf32), .Y(_1086_) );
OAI21X1 OAI21X1_1637 ( .A(_1085_), .B(_1039__bF_buf32), .C(_1086_), .Y(_26_) );
INVX2 INVX2_141 ( .A(bundlePid_i[7]), .Y(_1087_) );
NAND2X1 NAND2X1_706 ( .A(_3657__7_), .B(_1039__bF_buf45), .Y(_1088_) );
OAI21X1 OAI21X1_1638 ( .A(_1087_), .B(_1039__bF_buf45), .C(_1088_), .Y(_27_) );
INVX2 INVX2_142 ( .A(bundlePid_i[6]), .Y(_1089_) );
NAND2X1 NAND2X1_707 ( .A(_3657__6_), .B(_1039__bF_buf28), .Y(_1090_) );
OAI21X1 OAI21X1_1639 ( .A(_1089_), .B(_1039__bF_buf28), .C(_1090_), .Y(_28_) );
INVX2 INVX2_143 ( .A(bundlePid_i[5]), .Y(_1091_) );
NAND2X1 NAND2X1_708 ( .A(_3657__5_), .B(_1039__bF_buf10), .Y(_1092_) );
OAI21X1 OAI21X1_1640 ( .A(_1091_), .B(_1039__bF_buf10), .C(_1092_), .Y(_29_) );
INVX2 INVX2_144 ( .A(bundlePid_i[4]), .Y(_1093_) );
NAND2X1 NAND2X1_709 ( .A(_3657__4_), .B(_1039__bF_buf47), .Y(_1094_) );
OAI21X1 OAI21X1_1641 ( .A(_1093_), .B(_1039__bF_buf47), .C(_1094_), .Y(_30_) );
INVX2 INVX2_145 ( .A(bundlePid_i[3]), .Y(_1095_) );
NAND2X1 NAND2X1_710 ( .A(_3657__3_), .B(_1039__bF_buf40), .Y(_1096_) );
OAI21X1 OAI21X1_1642 ( .A(_1095_), .B(_1039__bF_buf40), .C(_1096_), .Y(_31_) );
NAND2X1 NAND2X1_711 ( .A(_3657__2_), .B(_1039__bF_buf49), .Y(_1097_) );
OAI21X1 OAI21X1_1643 ( .A(_1032_), .B(_1039__bF_buf49), .C(_1097_), .Y(_32_) );
NAND2X1 NAND2X1_712 ( .A(_3657__1_), .B(_1039__bF_buf12), .Y(_1098_) );
OAI21X1 OAI21X1_1644 ( .A(_1034_), .B(_1039__bF_buf12), .C(_1098_), .Y(_33_) );
NAND2X1 NAND2X1_713 ( .A(_3657__0_), .B(_1039__bF_buf20), .Y(_1099_) );
OAI21X1 OAI21X1_1645 ( .A(_1036_), .B(_1039__bF_buf20), .C(_1099_), .Y(_34_) );
INVX8 INVX8_5 ( .A(bundleLen_i[0]), .Y(_1100_) );
NOR2X1 NOR2X1_233 ( .A(_1100__bF_buf9_bF_buf1), .B(_1031__bF_buf44), .Y(_612_) );
INVX8 INVX8_6 ( .A(_612__bF_buf1), .Y(_1101_) );
OAI21X1 OAI21X1_1646 ( .A(_1100__bF_buf8_bF_buf3), .B(_1031__bF_buf47), .C(_3658__31_), .Y(_1102_) );
OAI21X1 OAI21X1_1647 ( .A(_1101__bF_buf7), .B(_1038_), .C(_1102_), .Y(_35_) );
OAI21X1 OAI21X1_1648 ( .A(_1100__bF_buf7_bF_buf1), .B(_1031__bF_buf72), .C(_3658__30_), .Y(_1103_) );
OAI21X1 OAI21X1_1649 ( .A(_1101__bF_buf29), .B(_1041_), .C(_1103_), .Y(_36_) );
OAI21X1 OAI21X1_1650 ( .A(_1100__bF_buf3), .B(_1031__bF_buf56), .C(_3658__29_), .Y(_1104_) );
OAI21X1 OAI21X1_1651 ( .A(_1101__bF_buf56), .B(_1043_), .C(_1104_), .Y(_37_) );
OAI21X1 OAI21X1_1652 ( .A(_1100__bF_buf5), .B(_1031__bF_buf11), .C(_3658__28_), .Y(_1105_) );
OAI21X1 OAI21X1_1653 ( .A(_1101__bF_buf41), .B(_1045_), .C(_1105_), .Y(_38_) );
OAI21X1 OAI21X1_1654 ( .A(_1100__bF_buf4), .B(_1031__bF_buf21), .C(_3658__27_), .Y(_1106_) );
OAI21X1 OAI21X1_1655 ( .A(_1101__bF_buf54), .B(_1047_), .C(_1106_), .Y(_39_) );
OAI21X1 OAI21X1_1656 ( .A(_1100__bF_buf2), .B(_1031__bF_buf50), .C(_3658__26_), .Y(_1107_) );
OAI21X1 OAI21X1_1657 ( .A(_1101__bF_buf25), .B(_1049_), .C(_1107_), .Y(_40_) );
OAI21X1 OAI21X1_1658 ( .A(_1100__bF_buf6), .B(_1031__bF_buf61), .C(_3658__25_), .Y(_1108_) );
OAI21X1 OAI21X1_1659 ( .A(_1101__bF_buf6), .B(_1051_), .C(_1108_), .Y(_41_) );
OAI21X1 OAI21X1_1660 ( .A(_1100__bF_buf12), .B(_1031__bF_buf27), .C(_3658__24_), .Y(_1109_) );
OAI21X1 OAI21X1_1661 ( .A(_1101__bF_buf11), .B(_1053_), .C(_1109_), .Y(_42_) );
OAI21X1 OAI21X1_1662 ( .A(_1100__bF_buf3), .B(_1031__bF_buf39), .C(_3658__23_), .Y(_1110_) );
OAI21X1 OAI21X1_1663 ( .A(_1101__bF_buf39), .B(_1055_), .C(_1110_), .Y(_43_) );
OAI21X1 OAI21X1_1664 ( .A(_1100__bF_buf14_bF_buf1), .B(_1031__bF_buf13), .C(_3658__22_), .Y(_1111_) );
OAI21X1 OAI21X1_1665 ( .A(_1101__bF_buf39), .B(_1057_), .C(_1111_), .Y(_44_) );
OAI21X1 OAI21X1_1666 ( .A(_1100__bF_buf13_bF_buf3), .B(_1031__bF_buf49), .C(_3658__21_), .Y(_1112_) );
OAI21X1 OAI21X1_1667 ( .A(_1101__bF_buf39), .B(_1059_), .C(_1112_), .Y(_45_) );
OAI21X1 OAI21X1_1668 ( .A(_1100__bF_buf12_bF_buf3), .B(_1031__bF_buf41), .C(_3658__20_), .Y(_1113_) );
OAI21X1 OAI21X1_1669 ( .A(_1101__bF_buf28), .B(_1061_), .C(_1113_), .Y(_46_) );
OAI21X1 OAI21X1_1670 ( .A(_1100__bF_buf11_bF_buf2), .B(_1031__bF_buf12), .C(_3658__19_), .Y(_1114_) );
OAI21X1 OAI21X1_1671 ( .A(_1101__bF_buf3), .B(_1063_), .C(_1114_), .Y(_47_) );
OAI21X1 OAI21X1_1672 ( .A(_1100__bF_buf10_bF_buf1), .B(_1031__bF_buf64), .C(_3658__18_), .Y(_1115_) );
OAI21X1 OAI21X1_1673 ( .A(_1101__bF_buf22), .B(_1065_), .C(_1115_), .Y(_48_) );
OAI21X1 OAI21X1_1674 ( .A(_1100__bF_buf9_bF_buf1), .B(_1031__bF_buf47), .C(_3658__17_), .Y(_1116_) );
OAI21X1 OAI21X1_1675 ( .A(_1101__bF_buf7), .B(_1067_), .C(_1116_), .Y(_49_) );
OAI21X1 OAI21X1_1676 ( .A(_1100__bF_buf8_bF_buf3), .B(_1031__bF_buf47), .C(_3658__16_), .Y(_1117_) );
OAI21X1 OAI21X1_1677 ( .A(_1101__bF_buf9), .B(_1069_), .C(_1117_), .Y(_50_) );
OAI21X1 OAI21X1_1678 ( .A(_1100__bF_buf7_bF_buf2), .B(_1031__bF_buf20), .C(_3658__15_), .Y(_1118_) );
OAI21X1 OAI21X1_1679 ( .A(_1101__bF_buf53), .B(_1071_), .C(_1118_), .Y(_51_) );
OAI21X1 OAI21X1_1680 ( .A(_1100__bF_buf3), .B(_1031__bF_buf70), .C(_3658__14_), .Y(_1119_) );
OAI21X1 OAI21X1_1681 ( .A(_1101__bF_buf1), .B(_1073_), .C(_1119_), .Y(_52_) );
OAI21X1 OAI21X1_1682 ( .A(_1100__bF_buf4), .B(_1031__bF_buf22), .C(_3658__13_), .Y(_1120_) );
OAI21X1 OAI21X1_1683 ( .A(_1101__bF_buf54), .B(_1075_), .C(_1120_), .Y(_53_) );
OAI21X1 OAI21X1_1684 ( .A(_1100__bF_buf4), .B(_1031__bF_buf26), .C(_3658__12_), .Y(_1121_) );
OAI21X1 OAI21X1_1685 ( .A(_1101__bF_buf3), .B(_1077_), .C(_1121_), .Y(_54_) );
OAI21X1 OAI21X1_1686 ( .A(_1100__bF_buf3), .B(_1031__bF_buf49), .C(_3658__11_), .Y(_1122_) );
OAI21X1 OAI21X1_1687 ( .A(_1101__bF_buf39), .B(_1079_), .C(_1122_), .Y(_55_) );
OAI21X1 OAI21X1_1688 ( .A(_1100__bF_buf4), .B(_1031__bF_buf36), .C(_3658__10_), .Y(_1123_) );
OAI21X1 OAI21X1_1689 ( .A(_1101__bF_buf43), .B(_1081_), .C(_1123_), .Y(_56_) );
OAI21X1 OAI21X1_1690 ( .A(_1100__bF_buf12), .B(_1031__bF_buf27), .C(_3658__9_), .Y(_1124_) );
OAI21X1 OAI21X1_1691 ( .A(_1101__bF_buf11), .B(_1083_), .C(_1124_), .Y(_57_) );
OAI21X1 OAI21X1_1692 ( .A(_1100__bF_buf3), .B(_1031__bF_buf56), .C(_3658__8_), .Y(_1125_) );
OAI21X1 OAI21X1_1693 ( .A(_1101__bF_buf56), .B(_1085_), .C(_1125_), .Y(_58_) );
OAI21X1 OAI21X1_1694 ( .A(_1100__bF_buf14_bF_buf2), .B(_1031__bF_buf29), .C(_3658__7_), .Y(_1126_) );
OAI21X1 OAI21X1_1695 ( .A(_1101__bF_buf30), .B(_1087_), .C(_1126_), .Y(_59_) );
OAI21X1 OAI21X1_1696 ( .A(_1100__bF_buf13_bF_buf0), .B(_1031__bF_buf54), .C(_3658__6_), .Y(_1127_) );
OAI21X1 OAI21X1_1697 ( .A(_1101__bF_buf32), .B(_1089_), .C(_1127_), .Y(_60_) );
OAI21X1 OAI21X1_1698 ( .A(_1100__bF_buf12_bF_buf1), .B(_1031__bF_buf75), .C(_3658__5_), .Y(_1128_) );
OAI21X1 OAI21X1_1699 ( .A(_1101__bF_buf39), .B(_1091_), .C(_1128_), .Y(_61_) );
OAI21X1 OAI21X1_1700 ( .A(_1100__bF_buf11_bF_buf3), .B(_1031__bF_buf9), .C(_3658__4_), .Y(_1129_) );
OAI21X1 OAI21X1_1701 ( .A(_1101__bF_buf11), .B(_1093_), .C(_1129_), .Y(_62_) );
OAI21X1 OAI21X1_1702 ( .A(_1100__bF_buf10_bF_buf3), .B(_1031__bF_buf26), .C(_3658__3_), .Y(_1130_) );
OAI21X1 OAI21X1_1703 ( .A(_1101__bF_buf0), .B(_1095_), .C(_1130_), .Y(_63_) );
OAI21X1 OAI21X1_1704 ( .A(_1100__bF_buf9_bF_buf0), .B(_1031__bF_buf57), .C(_3658__2_), .Y(_1131_) );
OAI21X1 OAI21X1_1705 ( .A(_1101__bF_buf35), .B(_1032_), .C(_1131_), .Y(_64_) );
OAI21X1 OAI21X1_1706 ( .A(_1100__bF_buf8_bF_buf1), .B(_1031__bF_buf0), .C(_3658__1_), .Y(_1132_) );
OAI21X1 OAI21X1_1707 ( .A(_1101__bF_buf16), .B(_1034_), .C(_1132_), .Y(_65_) );
OAI21X1 OAI21X1_1708 ( .A(_1100__bF_buf7_bF_buf2), .B(_1031__bF_buf68), .C(_3658__0_), .Y(_1133_) );
OAI21X1 OAI21X1_1709 ( .A(_1101__bF_buf6), .B(_1036_), .C(_1133_), .Y(_66_) );
NAND2X1 NAND2X1_714 ( .A(bundleLen_i[1]), .B(_612__bF_buf5), .Y(_1134_) );
INVX8 INVX8_7 ( .A(bundleLen_i[1]), .Y(_1135_) );
OAI21X1 OAI21X1_1710 ( .A(_1101__bF_buf14), .B(_1135__bF_buf2_bF_buf0), .C(_3659__31_), .Y(_1136_) );
OAI21X1 OAI21X1_1711 ( .A(_1038_), .B(_1134__bF_buf2), .C(_1136_), .Y(_67_) );
OAI21X1 OAI21X1_1712 ( .A(_1101__bF_buf47), .B(_1135__bF_buf1_bF_buf1), .C(_3659__30_), .Y(_1137_) );
OAI21X1 OAI21X1_1713 ( .A(_1041_), .B(_1134__bF_buf14), .C(_1137_), .Y(_68_) );
OAI21X1 OAI21X1_1714 ( .A(_1101__bF_buf42), .B(_1135__bF_buf11), .C(_3659__29_), .Y(_1138_) );
OAI21X1 OAI21X1_1715 ( .A(_1043_), .B(_1134__bF_buf10), .C(_1138_), .Y(_69_) );
OAI21X1 OAI21X1_1716 ( .A(_1101__bF_buf50), .B(_1135__bF_buf14_bF_buf2), .C(_3659__28_), .Y(_1139_) );
OAI21X1 OAI21X1_1717 ( .A(_1045_), .B(_1134__bF_buf5), .C(_1139_), .Y(_70_) );
OAI21X1 OAI21X1_1718 ( .A(_1101__bF_buf45), .B(_1135__bF_buf13_bF_buf2), .C(_3659__27_), .Y(_1140_) );
OAI21X1 OAI21X1_1719 ( .A(_1047_), .B(_1134__bF_buf1), .C(_1140_), .Y(_71_) );
OAI21X1 OAI21X1_1720 ( .A(_1101__bF_buf40), .B(_1135__bF_buf12_bF_buf1), .C(_3659__26_), .Y(_1141_) );
OAI21X1 OAI21X1_1721 ( .A(_1049_), .B(_1134__bF_buf0), .C(_1141_), .Y(_72_) );
OAI21X1 OAI21X1_1722 ( .A(_1101__bF_buf6), .B(_1135__bF_buf11_bF_buf1), .C(_3659__25_), .Y(_1142_) );
OAI21X1 OAI21X1_1723 ( .A(_1051_), .B(_1134__bF_buf1), .C(_1142_), .Y(_73_) );
OAI21X1 OAI21X1_1724 ( .A(_1101__bF_buf31), .B(_1135__bF_buf10_bF_buf1), .C(_3659__24_), .Y(_1143_) );
OAI21X1 OAI21X1_1725 ( .A(_1053_), .B(_1134__bF_buf11), .C(_1143_), .Y(_74_) );
OAI21X1 OAI21X1_1726 ( .A(_1101__bF_buf56), .B(_1135__bF_buf9_bF_buf2), .C(_3659__23_), .Y(_1144_) );
OAI21X1 OAI21X1_1727 ( .A(_1055_), .B(_1134__bF_buf10), .C(_1144_), .Y(_75_) );
OAI21X1 OAI21X1_1728 ( .A(_1101__bF_buf1), .B(_1135__bF_buf8_bF_buf3), .C(_3659__22_), .Y(_1145_) );
OAI21X1 OAI21X1_1729 ( .A(_1057_), .B(_1134__bF_buf2), .C(_1145_), .Y(_76_) );
OAI21X1 OAI21X1_1730 ( .A(_1101__bF_buf42), .B(_1135__bF_buf7_bF_buf1), .C(_3659__21_), .Y(_1146_) );
OAI21X1 OAI21X1_1731 ( .A(_1059_), .B(_1134__bF_buf10), .C(_1146_), .Y(_77_) );
OAI21X1 OAI21X1_1732 ( .A(_1101__bF_buf28), .B(_1135__bF_buf6_bF_buf1), .C(_3659__20_), .Y(_1147_) );
OAI21X1 OAI21X1_1733 ( .A(_1061_), .B(_1134__bF_buf7), .C(_1147_), .Y(_78_) );
OAI21X1 OAI21X1_1734 ( .A(_1101__bF_buf3), .B(_1135__bF_buf5_bF_buf0), .C(_3659__19_), .Y(_1148_) );
OAI21X1 OAI21X1_1735 ( .A(_1063_), .B(_1134__bF_buf7), .C(_1148_), .Y(_79_) );
OAI21X1 OAI21X1_1736 ( .A(_1101__bF_buf41), .B(_1135__bF_buf4_bF_buf2), .C(_3659__18_), .Y(_1149_) );
OAI21X1 OAI21X1_1737 ( .A(_1065_), .B(_1134__bF_buf11), .C(_1149_), .Y(_80_) );
OAI21X1 OAI21X1_1738 ( .A(_1101__bF_buf51), .B(_1135__bF_buf3_bF_buf0), .C(_3659__17_), .Y(_1150_) );
OAI21X1 OAI21X1_1739 ( .A(_1067_), .B(_1134__bF_buf2), .C(_1150_), .Y(_81_) );
OAI21X1 OAI21X1_1740 ( .A(_1101__bF_buf9), .B(_1135__bF_buf2_bF_buf2), .C(_3659__16_), .Y(_1151_) );
OAI21X1 OAI21X1_1741 ( .A(_1069_), .B(_1134__bF_buf2), .C(_1151_), .Y(_82_) );
OAI21X1 OAI21X1_1742 ( .A(_1101__bF_buf53), .B(_1135__bF_buf1_bF_buf1), .C(_3659__15_), .Y(_1152_) );
OAI21X1 OAI21X1_1743 ( .A(_1071_), .B(_1134__bF_buf13), .C(_1152_), .Y(_83_) );
OAI21X1 OAI21X1_1744 ( .A(_1101__bF_buf13), .B(_1135__bF_buf10), .C(_3659__14_), .Y(_1153_) );
OAI21X1 OAI21X1_1745 ( .A(_1073_), .B(_1134__bF_buf2), .C(_1153_), .Y(_84_) );
OAI21X1 OAI21X1_1746 ( .A(_1101__bF_buf54), .B(_1135__bF_buf14_bF_buf1), .C(_3659__13_), .Y(_1154_) );
OAI21X1 OAI21X1_1747 ( .A(_1075_), .B(_1134__bF_buf7), .C(_1154_), .Y(_85_) );
OAI21X1 OAI21X1_1748 ( .A(_1101__bF_buf37), .B(_1135__bF_buf13_bF_buf1), .C(_3659__12_), .Y(_1155_) );
OAI21X1 OAI21X1_1749 ( .A(_1077_), .B(_1134__bF_buf3), .C(_1155_), .Y(_86_) );
OAI21X1 OAI21X1_1750 ( .A(_1101__bF_buf35), .B(_1135__bF_buf12_bF_buf1), .C(_3659__11_), .Y(_1156_) );
OAI21X1 OAI21X1_1751 ( .A(_1079_), .B(_1134__bF_buf6), .C(_1156_), .Y(_87_) );
OAI21X1 OAI21X1_1752 ( .A(_1101__bF_buf28), .B(_1135__bF_buf11_bF_buf0), .C(_3659__10_), .Y(_1157_) );
OAI21X1 OAI21X1_1753 ( .A(_1081_), .B(_1134__bF_buf7), .C(_1157_), .Y(_88_) );
OAI21X1 OAI21X1_1754 ( .A(_1101__bF_buf20), .B(_1135__bF_buf10_bF_buf1), .C(_3659__9_), .Y(_1158_) );
OAI21X1 OAI21X1_1755 ( .A(_1083_), .B(_1134__bF_buf11), .C(_1158_), .Y(_89_) );
OAI21X1 OAI21X1_1756 ( .A(_1101__bF_buf56), .B(_1135__bF_buf9_bF_buf2), .C(_3659__8_), .Y(_1159_) );
OAI21X1 OAI21X1_1757 ( .A(_1085_), .B(_1134__bF_buf10), .C(_1159_), .Y(_90_) );
OAI21X1 OAI21X1_1758 ( .A(_1101__bF_buf41), .B(_1135__bF_buf8_bF_buf3), .C(_3659__7_), .Y(_1160_) );
OAI21X1 OAI21X1_1759 ( .A(_1087_), .B(_1134__bF_buf11), .C(_1160_), .Y(_91_) );
OAI21X1 OAI21X1_1760 ( .A(_1101__bF_buf32), .B(_1135__bF_buf7_bF_buf0), .C(_3659__6_), .Y(_1161_) );
OAI21X1 OAI21X1_1761 ( .A(_1089_), .B(_1134__bF_buf8), .C(_1161_), .Y(_92_) );
OAI21X1 OAI21X1_1762 ( .A(_1101__bF_buf56), .B(_1135__bF_buf6_bF_buf3), .C(_3659__5_), .Y(_1162_) );
OAI21X1 OAI21X1_1763 ( .A(_1091_), .B(_1134__bF_buf10), .C(_1162_), .Y(_93_) );
OAI21X1 OAI21X1_1764 ( .A(_1101__bF_buf30), .B(_1135__bF_buf5_bF_buf2), .C(_3659__4_), .Y(_1163_) );
OAI21X1 OAI21X1_1765 ( .A(_1093_), .B(_1134__bF_buf12), .C(_1163_), .Y(_94_) );
OAI21X1 OAI21X1_1766 ( .A(_1101__bF_buf0), .B(_1135__bF_buf4_bF_buf0), .C(_3659__3_), .Y(_1164_) );
OAI21X1 OAI21X1_1767 ( .A(_1095_), .B(_1134__bF_buf13), .C(_1164_), .Y(_95_) );
OAI21X1 OAI21X1_1768 ( .A(_1101__bF_buf17), .B(_1135__bF_buf3_bF_buf0), .C(_3659__2_), .Y(_1165_) );
OAI21X1 OAI21X1_1769 ( .A(_1032_), .B(_1134__bF_buf6), .C(_1165_), .Y(_96_) );
OAI21X1 OAI21X1_1770 ( .A(_1101__bF_buf48), .B(_1135__bF_buf2_bF_buf1), .C(_3659__1_), .Y(_1166_) );
OAI21X1 OAI21X1_1771 ( .A(_1034_), .B(_1134__bF_buf4), .C(_1166_), .Y(_97_) );
OAI21X1 OAI21X1_1772 ( .A(_1101__bF_buf16), .B(_1135__bF_buf1_bF_buf0), .C(_3659__0_), .Y(_1167_) );
OAI21X1 OAI21X1_1773 ( .A(_1036_), .B(_1134__bF_buf1), .C(_1167_), .Y(_98_) );
INVX2 INVX2_146 ( .A(bundleTid_i[63]), .Y(_1168_) );
NAND2X1 NAND2X1_715 ( .A(_3660__63_), .B(_1031__bF_buf9), .Y(_1169_) );
OAI21X1 OAI21X1_1774 ( .A(_1031__bF_buf54), .B(_1168_), .C(_1169_), .Y(_99_) );
INVX2 INVX2_147 ( .A(bundleTid_i[62]), .Y(_1170_) );
NAND2X1 NAND2X1_716 ( .A(_3660__62_), .B(_1031__bF_buf45), .Y(_1171_) );
OAI21X1 OAI21X1_1775 ( .A(_1031__bF_buf45), .B(_1170_), .C(_1171_), .Y(_100_) );
INVX2 INVX2_148 ( .A(bundleTid_i[61]), .Y(_1172_) );
NAND2X1 NAND2X1_717 ( .A(_3660__61_), .B(_1031__bF_buf15), .Y(_1173_) );
OAI21X1 OAI21X1_1776 ( .A(_1031__bF_buf51), .B(_1172_), .C(_1173_), .Y(_101_) );
INVX2 INVX2_149 ( .A(bundleTid_i[60]), .Y(_1174_) );
NAND2X1 NAND2X1_718 ( .A(_3660__60_), .B(_1031__bF_buf23), .Y(_1175_) );
OAI21X1 OAI21X1_1777 ( .A(_1031__bF_buf23), .B(_1174_), .C(_1175_), .Y(_102_) );
INVX2 INVX2_150 ( .A(bundleTid_i[59]), .Y(_1176_) );
NAND2X1 NAND2X1_719 ( .A(_3660__59_), .B(_1031__bF_buf3), .Y(_1177_) );
OAI21X1 OAI21X1_1778 ( .A(_1031__bF_buf3), .B(_1176_), .C(_1177_), .Y(_103_) );
INVX2 INVX2_151 ( .A(bundleTid_i[58]), .Y(_1178_) );
NAND2X1 NAND2X1_720 ( .A(_3660__58_), .B(_1031__bF_buf14), .Y(_1179_) );
OAI21X1 OAI21X1_1779 ( .A(_1031__bF_buf14), .B(_1178_), .C(_1179_), .Y(_104_) );
INVX2 INVX2_152 ( .A(bundleTid_i[57]), .Y(_1180_) );
NAND2X1 NAND2X1_721 ( .A(_3660__57_), .B(_1031__bF_buf44), .Y(_1181_) );
OAI21X1 OAI21X1_1780 ( .A(_1031__bF_buf44), .B(_1180_), .C(_1181_), .Y(_105_) );
INVX2 INVX2_153 ( .A(bundleTid_i[56]), .Y(_1182_) );
NAND2X1 NAND2X1_722 ( .A(_3660__56_), .B(_1031__bF_buf40), .Y(_1183_) );
OAI21X1 OAI21X1_1781 ( .A(_1031__bF_buf40), .B(_1182_), .C(_1183_), .Y(_106_) );
INVX2 INVX2_154 ( .A(bundleTid_i[55]), .Y(_1184_) );
NAND2X1 NAND2X1_723 ( .A(_3660__55_), .B(_1031__bF_buf73), .Y(_1185_) );
OAI21X1 OAI21X1_1782 ( .A(_1031__bF_buf73), .B(_1184_), .C(_1185_), .Y(_107_) );
INVX2 INVX2_155 ( .A(bundleTid_i[54]), .Y(_1186_) );
NAND2X1 NAND2X1_724 ( .A(_3660__54_), .B(_1031__bF_buf10), .Y(_1187_) );
OAI21X1 OAI21X1_1783 ( .A(_1031__bF_buf10), .B(_1186_), .C(_1187_), .Y(_108_) );
INVX2 INVX2_156 ( .A(bundleTid_i[53]), .Y(_1188_) );
NAND2X1 NAND2X1_725 ( .A(_3660__53_), .B(_1031__bF_buf62), .Y(_1189_) );
OAI21X1 OAI21X1_1784 ( .A(_1031__bF_buf62), .B(_1188_), .C(_1189_), .Y(_109_) );
INVX2 INVX2_157 ( .A(bundleTid_i[52]), .Y(_1190_) );
NAND2X1 NAND2X1_726 ( .A(_3660__52_), .B(_1031__bF_buf25), .Y(_1191_) );
OAI21X1 OAI21X1_1785 ( .A(_1031__bF_buf25), .B(_1190_), .C(_1191_), .Y(_110_) );
INVX2 INVX2_158 ( .A(bundleTid_i[51]), .Y(_1192_) );
NAND2X1 NAND2X1_727 ( .A(_3660__51_), .B(_1031__bF_buf66), .Y(_1193_) );
OAI21X1 OAI21X1_1786 ( .A(_1031__bF_buf66), .B(_1192_), .C(_1193_), .Y(_111_) );
INVX2 INVX2_159 ( .A(bundleTid_i[50]), .Y(_1194_) );
NAND2X1 NAND2X1_728 ( .A(_3660__50_), .B(_1031__bF_buf68), .Y(_1195_) );
OAI21X1 OAI21X1_1787 ( .A(_1031__bF_buf68), .B(_1194_), .C(_1195_), .Y(_112_) );
INVX2 INVX2_160 ( .A(bundleTid_i[49]), .Y(_1196_) );
NAND2X1 NAND2X1_729 ( .A(_3660__49_), .B(_1031__bF_buf47), .Y(_1197_) );
OAI21X1 OAI21X1_1788 ( .A(_1031__bF_buf8), .B(_1196_), .C(_1197_), .Y(_113_) );
INVX2 INVX2_161 ( .A(bundleTid_i[48]), .Y(_1198_) );
NAND2X1 NAND2X1_730 ( .A(_3660__48_), .B(_1031__bF_buf20), .Y(_1199_) );
OAI21X1 OAI21X1_1789 ( .A(_1031__bF_buf20), .B(_1198_), .C(_1199_), .Y(_114_) );
INVX2 INVX2_162 ( .A(bundleTid_i[47]), .Y(_1200_) );
NAND2X1 NAND2X1_731 ( .A(_3660__47_), .B(_1031__bF_buf54), .Y(_1201_) );
OAI21X1 OAI21X1_1790 ( .A(_1031__bF_buf54), .B(_1200_), .C(_1201_), .Y(_115_) );
INVX2 INVX2_163 ( .A(bundleTid_i[46]), .Y(_1202_) );
NAND2X1 NAND2X1_732 ( .A(_3660__46_), .B(_1031__bF_buf3), .Y(_1203_) );
OAI21X1 OAI21X1_1791 ( .A(_1031__bF_buf3), .B(_1202_), .C(_1203_), .Y(_116_) );
INVX2 INVX2_164 ( .A(bundleTid_i[45]), .Y(_1204_) );
NAND2X1 NAND2X1_733 ( .A(_3660__45_), .B(_1031__bF_buf70), .Y(_1205_) );
OAI21X1 OAI21X1_1792 ( .A(_1031__bF_buf70), .B(_1204_), .C(_1205_), .Y(_117_) );
INVX2 INVX2_165 ( .A(bundleTid_i[44]), .Y(_1206_) );
NAND2X1 NAND2X1_734 ( .A(_3660__44_), .B(_1031__bF_buf35), .Y(_1207_) );
OAI21X1 OAI21X1_1793 ( .A(_1031__bF_buf35), .B(_1206_), .C(_1207_), .Y(_118_) );
INVX2 INVX2_166 ( .A(bundleTid_i[43]), .Y(_1208_) );
NAND2X1 NAND2X1_735 ( .A(_3660__43_), .B(_1031__bF_buf5), .Y(_1209_) );
OAI21X1 OAI21X1_1794 ( .A(_1031__bF_buf5), .B(_1208_), .C(_1209_), .Y(_119_) );
INVX2 INVX2_167 ( .A(bundleTid_i[42]), .Y(_1210_) );
NAND2X1 NAND2X1_736 ( .A(_3660__42_), .B(_1031__bF_buf59), .Y(_1211_) );
OAI21X1 OAI21X1_1795 ( .A(_1031__bF_buf20), .B(_1210_), .C(_1211_), .Y(_120_) );
INVX2 INVX2_168 ( .A(bundleTid_i[41]), .Y(_1212_) );
NAND2X1 NAND2X1_737 ( .A(_3660__41_), .B(_1031__bF_buf13), .Y(_1213_) );
OAI21X1 OAI21X1_1796 ( .A(_1031__bF_buf13), .B(_1212_), .C(_1213_), .Y(_121_) );
INVX2 INVX2_169 ( .A(bundleTid_i[40]), .Y(_1214_) );
NAND2X1 NAND2X1_738 ( .A(_3660__40_), .B(_1031__bF_buf13), .Y(_1215_) );
OAI21X1 OAI21X1_1797 ( .A(_1031__bF_buf13), .B(_1214_), .C(_1215_), .Y(_122_) );
INVX2 INVX2_170 ( .A(bundleTid_i[39]), .Y(_1216_) );
NAND2X1 NAND2X1_739 ( .A(_3660__39_), .B(_1031__bF_buf27), .Y(_1217_) );
OAI21X1 OAI21X1_1798 ( .A(_1031__bF_buf27), .B(_1216_), .C(_1217_), .Y(_123_) );
INVX2 INVX2_171 ( .A(bundleTid_i[38]), .Y(_1218_) );
NAND2X1 NAND2X1_740 ( .A(_3660__38_), .B(_1031__bF_buf25), .Y(_1219_) );
OAI21X1 OAI21X1_1799 ( .A(_1031__bF_buf25), .B(_1218_), .C(_1219_), .Y(_124_) );
INVX2 INVX2_172 ( .A(bundleTid_i[37]), .Y(_1220_) );
NAND2X1 NAND2X1_741 ( .A(_3660__37_), .B(_1031__bF_buf25), .Y(_1221_) );
OAI21X1 OAI21X1_1800 ( .A(_1031__bF_buf25), .B(_1220_), .C(_1221_), .Y(_125_) );
INVX2 INVX2_173 ( .A(bundleTid_i[36]), .Y(_1222_) );
NAND2X1 NAND2X1_742 ( .A(_3660__36_), .B(_1031__bF_buf56), .Y(_1223_) );
OAI21X1 OAI21X1_1801 ( .A(_1031__bF_buf56), .B(_1222_), .C(_1223_), .Y(_126_) );
INVX2 INVX2_174 ( .A(bundleTid_i[35]), .Y(_1224_) );
NAND2X1 NAND2X1_743 ( .A(_3660__35_), .B(_1031__bF_buf45), .Y(_1225_) );
OAI21X1 OAI21X1_1802 ( .A(_1031__bF_buf45), .B(_1224_), .C(_1225_), .Y(_127_) );
INVX2 INVX2_175 ( .A(bundleTid_i[34]), .Y(_1226_) );
NAND2X1 NAND2X1_744 ( .A(_3660__34_), .B(_1031__bF_buf4), .Y(_1227_) );
OAI21X1 OAI21X1_1803 ( .A(_1031__bF_buf4), .B(_1226_), .C(_1227_), .Y(_128_) );
INVX2 INVX2_176 ( .A(bundleTid_i[33]), .Y(_1228_) );
NAND2X1 NAND2X1_745 ( .A(_3660__33_), .B(_1031__bF_buf52), .Y(_1229_) );
OAI21X1 OAI21X1_1804 ( .A(_1031__bF_buf52), .B(_1228_), .C(_1229_), .Y(_129_) );
INVX2 INVX2_177 ( .A(bundleTid_i[32]), .Y(_1230_) );
NAND2X1 NAND2X1_746 ( .A(_3660__32_), .B(_1031__bF_buf22), .Y(_1231_) );
OAI21X1 OAI21X1_1805 ( .A(_1031__bF_buf22), .B(_1230_), .C(_1231_), .Y(_130_) );
INVX2 INVX2_178 ( .A(bundleTid_i[31]), .Y(_1232_) );
NAND2X1 NAND2X1_747 ( .A(_3660__31_), .B(_1031__bF_buf68), .Y(_1233_) );
OAI21X1 OAI21X1_1806 ( .A(_1031__bF_buf68), .B(_1232_), .C(_1233_), .Y(_131_) );
INVX2 INVX2_179 ( .A(bundleTid_i[30]), .Y(_1234_) );
NAND2X1 NAND2X1_748 ( .A(_3660__30_), .B(_1031__bF_buf59), .Y(_1235_) );
OAI21X1 OAI21X1_1807 ( .A(_1031__bF_buf59), .B(_1234_), .C(_1235_), .Y(_132_) );
INVX2 INVX2_180 ( .A(bundleTid_i[29]), .Y(_1236_) );
NAND2X1 NAND2X1_749 ( .A(_3660__29_), .B(_1031__bF_buf72), .Y(_1237_) );
OAI21X1 OAI21X1_1808 ( .A(_1031__bF_buf72), .B(_1236_), .C(_1237_), .Y(_133_) );
INVX2 INVX2_181 ( .A(bundleTid_i[28]), .Y(_1238_) );
NAND2X1 NAND2X1_750 ( .A(_3660__28_), .B(_1031__bF_buf12), .Y(_1239_) );
OAI21X1 OAI21X1_1809 ( .A(_1031__bF_buf12), .B(_1238_), .C(_1239_), .Y(_134_) );
INVX2 INVX2_182 ( .A(bundleTid_i[27]), .Y(_1240_) );
NAND2X1 NAND2X1_751 ( .A(_3660__27_), .B(_1031__bF_buf77), .Y(_1241_) );
OAI21X1 OAI21X1_1810 ( .A(_1031__bF_buf77), .B(_1240_), .C(_1241_), .Y(_135_) );
INVX2 INVX2_183 ( .A(bundleTid_i[26]), .Y(_1242_) );
NAND2X1 NAND2X1_752 ( .A(_3660__26_), .B(_1031__bF_buf59), .Y(_1243_) );
OAI21X1 OAI21X1_1811 ( .A(_1031__bF_buf36), .B(_1242_), .C(_1243_), .Y(_136_) );
INVX2 INVX2_184 ( .A(bundleTid_i[25]), .Y(_1244_) );
NAND2X1 NAND2X1_753 ( .A(_3660__25_), .B(_1031__bF_buf75), .Y(_1245_) );
OAI21X1 OAI21X1_1812 ( .A(_1031__bF_buf66), .B(_1244_), .C(_1245_), .Y(_137_) );
INVX2 INVX2_185 ( .A(bundleTid_i[24]), .Y(_1246_) );
NAND2X1 NAND2X1_754 ( .A(_3660__24_), .B(_1031__bF_buf13), .Y(_1247_) );
OAI21X1 OAI21X1_1813 ( .A(_1031__bF_buf13), .B(_1246_), .C(_1247_), .Y(_138_) );
INVX2 INVX2_186 ( .A(bundleTid_i[23]), .Y(_1248_) );
NAND2X1 NAND2X1_755 ( .A(_3660__23_), .B(_1031__bF_buf34), .Y(_1249_) );
OAI21X1 OAI21X1_1814 ( .A(_1031__bF_buf74), .B(_1248_), .C(_1249_), .Y(_139_) );
INVX2 INVX2_187 ( .A(bundleTid_i[22]), .Y(_1250_) );
NAND2X1 NAND2X1_756 ( .A(_3660__22_), .B(_1031__bF_buf45), .Y(_1251_) );
OAI21X1 OAI21X1_1815 ( .A(_1031__bF_buf24), .B(_1250_), .C(_1251_), .Y(_140_) );
INVX2 INVX2_188 ( .A(bundleTid_i[21]), .Y(_1252_) );
NAND2X1 NAND2X1_757 ( .A(_3660__21_), .B(_1031__bF_buf4), .Y(_1253_) );
OAI21X1 OAI21X1_1816 ( .A(_1031__bF_buf4), .B(_1252_), .C(_1253_), .Y(_141_) );
INVX2 INVX2_189 ( .A(bundleTid_i[20]), .Y(_1254_) );
NAND2X1 NAND2X1_758 ( .A(_3660__20_), .B(_1031__bF_buf75), .Y(_1255_) );
OAI21X1 OAI21X1_1817 ( .A(_1031__bF_buf75), .B(_1254_), .C(_1255_), .Y(_142_) );
INVX2 INVX2_190 ( .A(bundleTid_i[19]), .Y(_1256_) );
NAND2X1 NAND2X1_759 ( .A(_3660__19_), .B(_1031__bF_buf52), .Y(_1257_) );
OAI21X1 OAI21X1_1818 ( .A(_1031__bF_buf52), .B(_1256_), .C(_1257_), .Y(_143_) );
INVX2 INVX2_191 ( .A(bundleTid_i[18]), .Y(_1258_) );
NAND2X1 NAND2X1_760 ( .A(_3660__18_), .B(_1031__bF_buf72), .Y(_1259_) );
OAI21X1 OAI21X1_1819 ( .A(_1031__bF_buf72), .B(_1258_), .C(_1259_), .Y(_144_) );
INVX2 INVX2_192 ( .A(bundleTid_i[17]), .Y(_1260_) );
NAND2X1 NAND2X1_761 ( .A(_3660__17_), .B(_1031__bF_buf61), .Y(_1261_) );
OAI21X1 OAI21X1_1820 ( .A(_1031__bF_buf61), .B(_1260_), .C(_1261_), .Y(_145_) );
INVX2 INVX2_193 ( .A(bundleTid_i[16]), .Y(_1262_) );
NAND2X1 NAND2X1_762 ( .A(_3660__16_), .B(_1031__bF_buf52), .Y(_1263_) );
OAI21X1 OAI21X1_1821 ( .A(_1031__bF_buf27), .B(_1262_), .C(_1263_), .Y(_146_) );
INVX2 INVX2_194 ( .A(bundleTid_i[15]), .Y(_1264_) );
NAND2X1 NAND2X1_763 ( .A(_3660__15_), .B(_1031__bF_buf11), .Y(_1265_) );
OAI21X1 OAI21X1_1822 ( .A(_1031__bF_buf11), .B(_1264_), .C(_1265_), .Y(_147_) );
INVX2 INVX2_195 ( .A(bundleTid_i[14]), .Y(_1266_) );
NAND2X1 NAND2X1_764 ( .A(_3660__14_), .B(_1031__bF_buf75), .Y(_1267_) );
OAI21X1 OAI21X1_1823 ( .A(_1031__bF_buf75), .B(_1266_), .C(_1267_), .Y(_148_) );
INVX2 INVX2_196 ( .A(bundleTid_i[13]), .Y(_1268_) );
NAND2X1 NAND2X1_765 ( .A(_3660__13_), .B(_1031__bF_buf29), .Y(_1269_) );
OAI21X1 OAI21X1_1824 ( .A(_1031__bF_buf29), .B(_1268_), .C(_1269_), .Y(_149_) );
INVX2 INVX2_197 ( .A(bundleTid_i[12]), .Y(_1270_) );
NAND2X1 NAND2X1_766 ( .A(_3660__12_), .B(_1031__bF_buf40), .Y(_1271_) );
OAI21X1 OAI21X1_1825 ( .A(_1031__bF_buf40), .B(_1270_), .C(_1271_), .Y(_150_) );
INVX2 INVX2_198 ( .A(bundleTid_i[11]), .Y(_1272_) );
NAND2X1 NAND2X1_767 ( .A(_3660__11_), .B(_1031__bF_buf55), .Y(_1273_) );
OAI21X1 OAI21X1_1826 ( .A(_1031__bF_buf55), .B(_1272_), .C(_1273_), .Y(_151_) );
INVX2 INVX2_199 ( .A(bundleTid_i[10]), .Y(_1274_) );
NAND2X1 NAND2X1_768 ( .A(_3660__10_), .B(_1031__bF_buf8), .Y(_1275_) );
OAI21X1 OAI21X1_1827 ( .A(_1031__bF_buf8), .B(_1274_), .C(_1275_), .Y(_152_) );
INVX2 INVX2_200 ( .A(bundleTid_i[9]), .Y(_1276_) );
NAND2X1 NAND2X1_769 ( .A(_3660__9_), .B(_1031__bF_buf36), .Y(_1277_) );
OAI21X1 OAI21X1_1828 ( .A(_1031__bF_buf36), .B(_1276_), .C(_1277_), .Y(_153_) );
INVX2 INVX2_201 ( .A(bundleTid_i[8]), .Y(_1278_) );
NAND2X1 NAND2X1_770 ( .A(_3660__8_), .B(_1031__bF_buf21), .Y(_1279_) );
OAI21X1 OAI21X1_1829 ( .A(_1031__bF_buf21), .B(_1278_), .C(_1279_), .Y(_154_) );
INVX2 INVX2_202 ( .A(bundleTid_i[7]), .Y(_1280_) );
NAND2X1 NAND2X1_771 ( .A(_3660__7_), .B(_1031__bF_buf27), .Y(_1281_) );
OAI21X1 OAI21X1_1830 ( .A(_1031__bF_buf27), .B(_1280_), .C(_1281_), .Y(_155_) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock_i_bF_buf64), .D(_0_), .Q(_3656__2_) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock_i_bF_buf10), .D(_1_), .Q(_3656__1_) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock_i_bF_buf36), .D(_2_), .Q(_3656__0_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock_i_bF_buf16), .D(_3_), .Q(_3657__31_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock_i_bF_buf37), .D(_4_), .Q(_3657__30_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(clock_i_bF_buf3), .D(_5_), .Q(_3657__29_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(clock_i_bF_buf51), .D(_6_), .Q(_3657__28_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(clock_i_bF_buf15), .D(_7_), .Q(_3657__27_) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(clock_i_bF_buf44), .D(_8_), .Q(_3657__26_) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(clock_i_bF_buf61), .D(_9_), .Q(_3657__25_) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(clock_i_bF_buf9), .D(_10_), .Q(_3657__24_) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(clock_i_bF_buf60), .D(_11_), .Q(_3657__23_) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(clock_i_bF_buf45), .D(_12_), .Q(_3657__22_) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(clock_i_bF_buf60), .D(_13_), .Q(_3657__21_) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(clock_i_bF_buf41), .D(_14_), .Q(_3657__20_) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(clock_i_bF_buf15), .D(_15_), .Q(_3657__19_) );
DFFPOSX1 DFFPOSX1_17 ( .CLK(clock_i_bF_buf53), .D(_16_), .Q(_3657__18_) );
DFFPOSX1 DFFPOSX1_18 ( .CLK(clock_i_bF_buf16), .D(_17_), .Q(_3657__17_) );
DFFPOSX1 DFFPOSX1_19 ( .CLK(clock_i_bF_buf45), .D(_18_), .Q(_3657__16_) );
DFFPOSX1 DFFPOSX1_20 ( .CLK(clock_i_bF_buf91), .D(_19_), .Q(_3657__15_) );
DFFPOSX1 DFFPOSX1_21 ( .CLK(clock_i_bF_buf7), .D(_20_), .Q(_3657__14_) );
DFFPOSX1 DFFPOSX1_22 ( .CLK(clock_i_bF_buf29), .D(_21_), .Q(_3657__13_) );
DFFPOSX1 DFFPOSX1_23 ( .CLK(clock_i_bF_buf10), .D(_22_), .Q(_3657__12_) );
DFFPOSX1 DFFPOSX1_24 ( .CLK(clock_i_bF_buf35), .D(_23_), .Q(_3657__11_) );
DFFPOSX1 DFFPOSX1_25 ( .CLK(clock_i_bF_buf38), .D(_24_), .Q(_3657__10_) );
DFFPOSX1 DFFPOSX1_26 ( .CLK(clock_i_bF_buf86), .D(_25_), .Q(_3657__9_) );
DFFPOSX1 DFFPOSX1_27 ( .CLK(clock_i_bF_buf70), .D(_26_), .Q(_3657__8_) );
DFFPOSX1 DFFPOSX1_28 ( .CLK(clock_i_bF_buf50), .D(_27_), .Q(_3657__7_) );
DFFPOSX1 DFFPOSX1_29 ( .CLK(clock_i_bF_buf55), .D(_28_), .Q(_3657__6_) );
DFFPOSX1 DFFPOSX1_30 ( .CLK(clock_i_bF_buf3), .D(_29_), .Q(_3657__5_) );
DFFPOSX1 DFFPOSX1_31 ( .CLK(clock_i_bF_buf100), .D(_30_), .Q(_3657__4_) );
DFFPOSX1 DFFPOSX1_32 ( .CLK(clock_i_bF_buf1), .D(_31_), .Q(_3657__3_) );
DFFPOSX1 DFFPOSX1_33 ( .CLK(clock_i_bF_buf64), .D(_32_), .Q(_3657__2_) );
DFFPOSX1 DFFPOSX1_34 ( .CLK(clock_i_bF_buf27), .D(_33_), .Q(_3657__1_) );
DFFPOSX1 DFFPOSX1_35 ( .CLK(clock_i_bF_buf61), .D(_34_), .Q(_3657__0_) );
DFFPOSX1 DFFPOSX1_36 ( .CLK(clock_i_bF_buf16), .D(_35_), .Q(_3658__31_) );
DFFPOSX1 DFFPOSX1_37 ( .CLK(clock_i_bF_buf37), .D(_36_), .Q(_3658__30_) );
DFFPOSX1 DFFPOSX1_38 ( .CLK(clock_i_bF_buf3), .D(_37_), .Q(_3658__29_) );
DFFPOSX1 DFFPOSX1_39 ( .CLK(clock_i_bF_buf95), .D(_38_), .Q(_3658__28_) );
DFFPOSX1 DFFPOSX1_40 ( .CLK(clock_i_bF_buf15), .D(_39_), .Q(_3658__27_) );
DFFPOSX1 DFFPOSX1_41 ( .CLK(clock_i_bF_buf44), .D(_40_), .Q(_3658__26_) );
DFFPOSX1 DFFPOSX1_42 ( .CLK(clock_i_bF_buf61), .D(_41_), .Q(_3658__25_) );
DFFPOSX1 DFFPOSX1_43 ( .CLK(clock_i_bF_buf9), .D(_42_), .Q(_3658__24_) );
DFFPOSX1 DFFPOSX1_44 ( .CLK(clock_i_bF_buf60), .D(_43_), .Q(_3658__23_) );
DFFPOSX1 DFFPOSX1_45 ( .CLK(clock_i_bF_buf60), .D(_44_), .Q(_3658__22_) );
DFFPOSX1 DFFPOSX1_46 ( .CLK(clock_i_bF_buf94), .D(_45_), .Q(_3658__21_) );
DFFPOSX1 DFFPOSX1_47 ( .CLK(clock_i_bF_buf38), .D(_46_), .Q(_3658__20_) );
DFFPOSX1 DFFPOSX1_48 ( .CLK(clock_i_bF_buf15), .D(_47_), .Q(_3658__19_) );
DFFPOSX1 DFFPOSX1_49 ( .CLK(clock_i_bF_buf25), .D(_48_), .Q(_3658__18_) );
DFFPOSX1 DFFPOSX1_50 ( .CLK(clock_i_bF_buf77), .D(_49_), .Q(_3658__17_) );
DFFPOSX1 DFFPOSX1_51 ( .CLK(clock_i_bF_buf13), .D(_50_), .Q(_3658__16_) );
DFFPOSX1 DFFPOSX1_52 ( .CLK(clock_i_bF_buf71), .D(_51_), .Q(_3658__15_) );
DFFPOSX1 DFFPOSX1_53 ( .CLK(clock_i_bF_buf7), .D(_52_), .Q(_3658__14_) );
DFFPOSX1 DFFPOSX1_54 ( .CLK(clock_i_bF_buf24), .D(_53_), .Q(_3658__13_) );
DFFPOSX1 DFFPOSX1_55 ( .CLK(clock_i_bF_buf57), .D(_54_), .Q(_3658__12_) );
DFFPOSX1 DFFPOSX1_56 ( .CLK(clock_i_bF_buf35), .D(_55_), .Q(_3658__11_) );
DFFPOSX1 DFFPOSX1_57 ( .CLK(clock_i_bF_buf41), .D(_56_), .Q(_3658__10_) );
DFFPOSX1 DFFPOSX1_58 ( .CLK(clock_i_bF_buf86), .D(_57_), .Q(_3658__9_) );
DFFPOSX1 DFFPOSX1_59 ( .CLK(clock_i_bF_buf70), .D(_58_), .Q(_3658__8_) );
DFFPOSX1 DFFPOSX1_60 ( .CLK(clock_i_bF_buf55), .D(_59_), .Q(_3658__7_) );
DFFPOSX1 DFFPOSX1_61 ( .CLK(clock_i_bF_buf55), .D(_60_), .Q(_3658__6_) );
DFFPOSX1 DFFPOSX1_62 ( .CLK(clock_i_bF_buf94), .D(_61_), .Q(_3658__5_) );
DFFPOSX1 DFFPOSX1_63 ( .CLK(clock_i_bF_buf55), .D(_62_), .Q(_3658__4_) );
DFFPOSX1 DFFPOSX1_64 ( .CLK(clock_i_bF_buf80), .D(_63_), .Q(_3658__3_) );
DFFPOSX1 DFFPOSX1_65 ( .CLK(clock_i_bF_buf33), .D(_64_), .Q(_3658__2_) );
DFFPOSX1 DFFPOSX1_66 ( .CLK(clock_i_bF_buf27), .D(_65_), .Q(_3658__1_) );
DFFPOSX1 DFFPOSX1_67 ( .CLK(clock_i_bF_buf36), .D(_66_), .Q(_3658__0_) );
DFFPOSX1 DFFPOSX1_68 ( .CLK(clock_i_bF_buf77), .D(_67_), .Q(_3659__31_) );
DFFPOSX1 DFFPOSX1_69 ( .CLK(clock_i_bF_buf28), .D(_68_), .Q(_3659__30_) );
DFFPOSX1 DFFPOSX1_70 ( .CLK(clock_i_bF_buf94), .D(_69_), .Q(_3659__29_) );
DFFPOSX1 DFFPOSX1_71 ( .CLK(clock_i_bF_buf67), .D(_70_), .Q(_3659__28_) );
DFFPOSX1 DFFPOSX1_72 ( .CLK(clock_i_bF_buf15), .D(_71_), .Q(_3659__27_) );
DFFPOSX1 DFFPOSX1_73 ( .CLK(clock_i_bF_buf44), .D(_72_), .Q(_3659__26_) );
DFFPOSX1 DFFPOSX1_74 ( .CLK(clock_i_bF_buf46), .D(_73_), .Q(_3659__25_) );
DFFPOSX1 DFFPOSX1_75 ( .CLK(clock_i_bF_buf9), .D(_74_), .Q(_3659__24_) );
DFFPOSX1 DFFPOSX1_76 ( .CLK(clock_i_bF_buf85), .D(_75_), .Q(_3659__23_) );
DFFPOSX1 DFFPOSX1_77 ( .CLK(clock_i_bF_buf7), .D(_76_), .Q(_3659__22_) );
DFFPOSX1 DFFPOSX1_78 ( .CLK(clock_i_bF_buf94), .D(_77_), .Q(_3659__21_) );
DFFPOSX1 DFFPOSX1_79 ( .CLK(clock_i_bF_buf80), .D(_78_), .Q(_3659__20_) );
DFFPOSX1 DFFPOSX1_80 ( .CLK(clock_i_bF_buf57), .D(_79_), .Q(_3659__19_) );
DFFPOSX1 DFFPOSX1_81 ( .CLK(clock_i_bF_buf47), .D(_80_), .Q(_3659__18_) );
DFFPOSX1 DFFPOSX1_82 ( .CLK(clock_i_bF_buf16), .D(_81_), .Q(_3659__17_) );
DFFPOSX1 DFFPOSX1_83 ( .CLK(clock_i_bF_buf16), .D(_82_), .Q(_3659__16_) );
DFFPOSX1 DFFPOSX1_84 ( .CLK(clock_i_bF_buf1), .D(_83_), .Q(_3659__15_) );
DFFPOSX1 DFFPOSX1_85 ( .CLK(clock_i_bF_buf75), .D(_84_), .Q(_3659__14_) );
DFFPOSX1 DFFPOSX1_86 ( .CLK(clock_i_bF_buf29), .D(_85_), .Q(_3659__13_) );
DFFPOSX1 DFFPOSX1_87 ( .CLK(clock_i_bF_buf83), .D(_86_), .Q(_3659__12_) );
DFFPOSX1 DFFPOSX1_88 ( .CLK(clock_i_bF_buf62), .D(_87_), .Q(_3659__11_) );
DFFPOSX1 DFFPOSX1_89 ( .CLK(clock_i_bF_buf38), .D(_88_), .Q(_3659__10_) );
DFFPOSX1 DFFPOSX1_90 ( .CLK(clock_i_bF_buf86), .D(_89_), .Q(_3659__9_) );
DFFPOSX1 DFFPOSX1_91 ( .CLK(clock_i_bF_buf70), .D(_90_), .Q(_3659__8_) );
DFFPOSX1 DFFPOSX1_92 ( .CLK(clock_i_bF_buf99), .D(_91_), .Q(_3659__7_) );
DFFPOSX1 DFFPOSX1_93 ( .CLK(clock_i_bF_buf52), .D(_92_), .Q(_3659__6_) );
DFFPOSX1 DFFPOSX1_94 ( .CLK(clock_i_bF_buf3), .D(_93_), .Q(_3659__5_) );
DFFPOSX1 DFFPOSX1_95 ( .CLK(clock_i_bF_buf0), .D(_94_), .Q(_3659__4_) );
DFFPOSX1 DFFPOSX1_96 ( .CLK(clock_i_bF_buf38), .D(_95_), .Q(_3659__3_) );
DFFPOSX1 DFFPOSX1_97 ( .CLK(clock_i_bF_buf76), .D(_96_), .Q(_3659__2_) );
DFFPOSX1 DFFPOSX1_98 ( .CLK(clock_i_bF_buf96), .D(_97_), .Q(_3659__1_) );
DFFPOSX1 DFFPOSX1_99 ( .CLK(clock_i_bF_buf36), .D(_98_), .Q(_3659__0_) );
DFFPOSX1 DFFPOSX1_100 ( .CLK(clock_i_bF_buf55), .D(_99_), .Q(_3660__63_) );
DFFPOSX1 DFFPOSX1_101 ( .CLK(clock_i_bF_buf31), .D(_100_), .Q(_3660__62_) );
DFFPOSX1 DFFPOSX1_102 ( .CLK(clock_i_bF_buf10), .D(_101_), .Q(_3660__61_) );
DFFPOSX1 DFFPOSX1_103 ( .CLK(clock_i_bF_buf8), .D(_102_), .Q(_3660__60_) );
DFFPOSX1 DFFPOSX1_104 ( .CLK(clock_i_bF_buf43), .D(_103_), .Q(_3660__59_) );
DFFPOSX1 DFFPOSX1_105 ( .CLK(clock_i_bF_buf31), .D(_104_), .Q(_3660__58_) );
DFFPOSX1 DFFPOSX1_106 ( .CLK(clock_i_bF_buf53), .D(_105_), .Q(_3660__57_) );
DFFPOSX1 DFFPOSX1_107 ( .CLK(clock_i_bF_buf76), .D(_106_), .Q(_3660__56_) );
DFFPOSX1 DFFPOSX1_108 ( .CLK(clock_i_bF_buf46), .D(_107_), .Q(_3660__55_) );
DFFPOSX1 DFFPOSX1_109 ( .CLK(clock_i_bF_buf101), .D(_108_), .Q(_3660__54_) );
DFFPOSX1 DFFPOSX1_110 ( .CLK(clock_i_bF_buf100), .D(_109_), .Q(_3660__53_) );
DFFPOSX1 DFFPOSX1_111 ( .CLK(clock_i_bF_buf88), .D(_110_), .Q(_3660__52_) );
DFFPOSX1 DFFPOSX1_112 ( .CLK(clock_i_bF_buf85), .D(_111_), .Q(_3660__51_) );
DFFPOSX1 DFFPOSX1_113 ( .CLK(clock_i_bF_buf46), .D(_112_), .Q(_3660__50_) );
DFFPOSX1 DFFPOSX1_114 ( .CLK(clock_i_bF_buf77), .D(_113_), .Q(_3660__49_) );
DFFPOSX1 DFFPOSX1_115 ( .CLK(clock_i_bF_buf63), .D(_114_), .Q(_3660__48_) );
DFFPOSX1 DFFPOSX1_116 ( .CLK(clock_i_bF_buf55), .D(_115_), .Q(_3660__47_) );
DFFPOSX1 DFFPOSX1_117 ( .CLK(clock_i_bF_buf43), .D(_116_), .Q(_3660__46_) );
DFFPOSX1 DFFPOSX1_118 ( .CLK(clock_i_bF_buf13), .D(_117_), .Q(_3660__45_) );
DFFPOSX1 DFFPOSX1_119 ( .CLK(clock_i_bF_buf90), .D(_118_), .Q(_3660__44_) );
DFFPOSX1 DFFPOSX1_120 ( .CLK(clock_i_bF_buf87), .D(_119_), .Q(_3660__43_) );
DFFPOSX1 DFFPOSX1_121 ( .CLK(clock_i_bF_buf63), .D(_120_), .Q(_3660__42_) );
DFFPOSX1 DFFPOSX1_122 ( .CLK(clock_i_bF_buf35), .D(_121_), .Q(_3660__41_) );
DFFPOSX1 DFFPOSX1_123 ( .CLK(clock_i_bF_buf35), .D(_122_), .Q(_3660__40_) );
DFFPOSX1 DFFPOSX1_124 ( .CLK(clock_i_bF_buf9), .D(_123_), .Q(_3660__39_) );
DFFPOSX1 DFFPOSX1_125 ( .CLK(clock_i_bF_buf99), .D(_124_), .Q(_3660__38_) );
DFFPOSX1 DFFPOSX1_126 ( .CLK(clock_i_bF_buf99), .D(_125_), .Q(_3660__37_) );
DFFPOSX1 DFFPOSX1_127 ( .CLK(clock_i_bF_buf70), .D(_126_), .Q(_3660__36_) );
DFFPOSX1 DFFPOSX1_128 ( .CLK(clock_i_bF_buf21), .D(_127_), .Q(_3660__35_) );
DFFPOSX1 DFFPOSX1_129 ( .CLK(clock_i_bF_buf40), .D(_128_), .Q(_3660__34_) );
DFFPOSX1 DFFPOSX1_130 ( .CLK(clock_i_bF_buf9), .D(_129_), .Q(_3660__33_) );
DFFPOSX1 DFFPOSX1_131 ( .CLK(clock_i_bF_buf24), .D(_130_), .Q(_3660__32_) );
DFFPOSX1 DFFPOSX1_132 ( .CLK(clock_i_bF_buf36), .D(_131_), .Q(_3660__31_) );
DFFPOSX1 DFFPOSX1_133 ( .CLK(clock_i_bF_buf63), .D(_132_), .Q(_3660__30_) );
DFFPOSX1 DFFPOSX1_134 ( .CLK(clock_i_bF_buf91), .D(_133_), .Q(_3660__29_) );
DFFPOSX1 DFFPOSX1_135 ( .CLK(clock_i_bF_buf29), .D(_134_), .Q(_3660__28_) );
DFFPOSX1 DFFPOSX1_136 ( .CLK(clock_i_bF_buf86), .D(_135_), .Q(_3660__27_) );
DFFPOSX1 DFFPOSX1_137 ( .CLK(clock_i_bF_buf63), .D(_136_), .Q(_3660__26_) );
DFFPOSX1 DFFPOSX1_138 ( .CLK(clock_i_bF_buf16), .D(_137_), .Q(_3660__25_) );
DFFPOSX1 DFFPOSX1_139 ( .CLK(clock_i_bF_buf35), .D(_138_), .Q(_3660__24_) );
DFFPOSX1 DFFPOSX1_140 ( .CLK(clock_i_bF_buf100), .D(_139_), .Q(_3660__23_) );
DFFPOSX1 DFFPOSX1_141 ( .CLK(clock_i_bF_buf21), .D(_140_), .Q(_3660__22_) );
DFFPOSX1 DFFPOSX1_142 ( .CLK(clock_i_bF_buf49), .D(_141_), .Q(_3660__21_) );
DFFPOSX1 DFFPOSX1_143 ( .CLK(clock_i_bF_buf94), .D(_142_), .Q(_3660__20_) );
DFFPOSX1 DFFPOSX1_144 ( .CLK(clock_i_bF_buf95), .D(_143_), .Q(_3660__19_) );
DFFPOSX1 DFFPOSX1_145 ( .CLK(clock_i_bF_buf91), .D(_144_), .Q(_3660__18_) );
DFFPOSX1 DFFPOSX1_146 ( .CLK(clock_i_bF_buf61), .D(_145_), .Q(_3660__17_) );
DFFPOSX1 DFFPOSX1_147 ( .CLK(clock_i_bF_buf86), .D(_146_), .Q(_3660__16_) );
DFFPOSX1 DFFPOSX1_148 ( .CLK(clock_i_bF_buf95), .D(_147_), .Q(_3660__15_) );
DFFPOSX1 DFFPOSX1_149 ( .CLK(clock_i_bF_buf81), .D(_148_), .Q(_3660__14_) );
DFFPOSX1 DFFPOSX1_150 ( .CLK(clock_i_bF_buf0), .D(_149_), .Q(_3660__13_) );
DFFPOSX1 DFFPOSX1_151 ( .CLK(clock_i_bF_buf76), .D(_150_), .Q(_3660__12_) );
DFFPOSX1 DFFPOSX1_152 ( .CLK(clock_i_bF_buf87), .D(_151_), .Q(_3660__11_) );
DFFPOSX1 DFFPOSX1_153 ( .CLK(clock_i_bF_buf7), .D(_152_), .Q(_3660__10_) );
DFFPOSX1 DFFPOSX1_154 ( .CLK(clock_i_bF_buf4), .D(_153_), .Q(_3660__9_) );
DFFPOSX1 DFFPOSX1_155 ( .CLK(clock_i_bF_buf15), .D(_154_), .Q(_3660__8_) );
DFFPOSX1 DFFPOSX1_156 ( .CLK(clock_i_bF_buf9), .D(_155_), .Q(_3660__7_) );
DFFPOSX1 DFFPOSX1_157 ( .CLK(clock_i_bF_buf59), .D(_156_), .Q(_3660__6_) );
DFFPOSX1 DFFPOSX1_158 ( .CLK(clock_i_bF_buf69), .D(_157_), .Q(_3660__5_) );
DFFPOSX1 DFFPOSX1_159 ( .CLK(clock_i_bF_buf51), .D(_158_), .Q(_3660__4_) );
DFFPOSX1 DFFPOSX1_160 ( .CLK(clock_i_bF_buf50), .D(_159_), .Q(_3660__3_) );
DFFPOSX1 DFFPOSX1_161 ( .CLK(clock_i_bF_buf42), .D(_160_), .Q(_3660__2_) );
DFFPOSX1 DFFPOSX1_162 ( .CLK(clock_i_bF_buf98), .D(_161_), .Q(_3660__1_) );
DFFPOSX1 DFFPOSX1_163 ( .CLK(clock_i_bF_buf64), .D(_162_), .Q(_3660__0_) );
DFFPOSX1 DFFPOSX1_164 ( .CLK(clock_i_bF_buf43), .D(_163_), .Q(_3661__63_) );
DFFPOSX1 DFFPOSX1_165 ( .CLK(clock_i_bF_buf40), .D(_164_), .Q(_3661__62_) );
DFFPOSX1 DFFPOSX1_166 ( .CLK(clock_i_bF_buf10), .D(_165_), .Q(_3661__61_) );
DFFPOSX1 DFFPOSX1_167 ( .CLK(clock_i_bF_buf61), .D(_166_), .Q(_3661__60_) );
DFFPOSX1 DFFPOSX1_168 ( .CLK(clock_i_bF_buf1), .D(_167_), .Q(_3661__59_) );
DFFPOSX1 DFFPOSX1_169 ( .CLK(clock_i_bF_buf65), .D(_168_), .Q(_3661__58_) );
DFFPOSX1 DFFPOSX1_170 ( .CLK(clock_i_bF_buf76), .D(_169_), .Q(_3661__57_) );
DFFPOSX1 DFFPOSX1_171 ( .CLK(clock_i_bF_buf76), .D(_170_), .Q(_3661__56_) );
DFFPOSX1 DFFPOSX1_172 ( .CLK(clock_i_bF_buf92), .D(_171_), .Q(_3661__55_) );
DFFPOSX1 DFFPOSX1_173 ( .CLK(clock_i_bF_buf101), .D(_172_), .Q(_3661__54_) );
DFFPOSX1 DFFPOSX1_174 ( .CLK(clock_i_bF_buf51), .D(_173_), .Q(_3661__53_) );
DFFPOSX1 DFFPOSX1_175 ( .CLK(clock_i_bF_buf88), .D(_174_), .Q(_3661__52_) );
DFFPOSX1 DFFPOSX1_176 ( .CLK(clock_i_bF_buf3), .D(_175_), .Q(_3661__51_) );
DFFPOSX1 DFFPOSX1_177 ( .CLK(clock_i_bF_buf92), .D(_176_), .Q(_3661__50_) );
DFFPOSX1 DFFPOSX1_178 ( .CLK(clock_i_bF_buf45), .D(_177_), .Q(_3661__49_) );
DFFPOSX1 DFFPOSX1_179 ( .CLK(clock_i_bF_buf90), .D(_178_), .Q(_3661__48_) );
DFFPOSX1 DFFPOSX1_180 ( .CLK(clock_i_bF_buf59), .D(_179_), .Q(_3661__47_) );
DFFPOSX1 DFFPOSX1_181 ( .CLK(clock_i_bF_buf28), .D(_180_), .Q(_3661__46_) );
DFFPOSX1 DFFPOSX1_182 ( .CLK(clock_i_bF_buf72), .D(_181_), .Q(_3661__45_) );
DFFPOSX1 DFFPOSX1_183 ( .CLK(clock_i_bF_buf4), .D(_182_), .Q(_3661__44_) );
DFFPOSX1 DFFPOSX1_184 ( .CLK(clock_i_bF_buf84), .D(_183_), .Q(_3661__43_) );
DFFPOSX1 DFFPOSX1_185 ( .CLK(clock_i_bF_buf38), .D(_184_), .Q(_3661__42_) );
DFFPOSX1 DFFPOSX1_186 ( .CLK(clock_i_bF_buf60), .D(_185_), .Q(_3661__41_) );
DFFPOSX1 DFFPOSX1_187 ( .CLK(clock_i_bF_buf60), .D(_186_), .Q(_3661__40_) );
DFFPOSX1 DFFPOSX1_188 ( .CLK(clock_i_bF_buf9), .D(_187_), .Q(_3661__39_) );
DFFPOSX1 DFFPOSX1_189 ( .CLK(clock_i_bF_buf99), .D(_188_), .Q(_3661__38_) );
DFFPOSX1 DFFPOSX1_190 ( .CLK(clock_i_bF_buf99), .D(_189_), .Q(_3661__37_) );
DFFPOSX1 DFFPOSX1_191 ( .CLK(clock_i_bF_buf85), .D(_190_), .Q(_3661__36_) );
DFFPOSX1 DFFPOSX1_192 ( .CLK(clock_i_bF_buf20), .D(_191_), .Q(_3661__35_) );
DFFPOSX1 DFFPOSX1_193 ( .CLK(clock_i_bF_buf26), .D(_192_), .Q(_3661__34_) );
DFFPOSX1 DFFPOSX1_194 ( .CLK(clock_i_bF_buf0), .D(_193_), .Q(_3661__33_) );
DFFPOSX1 DFFPOSX1_195 ( .CLK(clock_i_bF_buf24), .D(_194_), .Q(_3661__32_) );
DFFPOSX1 DFFPOSX1_196 ( .CLK(clock_i_bF_buf96), .D(_195_), .Q(_3661__31_) );
DFFPOSX1 DFFPOSX1_197 ( .CLK(clock_i_bF_buf4), .D(_196_), .Q(_3661__30_) );
DFFPOSX1 DFFPOSX1_198 ( .CLK(clock_i_bF_buf45), .D(_197_), .Q(_3661__29_) );
DFFPOSX1 DFFPOSX1_199 ( .CLK(clock_i_bF_buf29), .D(_198_), .Q(_3661__28_) );
DFFPOSX1 DFFPOSX1_200 ( .CLK(clock_i_bF_buf86), .D(_199_), .Q(_3661__27_) );
DFFPOSX1 DFFPOSX1_201 ( .CLK(clock_i_bF_buf4), .D(_200_), .Q(_3661__26_) );
DFFPOSX1 DFFPOSX1_202 ( .CLK(clock_i_bF_buf3), .D(_201_), .Q(_3661__25_) );
DFFPOSX1 DFFPOSX1_203 ( .CLK(clock_i_bF_buf62), .D(_202_), .Q(_3661__24_) );
DFFPOSX1 DFFPOSX1_204 ( .CLK(clock_i_bF_buf100), .D(_203_), .Q(_3661__23_) );
DFFPOSX1 DFFPOSX1_205 ( .CLK(clock_i_bF_buf64), .D(_204_), .Q(_3661__22_) );
DFFPOSX1 DFFPOSX1_206 ( .CLK(clock_i_bF_buf51), .D(_205_), .Q(_3661__21_) );
DFFPOSX1 DFFPOSX1_207 ( .CLK(clock_i_bF_buf60), .D(_206_), .Q(_3661__20_) );
DFFPOSX1 DFFPOSX1_208 ( .CLK(clock_i_bF_buf99), .D(_207_), .Q(_3661__19_) );
DFFPOSX1 DFFPOSX1_209 ( .CLK(clock_i_bF_buf28), .D(_208_), .Q(_3661__18_) );
DFFPOSX1 DFFPOSX1_210 ( .CLK(clock_i_bF_buf98), .D(_209_), .Q(_3661__17_) );
DFFPOSX1 DFFPOSX1_211 ( .CLK(clock_i_bF_buf9), .D(_210_), .Q(_3661__16_) );
DFFPOSX1 DFFPOSX1_212 ( .CLK(clock_i_bF_buf88), .D(_211_), .Q(_3661__15_) );
DFFPOSX1 DFFPOSX1_213 ( .CLK(clock_i_bF_buf35), .D(_212_), .Q(_3661__14_) );
DFFPOSX1 DFFPOSX1_214 ( .CLK(clock_i_bF_buf45), .D(_213_), .Q(_3661__13_) );
DFFPOSX1 DFFPOSX1_215 ( .CLK(clock_i_bF_buf76), .D(_214_), .Q(_3661__12_) );
DFFPOSX1 DFFPOSX1_216 ( .CLK(clock_i_bF_buf100), .D(_215_), .Q(_3661__11_) );
DFFPOSX1 DFFPOSX1_217 ( .CLK(clock_i_bF_buf88), .D(_216_), .Q(_3661__10_) );
DFFPOSX1 DFFPOSX1_218 ( .CLK(clock_i_bF_buf4), .D(_217_), .Q(_3661__9_) );
DFFPOSX1 DFFPOSX1_219 ( .CLK(clock_i_bF_buf15), .D(_218_), .Q(_3661__8_) );
DFFPOSX1 DFFPOSX1_220 ( .CLK(clock_i_bF_buf9), .D(_219_), .Q(_3661__7_) );
DFFPOSX1 DFFPOSX1_221 ( .CLK(clock_i_bF_buf55), .D(_220_), .Q(_3661__6_) );
DFFPOSX1 DFFPOSX1_222 ( .CLK(clock_i_bF_buf87), .D(_221_), .Q(_3661__5_) );
DFFPOSX1 DFFPOSX1_223 ( .CLK(clock_i_bF_buf51), .D(_222_), .Q(_3661__4_) );
DFFPOSX1 DFFPOSX1_224 ( .CLK(clock_i_bF_buf50), .D(_223_), .Q(_3661__3_) );
DFFPOSX1 DFFPOSX1_225 ( .CLK(clock_i_bF_buf24), .D(_224_), .Q(_3661__2_) );
DFFPOSX1 DFFPOSX1_226 ( .CLK(clock_i_bF_buf61), .D(_225_), .Q(_3661__1_) );
DFFPOSX1 DFFPOSX1_227 ( .CLK(clock_i_bF_buf44), .D(_226_), .Q(_3661__0_) );
DFFPOSX1 DFFPOSX1_228 ( .CLK(clock_i_bF_buf0), .D(_227_), .Q(_3662__63_) );
DFFPOSX1 DFFPOSX1_229 ( .CLK(clock_i_bF_buf75), .D(_228_), .Q(_3662__62_) );
DFFPOSX1 DFFPOSX1_230 ( .CLK(clock_i_bF_buf10), .D(_229_), .Q(_3662__61_) );
DFFPOSX1 DFFPOSX1_231 ( .CLK(clock_i_bF_buf57), .D(_230_), .Q(_3662__60_) );
DFFPOSX1 DFFPOSX1_232 ( .CLK(clock_i_bF_buf28), .D(_231_), .Q(_3662__59_) );
DFFPOSX1 DFFPOSX1_233 ( .CLK(clock_i_bF_buf65), .D(_232_), .Q(_3662__58_) );
DFFPOSX1 DFFPOSX1_234 ( .CLK(clock_i_bF_buf16), .D(_233_), .Q(_3662__57_) );
DFFPOSX1 DFFPOSX1_235 ( .CLK(clock_i_bF_buf76), .D(_234_), .Q(_3662__56_) );
DFFPOSX1 DFFPOSX1_236 ( .CLK(clock_i_bF_buf46), .D(_235_), .Q(_3662__55_) );
DFFPOSX1 DFFPOSX1_237 ( .CLK(clock_i_bF_buf37), .D(_236_), .Q(_3662__54_) );
DFFPOSX1 DFFPOSX1_238 ( .CLK(clock_i_bF_buf67), .D(_237_), .Q(_3662__53_) );
DFFPOSX1 DFFPOSX1_239 ( .CLK(clock_i_bF_buf88), .D(_238_), .Q(_3662__52_) );
DFFPOSX1 DFFPOSX1_240 ( .CLK(clock_i_bF_buf77), .D(_239_), .Q(_3662__51_) );
DFFPOSX1 DFFPOSX1_241 ( .CLK(clock_i_bF_buf92), .D(_240_), .Q(_3662__50_) );
DFFPOSX1 DFFPOSX1_242 ( .CLK(clock_i_bF_buf77), .D(_241_), .Q(_3662__49_) );
DFFPOSX1 DFFPOSX1_243 ( .CLK(clock_i_bF_buf90), .D(_242_), .Q(_3662__48_) );
DFFPOSX1 DFFPOSX1_244 ( .CLK(clock_i_bF_buf55), .D(_243_), .Q(_3662__47_) );
DFFPOSX1 DFFPOSX1_245 ( .CLK(clock_i_bF_buf28), .D(_244_), .Q(_3662__46_) );
DFFPOSX1 DFFPOSX1_246 ( .CLK(clock_i_bF_buf75), .D(_245_), .Q(_3662__45_) );
DFFPOSX1 DFFPOSX1_247 ( .CLK(clock_i_bF_buf79), .D(_246_), .Q(_3662__44_) );
DFFPOSX1 DFFPOSX1_248 ( .CLK(clock_i_bF_buf32), .D(_247_), .Q(_3662__43_) );
DFFPOSX1 DFFPOSX1_249 ( .CLK(clock_i_bF_buf4), .D(_248_), .Q(_3662__42_) );
DFFPOSX1 DFFPOSX1_250 ( .CLK(clock_i_bF_buf5), .D(_249_), .Q(_3662__41_) );
DFFPOSX1 DFFPOSX1_251 ( .CLK(clock_i_bF_buf16), .D(_250_), .Q(_3662__40_) );
DFFPOSX1 DFFPOSX1_252 ( .CLK(clock_i_bF_buf59), .D(_251_), .Q(_3662__39_) );
DFFPOSX1 DFFPOSX1_253 ( .CLK(clock_i_bF_buf67), .D(_252_), .Q(_3662__38_) );
DFFPOSX1 DFFPOSX1_254 ( .CLK(clock_i_bF_buf99), .D(_253_), .Q(_3662__37_) );
DFFPOSX1 DFFPOSX1_255 ( .CLK(clock_i_bF_buf70), .D(_254_), .Q(_3662__36_) );
DFFPOSX1 DFFPOSX1_256 ( .CLK(clock_i_bF_buf31), .D(_255_), .Q(_3662__35_) );
DFFPOSX1 DFFPOSX1_257 ( .CLK(clock_i_bF_buf40), .D(_256_), .Q(_3662__34_) );
DFFPOSX1 DFFPOSX1_258 ( .CLK(clock_i_bF_buf0), .D(_257_), .Q(_3662__33_) );
DFFPOSX1 DFFPOSX1_259 ( .CLK(clock_i_bF_buf24), .D(_258_), .Q(_3662__32_) );
DFFPOSX1 DFFPOSX1_260 ( .CLK(clock_i_bF_buf46), .D(_259_), .Q(_3662__31_) );
DFFPOSX1 DFFPOSX1_261 ( .CLK(clock_i_bF_buf63), .D(_260_), .Q(_3662__30_) );
DFFPOSX1 DFFPOSX1_262 ( .CLK(clock_i_bF_buf91), .D(_261_), .Q(_3662__29_) );
DFFPOSX1 DFFPOSX1_263 ( .CLK(clock_i_bF_buf29), .D(_262_), .Q(_3662__28_) );
DFFPOSX1 DFFPOSX1_264 ( .CLK(clock_i_bF_buf67), .D(_263_), .Q(_3662__27_) );
DFFPOSX1 DFFPOSX1_265 ( .CLK(clock_i_bF_buf32), .D(_264_), .Q(_3662__26_) );
DFFPOSX1 DFFPOSX1_266 ( .CLK(clock_i_bF_buf94), .D(_265_), .Q(_3662__25_) );
DFFPOSX1 DFFPOSX1_267 ( .CLK(clock_i_bF_buf62), .D(_266_), .Q(_3662__24_) );
DFFPOSX1 DFFPOSX1_268 ( .CLK(clock_i_bF_buf100), .D(_267_), .Q(_3662__23_) );
DFFPOSX1 DFFPOSX1_269 ( .CLK(clock_i_bF_buf65), .D(_268_), .Q(_3662__22_) );
DFFPOSX1 DFFPOSX1_270 ( .CLK(clock_i_bF_buf100), .D(_269_), .Q(_3662__21_) );
DFFPOSX1 DFFPOSX1_271 ( .CLK(clock_i_bF_buf45), .D(_270_), .Q(_3662__20_) );
DFFPOSX1 DFFPOSX1_272 ( .CLK(clock_i_bF_buf99), .D(_271_), .Q(_3662__19_) );
DFFPOSX1 DFFPOSX1_273 ( .CLK(clock_i_bF_buf0), .D(_272_), .Q(_3662__18_) );
DFFPOSX1 DFFPOSX1_274 ( .CLK(clock_i_bF_buf98), .D(_273_), .Q(_3662__17_) );
DFFPOSX1 DFFPOSX1_275 ( .CLK(clock_i_bF_buf86), .D(_274_), .Q(_3662__16_) );
DFFPOSX1 DFFPOSX1_276 ( .CLK(clock_i_bF_buf88), .D(_275_), .Q(_3662__15_) );
DFFPOSX1 DFFPOSX1_277 ( .CLK(clock_i_bF_buf62), .D(_276_), .Q(_3662__14_) );
DFFPOSX1 DFFPOSX1_278 ( .CLK(clock_i_bF_buf43), .D(_277_), .Q(_3662__13_) );
DFFPOSX1 DFFPOSX1_279 ( .CLK(clock_i_bF_buf64), .D(_278_), .Q(_3662__12_) );
DFFPOSX1 DFFPOSX1_280 ( .CLK(clock_i_bF_buf87), .D(_279_), .Q(_3662__11_) );
DFFPOSX1 DFFPOSX1_281 ( .CLK(clock_i_bF_buf7), .D(_280_), .Q(_3662__10_) );
DFFPOSX1 DFFPOSX1_282 ( .CLK(clock_i_bF_buf63), .D(_281_), .Q(_3662__9_) );
DFFPOSX1 DFFPOSX1_283 ( .CLK(clock_i_bF_buf15), .D(_282_), .Q(_3662__8_) );
DFFPOSX1 DFFPOSX1_284 ( .CLK(clock_i_bF_buf59), .D(_283_), .Q(_3662__7_) );
DFFPOSX1 DFFPOSX1_285 ( .CLK(clock_i_bF_buf59), .D(_284_), .Q(_3662__6_) );
DFFPOSX1 DFFPOSX1_286 ( .CLK(clock_i_bF_buf100), .D(_285_), .Q(_3662__5_) );
DFFPOSX1 DFFPOSX1_287 ( .CLK(clock_i_bF_buf51), .D(_286_), .Q(_3662__4_) );
DFFPOSX1 DFFPOSX1_288 ( .CLK(clock_i_bF_buf100), .D(_287_), .Q(_3662__3_) );
DFFPOSX1 DFFPOSX1_289 ( .CLK(clock_i_bF_buf47), .D(_288_), .Q(_3662__2_) );
DFFPOSX1 DFFPOSX1_290 ( .CLK(clock_i_bF_buf98), .D(_289_), .Q(_3662__1_) );
DFFPOSX1 DFFPOSX1_291 ( .CLK(clock_i_bF_buf33), .D(_290_), .Q(_3662__0_) );
DFFPOSX1 DFFPOSX1_292 ( .CLK(clock_i_bF_buf79), .D(_291_), .Q(_3663__63_) );
DFFPOSX1 DFFPOSX1_293 ( .CLK(clock_i_bF_buf25), .D(_292_), .Q(_3663__62_) );
DFFPOSX1 DFFPOSX1_294 ( .CLK(clock_i_bF_buf10), .D(_293_), .Q(_3663__61_) );
DFFPOSX1 DFFPOSX1_295 ( .CLK(clock_i_bF_buf14), .D(_294_), .Q(_3663__60_) );
DFFPOSX1 DFFPOSX1_296 ( .CLK(clock_i_bF_buf43), .D(_295_), .Q(_3663__59_) );
DFFPOSX1 DFFPOSX1_297 ( .CLK(clock_i_bF_buf21), .D(_296_), .Q(_3663__58_) );
DFFPOSX1 DFFPOSX1_298 ( .CLK(clock_i_bF_buf42), .D(_297_), .Q(_3663__57_) );
DFFPOSX1 DFFPOSX1_299 ( .CLK(clock_i_bF_buf76), .D(_298_), .Q(_3663__56_) );
DFFPOSX1 DFFPOSX1_300 ( .CLK(clock_i_bF_buf98), .D(_299_), .Q(_3663__55_) );
DFFPOSX1 DFFPOSX1_301 ( .CLK(clock_i_bF_buf73), .D(_300_), .Q(_3663__54_) );
DFFPOSX1 DFFPOSX1_302 ( .CLK(clock_i_bF_buf19), .D(_301_), .Q(_3663__53_) );
DFFPOSX1 DFFPOSX1_303 ( .CLK(clock_i_bF_buf88), .D(_302_), .Q(_3663__52_) );
DFFPOSX1 DFFPOSX1_304 ( .CLK(clock_i_bF_buf77), .D(_303_), .Q(_3663__51_) );
DFFPOSX1 DFFPOSX1_305 ( .CLK(clock_i_bF_buf36), .D(_304_), .Q(_3663__50_) );
DFFPOSX1 DFFPOSX1_306 ( .CLK(clock_i_bF_buf77), .D(_305_), .Q(_3663__49_) );
DFFPOSX1 DFFPOSX1_307 ( .CLK(clock_i_bF_buf28), .D(_306_), .Q(_3663__48_) );
DFFPOSX1 DFFPOSX1_308 ( .CLK(clock_i_bF_buf52), .D(_307_), .Q(_3663__47_) );
DFFPOSX1 DFFPOSX1_309 ( .CLK(clock_i_bF_buf37), .D(_308_), .Q(_3663__46_) );
DFFPOSX1 DFFPOSX1_310 ( .CLK(clock_i_bF_buf25), .D(_309_), .Q(_3663__45_) );
DFFPOSX1 DFFPOSX1_311 ( .CLK(clock_i_bF_buf30), .D(_310_), .Q(_3663__44_) );
DFFPOSX1 DFFPOSX1_312 ( .CLK(clock_i_bF_buf97), .D(_311_), .Q(_3663__43_) );
DFFPOSX1 DFFPOSX1_313 ( .CLK(clock_i_bF_buf80), .D(_312_), .Q(_3663__42_) );
DFFPOSX1 DFFPOSX1_314 ( .CLK(clock_i_bF_buf5), .D(_313_), .Q(_3663__41_) );
DFFPOSX1 DFFPOSX1_315 ( .CLK(clock_i_bF_buf16), .D(_314_), .Q(_3663__40_) );
DFFPOSX1 DFFPOSX1_316 ( .CLK(clock_i_bF_buf59), .D(_315_), .Q(_3663__39_) );
DFFPOSX1 DFFPOSX1_317 ( .CLK(clock_i_bF_buf75), .D(_316_), .Q(_3663__38_) );
DFFPOSX1 DFFPOSX1_318 ( .CLK(clock_i_bF_buf95), .D(_317_), .Q(_3663__37_) );
DFFPOSX1 DFFPOSX1_319 ( .CLK(clock_i_bF_buf85), .D(_318_), .Q(_3663__36_) );
DFFPOSX1 DFFPOSX1_320 ( .CLK(clock_i_bF_buf31), .D(_319_), .Q(_3663__35_) );
DFFPOSX1 DFFPOSX1_321 ( .CLK(clock_i_bF_buf53), .D(_320_), .Q(_3663__34_) );
DFFPOSX1 DFFPOSX1_322 ( .CLK(clock_i_bF_buf0), .D(_321_), .Q(_3663__33_) );
DFFPOSX1 DFFPOSX1_323 ( .CLK(clock_i_bF_buf38), .D(_322_), .Q(_3663__32_) );
DFFPOSX1 DFFPOSX1_324 ( .CLK(clock_i_bF_buf46), .D(_323_), .Q(_3663__31_) );
DFFPOSX1 DFFPOSX1_325 ( .CLK(clock_i_bF_buf4), .D(_324_), .Q(_3663__30_) );
DFFPOSX1 DFFPOSX1_326 ( .CLK(clock_i_bF_buf77), .D(_325_), .Q(_3663__29_) );
DFFPOSX1 DFFPOSX1_327 ( .CLK(clock_i_bF_buf80), .D(_326_), .Q(_3663__28_) );
DFFPOSX1 DFFPOSX1_328 ( .CLK(clock_i_bF_buf95), .D(_327_), .Q(_3663__27_) );
DFFPOSX1 DFFPOSX1_329 ( .CLK(clock_i_bF_buf32), .D(_328_), .Q(_3663__26_) );
DFFPOSX1 DFFPOSX1_330 ( .CLK(clock_i_bF_buf85), .D(_329_), .Q(_3663__25_) );
DFFPOSX1 DFFPOSX1_331 ( .CLK(clock_i_bF_buf76), .D(_330_), .Q(_3663__24_) );
DFFPOSX1 DFFPOSX1_332 ( .CLK(clock_i_bF_buf19), .D(_331_), .Q(_3663__23_) );
DFFPOSX1 DFFPOSX1_333 ( .CLK(clock_i_bF_buf81), .D(_332_), .Q(_3663__22_) );
DFFPOSX1 DFFPOSX1_334 ( .CLK(clock_i_bF_buf19), .D(_333_), .Q(_3663__21_) );
DFFPOSX1 DFFPOSX1_335 ( .CLK(clock_i_bF_buf75), .D(_334_), .Q(_3663__20_) );
DFFPOSX1 DFFPOSX1_336 ( .CLK(clock_i_bF_buf95), .D(_335_), .Q(_3663__19_) );
DFFPOSX1 DFFPOSX1_337 ( .CLK(clock_i_bF_buf0), .D(_336_), .Q(_3663__18_) );
DFFPOSX1 DFFPOSX1_338 ( .CLK(clock_i_bF_buf98), .D(_337_), .Q(_3663__17_) );
DFFPOSX1 DFFPOSX1_339 ( .CLK(clock_i_bF_buf95), .D(_338_), .Q(_3663__16_) );
DFFPOSX1 DFFPOSX1_340 ( .CLK(clock_i_bF_buf99), .D(_339_), .Q(_3663__15_) );
DFFPOSX1 DFFPOSX1_341 ( .CLK(clock_i_bF_buf94), .D(_340_), .Q(_3663__14_) );
DFFPOSX1 DFFPOSX1_342 ( .CLK(clock_i_bF_buf77), .D(_341_), .Q(_3663__13_) );
DFFPOSX1 DFFPOSX1_343 ( .CLK(clock_i_bF_buf33), .D(_342_), .Q(_3663__12_) );
DFFPOSX1 DFFPOSX1_344 ( .CLK(clock_i_bF_buf87), .D(_343_), .Q(_3663__11_) );
DFFPOSX1 DFFPOSX1_345 ( .CLK(clock_i_bF_buf7), .D(_344_), .Q(_3663__10_) );
DFFPOSX1 DFFPOSX1_346 ( .CLK(clock_i_bF_buf4), .D(_345_), .Q(_3663__9_) );
DFFPOSX1 DFFPOSX1_347 ( .CLK(clock_i_bF_buf98), .D(_346_), .Q(_3663__8_) );
DFFPOSX1 DFFPOSX1_348 ( .CLK(clock_i_bF_buf59), .D(_347_), .Q(_3663__7_) );
DFFPOSX1 DFFPOSX1_349 ( .CLK(clock_i_bF_buf55), .D(_348_), .Q(_3663__6_) );
DFFPOSX1 DFFPOSX1_350 ( .CLK(clock_i_bF_buf10), .D(_349_), .Q(_3663__5_) );
DFFPOSX1 DFFPOSX1_351 ( .CLK(clock_i_bF_buf25), .D(_350_), .Q(_3663__4_) );
DFFPOSX1 DFFPOSX1_352 ( .CLK(clock_i_bF_buf19), .D(_351_), .Q(_3663__3_) );
DFFPOSX1 DFFPOSX1_353 ( .CLK(clock_i_bF_buf80), .D(_352_), .Q(_3663__2_) );
DFFPOSX1 DFFPOSX1_354 ( .CLK(clock_i_bF_buf98), .D(_353_), .Q(_3663__1_) );
DFFPOSX1 DFFPOSX1_355 ( .CLK(clock_i_bF_buf44), .D(_354_), .Q(_3663__0_) );
DFFPOSX1 DFFPOSX1_356 ( .CLK(clock_i_bF_buf57), .D(_355_), .Q(_3652__63_) );
DFFPOSX1 DFFPOSX1_357 ( .CLK(clock_i_bF_buf57), .D(_356_), .Q(_3652__62_) );
DFFPOSX1 DFFPOSX1_358 ( .CLK(clock_i_bF_buf22), .D(_357_), .Q(_3652__61_) );
DFFPOSX1 DFFPOSX1_359 ( .CLK(clock_i_bF_buf98), .D(_358_), .Q(_3652__60_) );
DFFPOSX1 DFFPOSX1_360 ( .CLK(clock_i_bF_buf61), .D(_359_), .Q(_3652__59_) );
DFFPOSX1 DFFPOSX1_361 ( .CLK(clock_i_bF_buf36), .D(_360_), .Q(_3652__58_) );
DFFPOSX1 DFFPOSX1_362 ( .CLK(clock_i_bF_buf36), .D(_361_), .Q(_3652__57_) );
DFFPOSX1 DFFPOSX1_363 ( .CLK(clock_i_bF_buf36), .D(_362_), .Q(_3652__56_) );
DFFPOSX1 DFFPOSX1_364 ( .CLK(clock_i_bF_buf96), .D(_363_), .Q(_3652__55_) );
DFFPOSX1 DFFPOSX1_365 ( .CLK(clock_i_bF_buf96), .D(_364_), .Q(_3652__54_) );
DFFPOSX1 DFFPOSX1_366 ( .CLK(clock_i_bF_buf27), .D(_365_), .Q(_3652__53_) );
DFFPOSX1 DFFPOSX1_367 ( .CLK(clock_i_bF_buf96), .D(_366_), .Q(_3652__52_) );
DFFPOSX1 DFFPOSX1_368 ( .CLK(clock_i_bF_buf8), .D(_367_), .Q(_3652__51_) );
DFFPOSX1 DFFPOSX1_369 ( .CLK(clock_i_bF_buf56), .D(_368_), .Q(_3652__50_) );
DFFPOSX1 DFFPOSX1_370 ( .CLK(clock_i_bF_buf96), .D(_369_), .Q(_3652__49_) );
DFFPOSX1 DFFPOSX1_371 ( .CLK(clock_i_bF_buf89), .D(_370_), .Q(_3652__48_) );
DFFPOSX1 DFFPOSX1_372 ( .CLK(clock_i_bF_buf27), .D(_371_), .Q(_3652__47_) );
DFFPOSX1 DFFPOSX1_373 ( .CLK(clock_i_bF_buf54), .D(_372_), .Q(_3652__46_) );
DFFPOSX1 DFFPOSX1_374 ( .CLK(clock_i_bF_buf83), .D(_373_), .Q(_3652__45_) );
DFFPOSX1 DFFPOSX1_375 ( .CLK(clock_i_bF_buf101), .D(_374_), .Q(_3652__44_) );
DFFPOSX1 DFFPOSX1_376 ( .CLK(clock_i_bF_buf69), .D(_375_), .Q(_3652__43_) );
DFFPOSX1 DFFPOSX1_377 ( .CLK(clock_i_bF_buf84), .D(_376_), .Q(_3652__42_) );
DFFPOSX1 DFFPOSX1_378 ( .CLK(clock_i_bF_buf84), .D(_377_), .Q(_3652__41_) );
DFFPOSX1 DFFPOSX1_379 ( .CLK(clock_i_bF_buf84), .D(_378_), .Q(_3652__40_) );
DFFPOSX1 DFFPOSX1_380 ( .CLK(clock_i_bF_buf87), .D(_379_), .Q(_3652__39_) );
DFFPOSX1 DFFPOSX1_381 ( .CLK(clock_i_bF_buf52), .D(_380_), .Q(_3652__38_) );
DFFPOSX1 DFFPOSX1_382 ( .CLK(clock_i_bF_buf52), .D(_381_), .Q(_3652__37_) );
DFFPOSX1 DFFPOSX1_383 ( .CLK(clock_i_bF_buf69), .D(_382_), .Q(_3652__36_) );
DFFPOSX1 DFFPOSX1_384 ( .CLK(clock_i_bF_buf87), .D(_383_), .Q(_3652__35_) );
DFFPOSX1 DFFPOSX1_385 ( .CLK(clock_i_bF_buf39), .D(_384_), .Q(_3652__34_) );
DFFPOSX1 DFFPOSX1_386 ( .CLK(clock_i_bF_buf39), .D(_385_), .Q(_3652__33_) );
DFFPOSX1 DFFPOSX1_387 ( .CLK(clock_i_bF_buf87), .D(_386_), .Q(_3652__32_) );
DFFPOSX1 DFFPOSX1_388 ( .CLK(clock_i_bF_buf23), .D(_387_), .Q(_3652__31_) );
DFFPOSX1 DFFPOSX1_389 ( .CLK(clock_i_bF_buf58), .D(_388_), .Q(_3652__30_) );
DFFPOSX1 DFFPOSX1_390 ( .CLK(clock_i_bF_buf58), .D(_389_), .Q(_3652__29_) );
DFFPOSX1 DFFPOSX1_391 ( .CLK(clock_i_bF_buf10), .D(_390_), .Q(_3652__28_) );
DFFPOSX1 DFFPOSX1_392 ( .CLK(clock_i_bF_buf83), .D(_391_), .Q(_3652__27_) );
DFFPOSX1 DFFPOSX1_393 ( .CLK(clock_i_bF_buf78), .D(_392_), .Q(_3652__26_) );
DFFPOSX1 DFFPOSX1_394 ( .CLK(clock_i_bF_buf83), .D(_393_), .Q(_3652__25_) );
DFFPOSX1 DFFPOSX1_395 ( .CLK(clock_i_bF_buf97), .D(_394_), .Q(_3652__24_) );
DFFPOSX1 DFFPOSX1_396 ( .CLK(clock_i_bF_buf22), .D(_395_), .Q(_3652__23_) );
DFFPOSX1 DFFPOSX1_397 ( .CLK(clock_i_bF_buf18), .D(_396_), .Q(_3652__22_) );
DFFPOSX1 DFFPOSX1_398 ( .CLK(clock_i_bF_buf18), .D(_397_), .Q(_3652__21_) );
DFFPOSX1 DFFPOSX1_399 ( .CLK(clock_i_bF_buf2), .D(_398_), .Q(_3652__20_) );
DFFPOSX1 DFFPOSX1_400 ( .CLK(clock_i_bF_buf12), .D(_399_), .Q(_3652__19_) );
DFFPOSX1 DFFPOSX1_401 ( .CLK(clock_i_bF_buf12), .D(_400_), .Q(_3652__18_) );
DFFPOSX1 DFFPOSX1_402 ( .CLK(clock_i_bF_buf22), .D(_401_), .Q(_3652__17_) );
DFFPOSX1 DFFPOSX1_403 ( .CLK(clock_i_bF_buf80), .D(_402_), .Q(_3652__16_) );
DFFPOSX1 DFFPOSX1_404 ( .CLK(clock_i_bF_buf23), .D(_403_), .Q(_3652__15_) );
DFFPOSX1 DFFPOSX1_405 ( .CLK(clock_i_bF_buf2), .D(_404_), .Q(_3652__14_) );
DFFPOSX1 DFFPOSX1_406 ( .CLK(clock_i_bF_buf11), .D(_405_), .Q(_3652__13_) );
DFFPOSX1 DFFPOSX1_407 ( .CLK(clock_i_bF_buf11), .D(_406_), .Q(_3652__12_) );
DFFPOSX1 DFFPOSX1_408 ( .CLK(clock_i_bF_buf22), .D(_407_), .Q(_3652__11_) );
DFFPOSX1 DFFPOSX1_409 ( .CLK(clock_i_bF_buf18), .D(_408_), .Q(_3652__10_) );
DFFPOSX1 DFFPOSX1_410 ( .CLK(clock_i_bF_buf23), .D(_409_), .Q(_3652__9_) );
DFFPOSX1 DFFPOSX1_411 ( .CLK(clock_i_bF_buf96), .D(_410_), .Q(_3652__8_) );
DFFPOSX1 DFFPOSX1_412 ( .CLK(clock_i_bF_buf101), .D(_411_), .Q(_3652__7_) );
DFFPOSX1 DFFPOSX1_413 ( .CLK(clock_i_bF_buf73), .D(_412_), .Q(_3652__6_) );
DFFPOSX1 DFFPOSX1_414 ( .CLK(clock_i_bF_buf91), .D(_413_), .Q(_3652__5_) );
DFFPOSX1 DFFPOSX1_415 ( .CLK(clock_i_bF_buf91), .D(_414_), .Q(_3652__4_) );
DFFPOSX1 DFFPOSX1_416 ( .CLK(clock_i_bF_buf83), .D(_415_), .Q(_3652__3_) );
DFFPOSX1 DFFPOSX1_417 ( .CLK(clock_i_bF_buf78), .D(_416_), .Q(_3652__2_) );
DFFPOSX1 DFFPOSX1_418 ( .CLK(clock_i_bF_buf32), .D(_417_), .Q(_3652__1_) );
DFFPOSX1 DFFPOSX1_419 ( .CLK(clock_i_bF_buf58), .D(_418_), .Q(_3652__0_) );
DFFPOSX1 DFFPOSX1_420 ( .CLK(clock_i_bF_buf92), .D(_419_), .Q(_3653__63_) );
DFFPOSX1 DFFPOSX1_421 ( .CLK(clock_i_bF_buf8), .D(_420_), .Q(_3653__62_) );
DFFPOSX1 DFFPOSX1_422 ( .CLK(clock_i_bF_buf57), .D(_421_), .Q(_3653__61_) );
DFFPOSX1 DFFPOSX1_423 ( .CLK(clock_i_bF_buf8), .D(_422_), .Q(_3653__60_) );
DFFPOSX1 DFFPOSX1_424 ( .CLK(clock_i_bF_buf27), .D(_423_), .Q(_3653__59_) );
DFFPOSX1 DFFPOSX1_425 ( .CLK(clock_i_bF_buf36), .D(_424_), .Q(_3653__58_) );
DFFPOSX1 DFFPOSX1_426 ( .CLK(clock_i_bF_buf92), .D(_425_), .Q(_3653__57_) );
DFFPOSX1 DFFPOSX1_427 ( .CLK(clock_i_bF_buf27), .D(_426_), .Q(_3653__56_) );
DFFPOSX1 DFFPOSX1_428 ( .CLK(clock_i_bF_buf89), .D(_427_), .Q(_3653__55_) );
DFFPOSX1 DFFPOSX1_429 ( .CLK(clock_i_bF_buf89), .D(_428_), .Q(_3653__54_) );
DFFPOSX1 DFFPOSX1_430 ( .CLK(clock_i_bF_buf89), .D(_429_), .Q(_3653__53_) );
DFFPOSX1 DFFPOSX1_431 ( .CLK(clock_i_bF_buf27), .D(_430_), .Q(_3653__52_) );
DFFPOSX1 DFFPOSX1_432 ( .CLK(clock_i_bF_buf89), .D(_431_), .Q(_3653__51_) );
DFFPOSX1 DFFPOSX1_433 ( .CLK(clock_i_bF_buf89), .D(_432_), .Q(_3653__50_) );
DFFPOSX1 DFFPOSX1_434 ( .CLK(clock_i_bF_buf89), .D(_433_), .Q(_3653__49_) );
DFFPOSX1 DFFPOSX1_435 ( .CLK(clock_i_bF_buf89), .D(_434_), .Q(_3653__48_) );
DFFPOSX1 DFFPOSX1_436 ( .CLK(clock_i_bF_buf84), .D(_435_), .Q(_3653__47_) );
DFFPOSX1 DFFPOSX1_437 ( .CLK(clock_i_bF_buf78), .D(_436_), .Q(_3653__46_) );
DFFPOSX1 DFFPOSX1_438 ( .CLK(clock_i_bF_buf78), .D(_437_), .Q(_3653__45_) );
DFFPOSX1 DFFPOSX1_439 ( .CLK(clock_i_bF_buf101), .D(_438_), .Q(_3653__44_) );
DFFPOSX1 DFFPOSX1_440 ( .CLK(clock_i_bF_buf84), .D(_439_), .Q(_3653__43_) );
DFFPOSX1 DFFPOSX1_441 ( .CLK(clock_i_bF_buf84), .D(_440_), .Q(_3653__42_) );
DFFPOSX1 DFFPOSX1_442 ( .CLK(clock_i_bF_buf84), .D(_441_), .Q(_3653__41_) );
DFFPOSX1 DFFPOSX1_443 ( .CLK(clock_i_bF_buf84), .D(_442_), .Q(_3653__40_) );
DFFPOSX1 DFFPOSX1_444 ( .CLK(clock_i_bF_buf87), .D(_443_), .Q(_3653__39_) );
DFFPOSX1 DFFPOSX1_445 ( .CLK(clock_i_bF_buf52), .D(_444_), .Q(_3653__38_) );
DFFPOSX1 DFFPOSX1_446 ( .CLK(clock_i_bF_buf69), .D(_445_), .Q(_3653__37_) );
DFFPOSX1 DFFPOSX1_447 ( .CLK(clock_i_bF_buf69), .D(_446_), .Q(_3653__36_) );
DFFPOSX1 DFFPOSX1_448 ( .CLK(clock_i_bF_buf69), .D(_447_), .Q(_3653__35_) );
DFFPOSX1 DFFPOSX1_449 ( .CLK(clock_i_bF_buf69), .D(_448_), .Q(_3653__34_) );
DFFPOSX1 DFFPOSX1_450 ( .CLK(clock_i_bF_buf52), .D(_449_), .Q(_3653__33_) );
DFFPOSX1 DFFPOSX1_451 ( .CLK(clock_i_bF_buf39), .D(_450_), .Q(_3653__32_) );
DFFPOSX1 DFFPOSX1_452 ( .CLK(clock_i_bF_buf10), .D(_451_), .Q(_3653__31_) );
DFFPOSX1 DFFPOSX1_453 ( .CLK(clock_i_bF_buf58), .D(_452_), .Q(_3653__30_) );
DFFPOSX1 DFFPOSX1_454 ( .CLK(clock_i_bF_buf58), .D(_453_), .Q(_3653__29_) );
DFFPOSX1 DFFPOSX1_455 ( .CLK(clock_i_bF_buf58), .D(_454_), .Q(_3653__28_) );
DFFPOSX1 DFFPOSX1_456 ( .CLK(clock_i_bF_buf101), .D(_455_), .Q(_3653__27_) );
DFFPOSX1 DFFPOSX1_457 ( .CLK(clock_i_bF_buf93), .D(_456_), .Q(_3653__26_) );
DFFPOSX1 DFFPOSX1_458 ( .CLK(clock_i_bF_buf73), .D(_457_), .Q(_3653__25_) );
DFFPOSX1 DFFPOSX1_459 ( .CLK(clock_i_bF_buf97), .D(_458_), .Q(_3653__24_) );
DFFPOSX1 DFFPOSX1_460 ( .CLK(clock_i_bF_buf18), .D(_459_), .Q(_3653__23_) );
DFFPOSX1 DFFPOSX1_461 ( .CLK(clock_i_bF_buf18), .D(_460_), .Q(_3653__22_) );
DFFPOSX1 DFFPOSX1_462 ( .CLK(clock_i_bF_buf12), .D(_461_), .Q(_3653__21_) );
DFFPOSX1 DFFPOSX1_463 ( .CLK(clock_i_bF_buf80), .D(_462_), .Q(_3653__20_) );
DFFPOSX1 DFFPOSX1_464 ( .CLK(clock_i_bF_buf54), .D(_463_), .Q(_3653__19_) );
DFFPOSX1 DFFPOSX1_465 ( .CLK(clock_i_bF_buf27), .D(_464_), .Q(_3653__18_) );
DFFPOSX1 DFFPOSX1_466 ( .CLK(clock_i_bF_buf54), .D(_465_), .Q(_3653__17_) );
DFFPOSX1 DFFPOSX1_467 ( .CLK(clock_i_bF_buf54), .D(_466_), .Q(_3653__16_) );
DFFPOSX1 DFFPOSX1_468 ( .CLK(clock_i_bF_buf30), .D(_467_), .Q(_3653__15_) );
DFFPOSX1 DFFPOSX1_469 ( .CLK(clock_i_bF_buf80), .D(_468_), .Q(_3653__14_) );
DFFPOSX1 DFFPOSX1_470 ( .CLK(clock_i_bF_buf2), .D(_469_), .Q(_3653__13_) );
DFFPOSX1 DFFPOSX1_471 ( .CLK(clock_i_bF_buf11), .D(_470_), .Q(_3653__12_) );
DFFPOSX1 DFFPOSX1_472 ( .CLK(clock_i_bF_buf54), .D(_471_), .Q(_3653__11_) );
DFFPOSX1 DFFPOSX1_473 ( .CLK(clock_i_bF_buf96), .D(_472_), .Q(_3653__10_) );
DFFPOSX1 DFFPOSX1_474 ( .CLK(clock_i_bF_buf54), .D(_473_), .Q(_3653__9_) );
DFFPOSX1 DFFPOSX1_475 ( .CLK(clock_i_bF_buf54), .D(_474_), .Q(_3653__8_) );
DFFPOSX1 DFFPOSX1_476 ( .CLK(clock_i_bF_buf93), .D(_475_), .Q(_3653__7_) );
DFFPOSX1 DFFPOSX1_477 ( .CLK(clock_i_bF_buf93), .D(_476_), .Q(_3653__6_) );
DFFPOSX1 DFFPOSX1_478 ( .CLK(clock_i_bF_buf97), .D(_477_), .Q(_3653__5_) );
DFFPOSX1 DFFPOSX1_479 ( .CLK(clock_i_bF_buf73), .D(_478_), .Q(_3653__4_) );
DFFPOSX1 DFFPOSX1_480 ( .CLK(clock_i_bF_buf93), .D(_479_), .Q(_3653__3_) );
DFFPOSX1 DFFPOSX1_481 ( .CLK(clock_i_bF_buf83), .D(_480_), .Q(_3653__2_) );
DFFPOSX1 DFFPOSX1_482 ( .CLK(clock_i_bF_buf83), .D(_481_), .Q(_3653__1_) );
DFFPOSX1 DFFPOSX1_483 ( .CLK(clock_i_bF_buf37), .D(_482_), .Q(_3653__0_) );
DFFPOSX1 DFFPOSX1_484 ( .CLK(clock_i_bF_buf57), .D(_483_), .Q(_3654__63_) );
DFFPOSX1 DFFPOSX1_485 ( .CLK(clock_i_bF_buf8), .D(_484_), .Q(_3654__62_) );
DFFPOSX1 DFFPOSX1_486 ( .CLK(clock_i_bF_buf57), .D(_485_), .Q(_3654__61_) );
DFFPOSX1 DFFPOSX1_487 ( .CLK(clock_i_bF_buf8), .D(_486_), .Q(_3654__60_) );
DFFPOSX1 DFFPOSX1_488 ( .CLK(clock_i_bF_buf36), .D(_487_), .Q(_3654__59_) );
DFFPOSX1 DFFPOSX1_489 ( .CLK(clock_i_bF_buf8), .D(_488_), .Q(_3654__58_) );
DFFPOSX1 DFFPOSX1_490 ( .CLK(clock_i_bF_buf56), .D(_489_), .Q(_3654__57_) );
DFFPOSX1 DFFPOSX1_491 ( .CLK(clock_i_bF_buf8), .D(_490_), .Q(_3654__56_) );
DFFPOSX1 DFFPOSX1_492 ( .CLK(clock_i_bF_buf56), .D(_491_), .Q(_3654__55_) );
DFFPOSX1 DFFPOSX1_493 ( .CLK(clock_i_bF_buf2), .D(_492_), .Q(_3654__54_) );
DFFPOSX1 DFFPOSX1_494 ( .CLK(clock_i_bF_buf27), .D(_493_), .Q(_3654__53_) );
DFFPOSX1 DFFPOSX1_495 ( .CLK(clock_i_bF_buf12), .D(_494_), .Q(_3654__52_) );
DFFPOSX1 DFFPOSX1_496 ( .CLK(clock_i_bF_buf56), .D(_495_), .Q(_3654__51_) );
DFFPOSX1 DFFPOSX1_497 ( .CLK(clock_i_bF_buf56), .D(_496_), .Q(_3654__50_) );
DFFPOSX1 DFFPOSX1_498 ( .CLK(clock_i_bF_buf22), .D(_497_), .Q(_3654__49_) );
DFFPOSX1 DFFPOSX1_499 ( .CLK(clock_i_bF_buf12), .D(_498_), .Q(_3654__48_) );
DFFPOSX1 DFFPOSX1_500 ( .CLK(clock_i_bF_buf56), .D(_499_), .Q(_3654__47_) );
DFFPOSX1 DFFPOSX1_501 ( .CLK(clock_i_bF_buf22), .D(_500_), .Q(_3654__46_) );
DFFPOSX1 DFFPOSX1_502 ( .CLK(clock_i_bF_buf39), .D(_501_), .Q(_3654__45_) );
DFFPOSX1 DFFPOSX1_503 ( .CLK(clock_i_bF_buf14), .D(_502_), .Q(_3654__44_) );
DFFPOSX1 DFFPOSX1_504 ( .CLK(clock_i_bF_buf14), .D(_503_), .Q(_3654__43_) );
DFFPOSX1 DFFPOSX1_505 ( .CLK(clock_i_bF_buf84), .D(_504_), .Q(_3654__42_) );
DFFPOSX1 DFFPOSX1_506 ( .CLK(clock_i_bF_buf58), .D(_505_), .Q(_3654__41_) );
DFFPOSX1 DFFPOSX1_507 ( .CLK(clock_i_bF_buf69), .D(_506_), .Q(_3654__40_) );
DFFPOSX1 DFFPOSX1_508 ( .CLK(clock_i_bF_buf69), .D(_507_), .Q(_3654__39_) );
DFFPOSX1 DFFPOSX1_509 ( .CLK(clock_i_bF_buf42), .D(_508_), .Q(_3654__38_) );
DFFPOSX1 DFFPOSX1_510 ( .CLK(clock_i_bF_buf52), .D(_509_), .Q(_3654__37_) );
DFFPOSX1 DFFPOSX1_511 ( .CLK(clock_i_bF_buf39), .D(_510_), .Q(_3654__36_) );
DFFPOSX1 DFFPOSX1_512 ( .CLK(clock_i_bF_buf14), .D(_511_), .Q(_3654__35_) );
DFFPOSX1 DFFPOSX1_513 ( .CLK(clock_i_bF_buf39), .D(_512_), .Q(_3654__34_) );
DFFPOSX1 DFFPOSX1_514 ( .CLK(clock_i_bF_buf39), .D(_513_), .Q(_3654__33_) );
DFFPOSX1 DFFPOSX1_515 ( .CLK(clock_i_bF_buf55), .D(_514_), .Q(_3654__32_) );
DFFPOSX1 DFFPOSX1_516 ( .CLK(clock_i_bF_buf14), .D(_515_), .Q(_3654__31_) );
DFFPOSX1 DFFPOSX1_517 ( .CLK(clock_i_bF_buf54), .D(_516_), .Q(_3654__30_) );
DFFPOSX1 DFFPOSX1_518 ( .CLK(clock_i_bF_buf54), .D(_517_), .Q(_3654__29_) );
DFFPOSX1 DFFPOSX1_519 ( .CLK(clock_i_bF_buf12), .D(_518_), .Q(_3654__28_) );
DFFPOSX1 DFFPOSX1_520 ( .CLK(clock_i_bF_buf93), .D(_519_), .Q(_3654__27_) );
DFFPOSX1 DFFPOSX1_521 ( .CLK(clock_i_bF_buf23), .D(_520_), .Q(_3654__26_) );
DFFPOSX1 DFFPOSX1_522 ( .CLK(clock_i_bF_buf69), .D(_521_), .Q(_3654__25_) );
DFFPOSX1 DFFPOSX1_523 ( .CLK(clock_i_bF_buf58), .D(_522_), .Q(_3654__24_) );
DFFPOSX1 DFFPOSX1_524 ( .CLK(clock_i_bF_buf58), .D(_523_), .Q(_3654__23_) );
DFFPOSX1 DFFPOSX1_525 ( .CLK(clock_i_bF_buf11), .D(_524_), .Q(_3654__22_) );
DFFPOSX1 DFFPOSX1_526 ( .CLK(clock_i_bF_buf2), .D(_525_), .Q(_3654__21_) );
DFFPOSX1 DFFPOSX1_527 ( .CLK(clock_i_bF_buf18), .D(_526_), .Q(_3654__20_) );
DFFPOSX1 DFFPOSX1_528 ( .CLK(clock_i_bF_buf22), .D(_527_), .Q(_3654__19_) );
DFFPOSX1 DFFPOSX1_529 ( .CLK(clock_i_bF_buf23), .D(_528_), .Q(_3654__18_) );
DFFPOSX1 DFFPOSX1_530 ( .CLK(clock_i_bF_buf12), .D(_529_), .Q(_3654__17_) );
DFFPOSX1 DFFPOSX1_531 ( .CLK(clock_i_bF_buf12), .D(_530_), .Q(_3654__16_) );
DFFPOSX1 DFFPOSX1_532 ( .CLK(clock_i_bF_buf23), .D(_531_), .Q(_3654__15_) );
DFFPOSX1 DFFPOSX1_533 ( .CLK(clock_i_bF_buf15), .D(_532_), .Q(_3654__14_) );
DFFPOSX1 DFFPOSX1_534 ( .CLK(clock_i_bF_buf2), .D(_533_), .Q(_3654__13_) );
DFFPOSX1 DFFPOSX1_535 ( .CLK(clock_i_bF_buf11), .D(_534_), .Q(_3654__12_) );
DFFPOSX1 DFFPOSX1_536 ( .CLK(clock_i_bF_buf2), .D(_535_), .Q(_3654__11_) );
DFFPOSX1 DFFPOSX1_537 ( .CLK(clock_i_bF_buf11), .D(_536_), .Q(_3654__10_) );
DFFPOSX1 DFFPOSX1_538 ( .CLK(clock_i_bF_buf23), .D(_537_), .Q(_3654__9_) );
DFFPOSX1 DFFPOSX1_539 ( .CLK(clock_i_bF_buf18), .D(_538_), .Q(_3654__8_) );
DFFPOSX1 DFFPOSX1_540 ( .CLK(clock_i_bF_buf93), .D(_539_), .Q(_3654__7_) );
DFFPOSX1 DFFPOSX1_541 ( .CLK(clock_i_bF_buf30), .D(_540_), .Q(_3654__6_) );
DFFPOSX1 DFFPOSX1_542 ( .CLK(clock_i_bF_buf30), .D(_541_), .Q(_3654__5_) );
DFFPOSX1 DFFPOSX1_543 ( .CLK(clock_i_bF_buf91), .D(_542_), .Q(_3654__4_) );
DFFPOSX1 DFFPOSX1_544 ( .CLK(clock_i_bF_buf73), .D(_543_), .Q(_3654__3_) );
DFFPOSX1 DFFPOSX1_545 ( .CLK(clock_i_bF_buf32), .D(_544_), .Q(_3654__2_) );
DFFPOSX1 DFFPOSX1_546 ( .CLK(clock_i_bF_buf32), .D(_545_), .Q(_3654__1_) );
DFFPOSX1 DFFPOSX1_547 ( .CLK(clock_i_bF_buf73), .D(_546_), .Q(_3654__0_) );
DFFPOSX1 DFFPOSX1_548 ( .CLK(clock_i_bF_buf80), .D(_547_), .Q(_3655__63_) );
DFFPOSX1 DFFPOSX1_549 ( .CLK(clock_i_bF_buf54), .D(_548_), .Q(_3655__62_) );
DFFPOSX1 DFFPOSX1_550 ( .CLK(clock_i_bF_buf22), .D(_549_), .Q(_3655__61_) );
DFFPOSX1 DFFPOSX1_551 ( .CLK(clock_i_bF_buf80), .D(_550_), .Q(_3655__60_) );
DFFPOSX1 DFFPOSX1_552 ( .CLK(clock_i_bF_buf8), .D(_551_), .Q(_3655__59_) );
DFFPOSX1 DFFPOSX1_553 ( .CLK(clock_i_bF_buf61), .D(_552_), .Q(_3655__58_) );
DFFPOSX1 DFFPOSX1_554 ( .CLK(clock_i_bF_buf8), .D(_553_), .Q(_3655__57_) );
DFFPOSX1 DFFPOSX1_555 ( .CLK(clock_i_bF_buf11), .D(_554_), .Q(_3655__56_) );
DFFPOSX1 DFFPOSX1_556 ( .CLK(clock_i_bF_buf89), .D(_555_), .Q(_3655__55_) );
DFFPOSX1 DFFPOSX1_557 ( .CLK(clock_i_bF_buf56), .D(_556_), .Q(_3655__54_) );
DFFPOSX1 DFFPOSX1_558 ( .CLK(clock_i_bF_buf56), .D(_557_), .Q(_3655__53_) );
DFFPOSX1 DFFPOSX1_559 ( .CLK(clock_i_bF_buf57), .D(_558_), .Q(_3655__52_) );
DFFPOSX1 DFFPOSX1_560 ( .CLK(clock_i_bF_buf12), .D(_559_), .Q(_3655__51_) );
DFFPOSX1 DFFPOSX1_561 ( .CLK(clock_i_bF_buf56), .D(_560_), .Q(_3655__50_) );
DFFPOSX1 DFFPOSX1_562 ( .CLK(clock_i_bF_buf56), .D(_561_), .Q(_3655__49_) );
DFFPOSX1 DFFPOSX1_563 ( .CLK(clock_i_bF_buf11), .D(_562_), .Q(_3655__48_) );
DFFPOSX1 DFFPOSX1_564 ( .CLK(clock_i_bF_buf23), .D(_563_), .Q(_3655__47_) );
DFFPOSX1 DFFPOSX1_565 ( .CLK(clock_i_bF_buf14), .D(_564_), .Q(_3655__46_) );
DFFPOSX1 DFFPOSX1_566 ( .CLK(clock_i_bF_buf14), .D(_565_), .Q(_3655__45_) );
DFFPOSX1 DFFPOSX1_567 ( .CLK(clock_i_bF_buf101), .D(_566_), .Q(_3655__44_) );
DFFPOSX1 DFFPOSX1_568 ( .CLK(clock_i_bF_buf14), .D(_567_), .Q(_3655__43_) );
DFFPOSX1 DFFPOSX1_569 ( .CLK(clock_i_bF_buf78), .D(_568_), .Q(_3655__42_) );
DFFPOSX1 DFFPOSX1_570 ( .CLK(clock_i_bF_buf78), .D(_569_), .Q(_3655__41_) );
DFFPOSX1 DFFPOSX1_571 ( .CLK(clock_i_bF_buf58), .D(_570_), .Q(_3655__40_) );
DFFPOSX1 DFFPOSX1_572 ( .CLK(clock_i_bF_buf39), .D(_571_), .Q(_3655__39_) );
DFFPOSX1 DFFPOSX1_573 ( .CLK(clock_i_bF_buf42), .D(_572_), .Q(_3655__38_) );
DFFPOSX1 DFFPOSX1_574 ( .CLK(clock_i_bF_buf39), .D(_573_), .Q(_3655__37_) );
DFFPOSX1 DFFPOSX1_575 ( .CLK(clock_i_bF_buf101), .D(_574_), .Q(_3655__36_) );
DFFPOSX1 DFFPOSX1_576 ( .CLK(clock_i_bF_buf14), .D(_575_), .Q(_3655__35_) );
DFFPOSX1 DFFPOSX1_577 ( .CLK(clock_i_bF_buf39), .D(_576_), .Q(_3655__34_) );
DFFPOSX1 DFFPOSX1_578 ( .CLK(clock_i_bF_buf101), .D(_577_), .Q(_3655__33_) );
DFFPOSX1 DFFPOSX1_579 ( .CLK(clock_i_bF_buf42), .D(_578_), .Q(_3655__32_) );
DFFPOSX1 DFFPOSX1_580 ( .CLK(clock_i_bF_buf93), .D(_579_), .Q(_3655__31_) );
DFFPOSX1 DFFPOSX1_581 ( .CLK(clock_i_bF_buf78), .D(_580_), .Q(_3655__30_) );
DFFPOSX1 DFFPOSX1_582 ( .CLK(clock_i_bF_buf93), .D(_581_), .Q(_3655__29_) );
DFFPOSX1 DFFPOSX1_583 ( .CLK(clock_i_bF_buf83), .D(_582_), .Q(_3655__28_) );
DFFPOSX1 DFFPOSX1_584 ( .CLK(clock_i_bF_buf93), .D(_583_), .Q(_3655__27_) );
DFFPOSX1 DFFPOSX1_585 ( .CLK(clock_i_bF_buf79), .D(_584_), .Q(_3655__26_) );
DFFPOSX1 DFFPOSX1_586 ( .CLK(clock_i_bF_buf14), .D(_585_), .Q(_3655__25_) );
DFFPOSX1 DFFPOSX1_587 ( .CLK(clock_i_bF_buf93), .D(_586_), .Q(_3655__24_) );
DFFPOSX1 DFFPOSX1_588 ( .CLK(clock_i_bF_buf101), .D(_587_), .Q(_3655__23_) );
DFFPOSX1 DFFPOSX1_589 ( .CLK(clock_i_bF_buf22), .D(_588_), .Q(_3655__22_) );
DFFPOSX1 DFFPOSX1_590 ( .CLK(clock_i_bF_buf22), .D(_589_), .Q(_3655__21_) );
DFFPOSX1 DFFPOSX1_591 ( .CLK(clock_i_bF_buf2), .D(_590_), .Q(_3655__20_) );
DFFPOSX1 DFFPOSX1_592 ( .CLK(clock_i_bF_buf18), .D(_591_), .Q(_3655__19_) );
DFFPOSX1 DFFPOSX1_593 ( .CLK(clock_i_bF_buf78), .D(_592_), .Q(_3655__18_) );
DFFPOSX1 DFFPOSX1_594 ( .CLK(clock_i_bF_buf12), .D(_593_), .Q(_3655__17_) );
DFFPOSX1 DFFPOSX1_595 ( .CLK(clock_i_bF_buf30), .D(_594_), .Q(_3655__16_) );
DFFPOSX1 DFFPOSX1_596 ( .CLK(clock_i_bF_buf2), .D(_595_), .Q(_3655__15_) );
DFFPOSX1 DFFPOSX1_597 ( .CLK(clock_i_bF_buf23), .D(_596_), .Q(_3655__14_) );
DFFPOSX1 DFFPOSX1_598 ( .CLK(clock_i_bF_buf2), .D(_597_), .Q(_3655__13_) );
DFFPOSX1 DFFPOSX1_599 ( .CLK(clock_i_bF_buf30), .D(_598_), .Q(_3655__12_) );
DFFPOSX1 DFFPOSX1_600 ( .CLK(clock_i_bF_buf30), .D(_599_), .Q(_3655__11_) );
DFFPOSX1 DFFPOSX1_601 ( .CLK(clock_i_bF_buf78), .D(_600_), .Q(_3655__10_) );
DFFPOSX1 DFFPOSX1_602 ( .CLK(clock_i_bF_buf23), .D(_601_), .Q(_3655__9_) );
DFFPOSX1 DFFPOSX1_603 ( .CLK(clock_i_bF_buf42), .D(_602_), .Q(_3655__8_) );
DFFPOSX1 DFFPOSX1_604 ( .CLK(clock_i_bF_buf52), .D(_603_), .Q(_3655__7_) );
DFFPOSX1 DFFPOSX1_605 ( .CLK(clock_i_bF_buf83), .D(_604_), .Q(_3655__6_) );
DFFPOSX1 DFFPOSX1_606 ( .CLK(clock_i_bF_buf97), .D(_605_), .Q(_3655__5_) );
DFFPOSX1 DFFPOSX1_607 ( .CLK(clock_i_bF_buf83), .D(_606_), .Q(_3655__4_) );
DFFPOSX1 DFFPOSX1_608 ( .CLK(clock_i_bF_buf78), .D(_607_), .Q(_3655__3_) );
DFFPOSX1 DFFPOSX1_609 ( .CLK(clock_i_bF_buf73), .D(_608_), .Q(_3655__2_) );
DFFPOSX1 DFFPOSX1_610 ( .CLK(clock_i_bF_buf73), .D(_609_), .Q(_3655__1_) );
DFFPOSX1 DFFPOSX1_611 ( .CLK(clock_i_bF_buf93), .D(_610_), .Q(_3655__0_) );
DFFPOSX1 DFFPOSX1_612 ( .CLK(clock_i_bF_buf92), .D(enable_i_bF_buf6), .Q(_3640_) );
DFFPOSX1 DFFPOSX1_613 ( .CLK(clock_i_bF_buf35), .D(_611__bF_buf2), .Q(_3641_) );
DFFPOSX1 DFFPOSX1_614 ( .CLK(clock_i_bF_buf26), .D(_612__bF_buf2), .Q(_3642_) );
DFFPOSX1 DFFPOSX1_615 ( .CLK(clock_i_bF_buf35), .D(_613__bF_buf4), .Q(_3643_) );
DFFPOSX1 DFFPOSX1_616 ( .CLK(clock_i_bF_buf20), .D(_614_), .Q(_3644__31_) );
DFFPOSX1 DFFPOSX1_617 ( .CLK(clock_i_bF_buf15), .D(_615_), .Q(_3644__30_) );
DFFPOSX1 DFFPOSX1_618 ( .CLK(clock_i_bF_buf21), .D(_616_), .Q(_3644__29_) );
DFFPOSX1 DFFPOSX1_619 ( .CLK(clock_i_bF_buf96), .D(_617_), .Q(_3644__28_) );
DFFPOSX1 DFFPOSX1_620 ( .CLK(clock_i_bF_buf48), .D(_618_), .Q(_3644__27_) );
DFFPOSX1 DFFPOSX1_621 ( .CLK(clock_i_bF_buf24), .D(_619_), .Q(_3644__26_) );
DFFPOSX1 DFFPOSX1_622 ( .CLK(clock_i_bF_buf96), .D(_620_), .Q(_3644__25_) );
DFFPOSX1 DFFPOSX1_623 ( .CLK(clock_i_bF_buf44), .D(_621_), .Q(_3644__24_) );
DFFPOSX1 DFFPOSX1_624 ( .CLK(clock_i_bF_buf41), .D(_622_), .Q(_3644__23_) );
DFFPOSX1 DFFPOSX1_625 ( .CLK(clock_i_bF_buf92), .D(_623_), .Q(_3644__22_) );
DFFPOSX1 DFFPOSX1_626 ( .CLK(clock_i_bF_buf48), .D(_624_), .Q(_3644__21_) );
DFFPOSX1 DFFPOSX1_627 ( .CLK(clock_i_bF_buf35), .D(_625_), .Q(_3644__20_) );
DFFPOSX1 DFFPOSX1_628 ( .CLK(clock_i_bF_buf31), .D(_626_), .Q(_3644__19_) );
DFFPOSX1 DFFPOSX1_629 ( .CLK(clock_i_bF_buf20), .D(_627_), .Q(_3644__18_) );
DFFPOSX1 DFFPOSX1_630 ( .CLK(clock_i_bF_buf41), .D(_628_), .Q(_3644__17_) );
DFFPOSX1 DFFPOSX1_631 ( .CLK(clock_i_bF_buf92), .D(_629_), .Q(_3644__16_) );
DFFPOSX1 DFFPOSX1_632 ( .CLK(clock_i_bF_buf41), .D(_630_), .Q(_3644__15_) );
DFFPOSX1 DFFPOSX1_633 ( .CLK(clock_i_bF_buf41), .D(_631_), .Q(_3644__14_) );
DFFPOSX1 DFFPOSX1_634 ( .CLK(clock_i_bF_buf88), .D(_632_), .Q(_3644__13_) );
DFFPOSX1 DFFPOSX1_635 ( .CLK(clock_i_bF_buf20), .D(_633_), .Q(_3644__12_) );
DFFPOSX1 DFFPOSX1_636 ( .CLK(clock_i_bF_buf6), .D(_634_), .Q(_3644__11_) );
DFFPOSX1 DFFPOSX1_637 ( .CLK(clock_i_bF_buf92), .D(_635_), .Q(_3644__10_) );
DFFPOSX1 DFFPOSX1_638 ( .CLK(clock_i_bF_buf20), .D(_636_), .Q(_3644__9_) );
DFFPOSX1 DFFPOSX1_639 ( .CLK(clock_i_bF_buf6), .D(_637_), .Q(_3644__8_) );
DFFPOSX1 DFFPOSX1_640 ( .CLK(clock_i_bF_buf3), .D(_638_), .Q(_3644__7_) );
DFFPOSX1 DFFPOSX1_641 ( .CLK(clock_i_bF_buf20), .D(_639_), .Q(_3644__6_) );
DFFPOSX1 DFFPOSX1_642 ( .CLK(clock_i_bF_buf20), .D(_640_), .Q(_3644__5_) );
DFFPOSX1 DFFPOSX1_643 ( .CLK(clock_i_bF_buf31), .D(_641_), .Q(_3644__4_) );
DFFPOSX1 DFFPOSX1_644 ( .CLK(clock_i_bF_buf92), .D(_642_), .Q(_3644__3_) );
DFFPOSX1 DFFPOSX1_645 ( .CLK(clock_i_bF_buf6), .D(_643_), .Q(_3644__2_) );
DFFPOSX1 DFFPOSX1_646 ( .CLK(clock_i_bF_buf48), .D(_644_), .Q(_3644__1_) );
DFFPOSX1 DFFPOSX1_647 ( .CLK(clock_i_bF_buf48), .D(_645_), .Q(_3644__0_) );
DFFPOSX1 DFFPOSX1_648 ( .CLK(clock_i_bF_buf98), .D(_646_), .Q(_3645__31_) );
DFFPOSX1 DFFPOSX1_649 ( .CLK(clock_i_bF_buf38), .D(_647_), .Q(_3645__30_) );
DFFPOSX1 DFFPOSX1_650 ( .CLK(clock_i_bF_buf24), .D(_648_), .Q(_3645__29_) );
DFFPOSX1 DFFPOSX1_651 ( .CLK(clock_i_bF_buf70), .D(_649_), .Q(_3645__28_) );
DFFPOSX1 DFFPOSX1_652 ( .CLK(clock_i_bF_buf61), .D(_650_), .Q(_3645__27_) );
DFFPOSX1 DFFPOSX1_653 ( .CLK(clock_i_bF_buf20), .D(_651_), .Q(_3645__26_) );
DFFPOSX1 DFFPOSX1_654 ( .CLK(clock_i_bF_buf70), .D(_652_), .Q(_3645__25_) );
DFFPOSX1 DFFPOSX1_655 ( .CLK(clock_i_bF_buf6), .D(_653_), .Q(_3645__24_) );
DFFPOSX1 DFFPOSX1_656 ( .CLK(clock_i_bF_buf63), .D(_654_), .Q(_3645__23_) );
DFFPOSX1 DFFPOSX1_657 ( .CLK(clock_i_bF_buf48), .D(_655_), .Q(_3645__22_) );
DFFPOSX1 DFFPOSX1_658 ( .CLK(clock_i_bF_buf50), .D(_656_), .Q(_3645__21_) );
DFFPOSX1 DFFPOSX1_659 ( .CLK(clock_i_bF_buf48), .D(_657_), .Q(_3645__20_) );
DFFPOSX1 DFFPOSX1_660 ( .CLK(clock_i_bF_buf60), .D(_658_), .Q(_3645__19_) );
DFFPOSX1 DFFPOSX1_661 ( .CLK(clock_i_bF_buf70), .D(_659_), .Q(_3645__18_) );
DFFPOSX1 DFFPOSX1_662 ( .CLK(clock_i_bF_buf63), .D(_660_), .Q(_3645__17_) );
DFFPOSX1 DFFPOSX1_663 ( .CLK(clock_i_bF_buf20), .D(_661_), .Q(_3645__16_) );
DFFPOSX1 DFFPOSX1_664 ( .CLK(clock_i_bF_buf6), .D(_662_), .Q(_3645__15_) );
DFFPOSX1 DFFPOSX1_665 ( .CLK(clock_i_bF_buf27), .D(_663_), .Q(_3645__14_) );
DFFPOSX1 DFFPOSX1_666 ( .CLK(clock_i_bF_buf44), .D(_664_), .Q(_3645__13_) );
DFFPOSX1 DFFPOSX1_667 ( .CLK(clock_i_bF_buf51), .D(_665_), .Q(_3645__12_) );
DFFPOSX1 DFFPOSX1_668 ( .CLK(clock_i_bF_buf6), .D(_666_), .Q(_3645__11_) );
DFFPOSX1 DFFPOSX1_669 ( .CLK(clock_i_bF_buf21), .D(_667_), .Q(_3645__10_) );
DFFPOSX1 DFFPOSX1_670 ( .CLK(clock_i_bF_buf7), .D(_668_), .Q(_3645__9_) );
DFFPOSX1 DFFPOSX1_671 ( .CLK(clock_i_bF_buf92), .D(_669_), .Q(_3645__8_) );
DFFPOSX1 DFFPOSX1_672 ( .CLK(clock_i_bF_buf1), .D(_670_), .Q(_3645__7_) );
DFFPOSX1 DFFPOSX1_673 ( .CLK(clock_i_bF_buf20), .D(_671_), .Q(_3645__6_) );
DFFPOSX1 DFFPOSX1_674 ( .CLK(clock_i_bF_buf48), .D(_672_), .Q(_3645__5_) );
DFFPOSX1 DFFPOSX1_675 ( .CLK(clock_i_bF_buf89), .D(_673_), .Q(_3645__4_) );
DFFPOSX1 DFFPOSX1_676 ( .CLK(clock_i_bF_buf49), .D(_674_), .Q(_3645__3_) );
DFFPOSX1 DFFPOSX1_677 ( .CLK(clock_i_bF_buf21), .D(_675_), .Q(_3645__2_) );
DFFPOSX1 DFFPOSX1_678 ( .CLK(clock_i_bF_buf51), .D(_676_), .Q(_3645__1_) );
DFFPOSX1 DFFPOSX1_679 ( .CLK(clock_i_bF_buf6), .D(_677_), .Q(_3645__0_) );
DFFPOSX1 DFFPOSX1_680 ( .CLK(clock_i_bF_buf1), .D(_678_), .Q(_3646__31_) );
DFFPOSX1 DFFPOSX1_681 ( .CLK(clock_i_bF_buf60), .D(_679_), .Q(_3646__30_) );
DFFPOSX1 DFFPOSX1_682 ( .CLK(clock_i_bF_buf46), .D(_680_), .Q(_3646__29_) );
DFFPOSX1 DFFPOSX1_683 ( .CLK(clock_i_bF_buf63), .D(_681_), .Q(_3646__28_) );
DFFPOSX1 DFFPOSX1_684 ( .CLK(clock_i_bF_buf65), .D(_682_), .Q(_3646__27_) );
DFFPOSX1 DFFPOSX1_685 ( .CLK(clock_i_bF_buf44), .D(_683_), .Q(_3646__26_) );
DFFPOSX1 DFFPOSX1_686 ( .CLK(clock_i_bF_buf65), .D(_684_), .Q(_3646__25_) );
DFFPOSX1 DFFPOSX1_687 ( .CLK(clock_i_bF_buf62), .D(_685_), .Q(_3646__24_) );
DFFPOSX1 DFFPOSX1_688 ( .CLK(clock_i_bF_buf41), .D(_686_), .Q(_3646__23_) );
DFFPOSX1 DFFPOSX1_689 ( .CLK(clock_i_bF_buf50), .D(_687_), .Q(_3646__22_) );
DFFPOSX1 DFFPOSX1_690 ( .CLK(clock_i_bF_buf63), .D(_688_), .Q(_3646__21_) );
DFFPOSX1 DFFPOSX1_691 ( .CLK(clock_i_bF_buf70), .D(_689_), .Q(_3646__20_) );
DFFPOSX1 DFFPOSX1_692 ( .CLK(clock_i_bF_buf41), .D(_690_), .Q(_3646__19_) );
DFFPOSX1 DFFPOSX1_693 ( .CLK(clock_i_bF_buf48), .D(_691_), .Q(_3646__18_) );
DFFPOSX1 DFFPOSX1_694 ( .CLK(clock_i_bF_buf6), .D(_692_), .Q(_3646__17_) );
DFFPOSX1 DFFPOSX1_695 ( .CLK(clock_i_bF_buf62), .D(_693_), .Q(_3646__16_) );
DFFPOSX1 DFFPOSX1_696 ( .CLK(clock_i_bF_buf62), .D(_694_), .Q(_3646__15_) );
DFFPOSX1 DFFPOSX1_697 ( .CLK(clock_i_bF_buf50), .D(_695_), .Q(_3646__14_) );
DFFPOSX1 DFFPOSX1_698 ( .CLK(clock_i_bF_buf6), .D(_696_), .Q(_3646__13_) );
DFFPOSX1 DFFPOSX1_699 ( .CLK(clock_i_bF_buf65), .D(_697_), .Q(_3646__12_) );
DFFPOSX1 DFFPOSX1_700 ( .CLK(clock_i_bF_buf77), .D(_698_), .Q(_3646__11_) );
DFFPOSX1 DFFPOSX1_701 ( .CLK(clock_i_bF_buf71), .D(_699_), .Q(_3646__10_) );
DFFPOSX1 DFFPOSX1_702 ( .CLK(clock_i_bF_buf62), .D(_700_), .Q(_3646__9_) );
DFFPOSX1 DFFPOSX1_703 ( .CLK(clock_i_bF_buf100), .D(_701_), .Q(_3646__8_) );
DFFPOSX1 DFFPOSX1_704 ( .CLK(clock_i_bF_buf6), .D(_702_), .Q(_3646__7_) );
DFFPOSX1 DFFPOSX1_705 ( .CLK(clock_i_bF_buf65), .D(_703_), .Q(_3646__6_) );
DFFPOSX1 DFFPOSX1_706 ( .CLK(clock_i_bF_buf48), .D(_704_), .Q(_3646__5_) );
DFFPOSX1 DFFPOSX1_707 ( .CLK(clock_i_bF_buf48), .D(_705_), .Q(_3646__4_) );
DFFPOSX1 DFFPOSX1_708 ( .CLK(clock_i_bF_buf96), .D(_706_), .Q(_3646__3_) );
DFFPOSX1 DFFPOSX1_709 ( .CLK(clock_i_bF_buf46), .D(_707_), .Q(_3646__2_) );
DFFPOSX1 DFFPOSX1_710 ( .CLK(clock_i_bF_buf3), .D(_708_), .Q(_3646__1_) );
DFFPOSX1 DFFPOSX1_711 ( .CLK(clock_i_bF_buf7), .D(_709_), .Q(_3646__0_) );
DFFPOSX1 DFFPOSX1_712 ( .CLK(clock_i_bF_buf100), .D(_710_), .Q(_3647__31_) );
DFFPOSX1 DFFPOSX1_713 ( .CLK(clock_i_bF_buf85), .D(_711_), .Q(_3647__30_) );
DFFPOSX1 DFFPOSX1_714 ( .CLK(clock_i_bF_buf76), .D(_712_), .Q(_3647__29_) );
DFFPOSX1 DFFPOSX1_715 ( .CLK(clock_i_bF_buf0), .D(_713_), .Q(_3647__28_) );
DFFPOSX1 DFFPOSX1_716 ( .CLK(clock_i_bF_buf81), .D(_714_), .Q(_3647__27_) );
DFFPOSX1 DFFPOSX1_717 ( .CLK(clock_i_bF_buf40), .D(_715_), .Q(_3647__26_) );
DFFPOSX1 DFFPOSX1_718 ( .CLK(clock_i_bF_buf85), .D(_716_), .Q(_3647__25_) );
DFFPOSX1 DFFPOSX1_719 ( .CLK(clock_i_bF_buf31), .D(_717_), .Q(_3647__24_) );
DFFPOSX1 DFFPOSX1_720 ( .CLK(clock_i_bF_buf87), .D(_718_), .Q(_3647__23_) );
DFFPOSX1 DFFPOSX1_721 ( .CLK(clock_i_bF_buf4), .D(_719_), .Q(_3647__22_) );
DFFPOSX1 DFFPOSX1_722 ( .CLK(clock_i_bF_buf41), .D(_720_), .Q(_3647__21_) );
DFFPOSX1 DFFPOSX1_723 ( .CLK(clock_i_bF_buf10), .D(_721_), .Q(_3647__20_) );
DFFPOSX1 DFFPOSX1_724 ( .CLK(clock_i_bF_buf44), .D(_722_), .Q(_3647__19_) );
DFFPOSX1 DFFPOSX1_725 ( .CLK(clock_i_bF_buf59), .D(_723_), .Q(_3647__18_) );
DFFPOSX1 DFFPOSX1_726 ( .CLK(clock_i_bF_buf21), .D(_724_), .Q(_3647__17_) );
DFFPOSX1 DFFPOSX1_727 ( .CLK(clock_i_bF_buf64), .D(_725_), .Q(_3647__16_) );
DFFPOSX1 DFFPOSX1_728 ( .CLK(clock_i_bF_buf64), .D(_726_), .Q(_3647__15_) );
DFFPOSX1 DFFPOSX1_729 ( .CLK(clock_i_bF_buf24), .D(_727_), .Q(_3647__14_) );
DFFPOSX1 DFFPOSX1_730 ( .CLK(clock_i_bF_buf46), .D(_728_), .Q(_3647__13_) );
DFFPOSX1 DFFPOSX1_731 ( .CLK(clock_i_bF_buf21), .D(_729_), .Q(_3647__12_) );
DFFPOSX1 DFFPOSX1_732 ( .CLK(clock_i_bF_buf31), .D(_730_), .Q(_3647__11_) );
DFFPOSX1 DFFPOSX1_733 ( .CLK(clock_i_bF_buf25), .D(_731_), .Q(_3647__10_) );
DFFPOSX1 DFFPOSX1_734 ( .CLK(clock_i_bF_buf19), .D(_732_), .Q(_3647__9_) );
DFFPOSX1 DFFPOSX1_735 ( .CLK(clock_i_bF_buf29), .D(_733_), .Q(_3647__8_) );
DFFPOSX1 DFFPOSX1_736 ( .CLK(clock_i_bF_buf41), .D(_734_), .Q(_3647__7_) );
DFFPOSX1 DFFPOSX1_737 ( .CLK(clock_i_bF_buf38), .D(_735_), .Q(_3647__6_) );
DFFPOSX1 DFFPOSX1_738 ( .CLK(clock_i_bF_buf65), .D(_736_), .Q(_3647__5_) );
DFFPOSX1 DFFPOSX1_739 ( .CLK(clock_i_bF_buf46), .D(_737_), .Q(_3647__4_) );
DFFPOSX1 DFFPOSX1_740 ( .CLK(clock_i_bF_buf43), .D(_738_), .Q(_3647__3_) );
DFFPOSX1 DFFPOSX1_741 ( .CLK(clock_i_bF_buf85), .D(_739_), .Q(_3647__2_) );
DFFPOSX1 DFFPOSX1_742 ( .CLK(clock_i_bF_buf45), .D(_740_), .Q(_3647__1_) );
DFFPOSX1 DFFPOSX1_743 ( .CLK(clock_i_bF_buf64), .D(_741_), .Q(_3647__0_) );
DFFPOSX1 DFFPOSX1_744 ( .CLK(clock_i_bF_buf85), .D(_742_), .Q(_3636__63_) );
DFFPOSX1 DFFPOSX1_745 ( .CLK(clock_i_bF_buf29), .D(_743_), .Q(_3636__62_) );
DFFPOSX1 DFFPOSX1_746 ( .CLK(clock_i_bF_buf90), .D(_744_), .Q(_3636__61_) );
DFFPOSX1 DFFPOSX1_747 ( .CLK(clock_i_bF_buf28), .D(_745_), .Q(_3636__60_) );
DFFPOSX1 DFFPOSX1_748 ( .CLK(clock_i_bF_buf71), .D(_746_), .Q(_3636__59_) );
DFFPOSX1 DFFPOSX1_749 ( .CLK(clock_i_bF_buf71), .D(_747_), .Q(_3636__58_) );
DFFPOSX1 DFFPOSX1_750 ( .CLK(clock_i_bF_buf71), .D(_748_), .Q(_3636__57_) );
DFFPOSX1 DFFPOSX1_751 ( .CLK(clock_i_bF_buf90), .D(_749_), .Q(_3636__56_) );
DFFPOSX1 DFFPOSX1_752 ( .CLK(clock_i_bF_buf90), .D(_750_), .Q(_3636__55_) );
DFFPOSX1 DFFPOSX1_753 ( .CLK(clock_i_bF_buf90), .D(_751_), .Q(_3636__54_) );
DFFPOSX1 DFFPOSX1_754 ( .CLK(clock_i_bF_buf97), .D(_752_), .Q(_3636__53_) );
DFFPOSX1 DFFPOSX1_755 ( .CLK(clock_i_bF_buf37), .D(_753_), .Q(_3636__52_) );
DFFPOSX1 DFFPOSX1_756 ( .CLK(clock_i_bF_buf37), .D(_754_), .Q(_3636__51_) );
DFFPOSX1 DFFPOSX1_757 ( .CLK(clock_i_bF_buf32), .D(_755_), .Q(_3636__50_) );
DFFPOSX1 DFFPOSX1_758 ( .CLK(clock_i_bF_buf43), .D(_756_), .Q(_3636__49_) );
DFFPOSX1 DFFPOSX1_759 ( .CLK(clock_i_bF_buf43), .D(_757_), .Q(_3636__48_) );
DFFPOSX1 DFFPOSX1_760 ( .CLK(clock_i_bF_buf79), .D(_758_), .Q(_3636__47_) );
DFFPOSX1 DFFPOSX1_761 ( .CLK(clock_i_bF_buf0), .D(_759_), .Q(_3636__46_) );
DFFPOSX1 DFFPOSX1_762 ( .CLK(clock_i_bF_buf47), .D(_760_), .Q(_3636__45_) );
DFFPOSX1 DFFPOSX1_763 ( .CLK(clock_i_bF_buf42), .D(_761_), .Q(_3636__44_) );
DFFPOSX1 DFFPOSX1_764 ( .CLK(clock_i_bF_buf19), .D(_762_), .Q(_3636__43_) );
DFFPOSX1 DFFPOSX1_765 ( .CLK(clock_i_bF_buf19), .D(_763_), .Q(_3636__42_) );
DFFPOSX1 DFFPOSX1_766 ( .CLK(clock_i_bF_buf51), .D(_764_), .Q(_3636__41_) );
DFFPOSX1 DFFPOSX1_767 ( .CLK(clock_i_bF_buf50), .D(_765_), .Q(_3636__40_) );
DFFPOSX1 DFFPOSX1_768 ( .CLK(clock_i_bF_buf19), .D(_766_), .Q(_3636__39_) );
DFFPOSX1 DFFPOSX1_769 ( .CLK(clock_i_bF_buf42), .D(_767_), .Q(_3636__38_) );
DFFPOSX1 DFFPOSX1_770 ( .CLK(clock_i_bF_buf67), .D(_768_), .Q(_3636__37_) );
DFFPOSX1 DFFPOSX1_771 ( .CLK(clock_i_bF_buf47), .D(_769_), .Q(_3636__36_) );
DFFPOSX1 DFFPOSX1_772 ( .CLK(clock_i_bF_buf47), .D(_770_), .Q(_3636__35_) );
DFFPOSX1 DFFPOSX1_773 ( .CLK(clock_i_bF_buf95), .D(_771_), .Q(_3636__34_) );
DFFPOSX1 DFFPOSX1_774 ( .CLK(clock_i_bF_buf88), .D(_772_), .Q(_3636__33_) );
DFFPOSX1 DFFPOSX1_775 ( .CLK(clock_i_bF_buf13), .D(_773_), .Q(_3636__32_) );
DFFPOSX1 DFFPOSX1_776 ( .CLK(clock_i_bF_buf13), .D(_774_), .Q(_3636__31_) );
DFFPOSX1 DFFPOSX1_777 ( .CLK(clock_i_bF_buf13), .D(_775_), .Q(_3636__30_) );
DFFPOSX1 DFFPOSX1_778 ( .CLK(clock_i_bF_buf53), .D(_776_), .Q(_3636__29_) );
DFFPOSX1 DFFPOSX1_779 ( .CLK(clock_i_bF_buf40), .D(_777_), .Q(_3636__28_) );
DFFPOSX1 DFFPOSX1_780 ( .CLK(clock_i_bF_buf74), .D(_778_), .Q(_3636__27_) );
DFFPOSX1 DFFPOSX1_781 ( .CLK(clock_i_bF_buf25), .D(_779_), .Q(_3636__26_) );
DFFPOSX1 DFFPOSX1_782 ( .CLK(clock_i_bF_buf49), .D(_780_), .Q(_3636__25_) );
DFFPOSX1 DFFPOSX1_783 ( .CLK(clock_i_bF_buf49), .D(_781_), .Q(_3636__24_) );
DFFPOSX1 DFFPOSX1_784 ( .CLK(clock_i_bF_buf49), .D(_782_), .Q(_3636__23_) );
DFFPOSX1 DFFPOSX1_785 ( .CLK(clock_i_bF_buf49), .D(_783_), .Q(_3636__22_) );
DFFPOSX1 DFFPOSX1_786 ( .CLK(clock_i_bF_buf66), .D(_784_), .Q(_3636__21_) );
DFFPOSX1 DFFPOSX1_787 ( .CLK(clock_i_bF_buf53), .D(_785_), .Q(_3636__20_) );
DFFPOSX1 DFFPOSX1_788 ( .CLK(clock_i_bF_buf81), .D(_786_), .Q(_3636__19_) );
DFFPOSX1 DFFPOSX1_789 ( .CLK(clock_i_bF_buf34), .D(_787_), .Q(_3636__18_) );
DFFPOSX1 DFFPOSX1_790 ( .CLK(clock_i_bF_buf72), .D(_788_), .Q(_3636__17_) );
DFFPOSX1 DFFPOSX1_791 ( .CLK(clock_i_bF_buf72), .D(_789_), .Q(_3636__16_) );
DFFPOSX1 DFFPOSX1_792 ( .CLK(clock_i_bF_buf35), .D(_790_), .Q(_3636__15_) );
DFFPOSX1 DFFPOSX1_793 ( .CLK(clock_i_bF_buf34), .D(_791_), .Q(_3636__14_) );
DFFPOSX1 DFFPOSX1_794 ( .CLK(clock_i_bF_buf26), .D(_792_), .Q(_3636__13_) );
DFFPOSX1 DFFPOSX1_795 ( .CLK(clock_i_bF_buf26), .D(_793_), .Q(_3636__12_) );
DFFPOSX1 DFFPOSX1_796 ( .CLK(clock_i_bF_buf26), .D(_794_), .Q(_3636__11_) );
DFFPOSX1 DFFPOSX1_797 ( .CLK(clock_i_bF_buf64), .D(_795_), .Q(_3636__10_) );
DFFPOSX1 DFFPOSX1_798 ( .CLK(clock_i_bF_buf65), .D(_796_), .Q(_3636__9_) );
DFFPOSX1 DFFPOSX1_799 ( .CLK(clock_i_bF_buf82), .D(_797_), .Q(_3636__8_) );
DFFPOSX1 DFFPOSX1_800 ( .CLK(clock_i_bF_buf31), .D(_798_), .Q(_3636__7_) );
DFFPOSX1 DFFPOSX1_801 ( .CLK(clock_i_bF_buf31), .D(_799_), .Q(_3636__6_) );
DFFPOSX1 DFFPOSX1_802 ( .CLK(clock_i_bF_buf5), .D(_800_), .Q(_3636__5_) );
DFFPOSX1 DFFPOSX1_803 ( .CLK(clock_i_bF_buf5), .D(_801_), .Q(_3636__4_) );
DFFPOSX1 DFFPOSX1_804 ( .CLK(clock_i_bF_buf33), .D(_802_), .Q(_3636__3_) );
DFFPOSX1 DFFPOSX1_805 ( .CLK(clock_i_bF_buf82), .D(_803_), .Q(_3636__2_) );
DFFPOSX1 DFFPOSX1_806 ( .CLK(clock_i_bF_buf72), .D(_804_), .Q(_3636__1_) );
DFFPOSX1 DFFPOSX1_807 ( .CLK(clock_i_bF_buf72), .D(_805_), .Q(_3636__0_) );
DFFPOSX1 DFFPOSX1_808 ( .CLK(clock_i_bF_buf85), .D(_806_), .Q(_3637__63_) );
DFFPOSX1 DFFPOSX1_809 ( .CLK(clock_i_bF_buf24), .D(_807_), .Q(_3637__62_) );
DFFPOSX1 DFFPOSX1_810 ( .CLK(clock_i_bF_buf1), .D(_808_), .Q(_3637__61_) );
DFFPOSX1 DFFPOSX1_811 ( .CLK(clock_i_bF_buf95), .D(_809_), .Q(_3637__60_) );
DFFPOSX1 DFFPOSX1_812 ( .CLK(clock_i_bF_buf1), .D(_810_), .Q(_3637__59_) );
DFFPOSX1 DFFPOSX1_813 ( .CLK(clock_i_bF_buf90), .D(_811_), .Q(_3637__58_) );
DFFPOSX1 DFFPOSX1_814 ( .CLK(clock_i_bF_buf90), .D(_812_), .Q(_3637__57_) );
DFFPOSX1 DFFPOSX1_815 ( .CLK(clock_i_bF_buf1), .D(_813_), .Q(_3637__56_) );
DFFPOSX1 DFFPOSX1_816 ( .CLK(clock_i_bF_buf28), .D(_814_), .Q(_3637__55_) );
DFFPOSX1 DFFPOSX1_817 ( .CLK(clock_i_bF_buf18), .D(_815_), .Q(_3637__54_) );
DFFPOSX1 DFFPOSX1_818 ( .CLK(clock_i_bF_buf73), .D(_816_), .Q(_3637__53_) );
DFFPOSX1 DFFPOSX1_819 ( .CLK(clock_i_bF_buf97), .D(_817_), .Q(_3637__52_) );
DFFPOSX1 DFFPOSX1_820 ( .CLK(clock_i_bF_buf91), .D(_818_), .Q(_3637__51_) );
DFFPOSX1 DFFPOSX1_821 ( .CLK(clock_i_bF_buf37), .D(_819_), .Q(_3637__50_) );
DFFPOSX1 DFFPOSX1_822 ( .CLK(clock_i_bF_buf32), .D(_820_), .Q(_3637__49_) );
DFFPOSX1 DFFPOSX1_823 ( .CLK(clock_i_bF_buf43), .D(_821_), .Q(_3637__48_) );
DFFPOSX1 DFFPOSX1_824 ( .CLK(clock_i_bF_buf79), .D(_822_), .Q(_3637__47_) );
DFFPOSX1 DFFPOSX1_825 ( .CLK(clock_i_bF_buf79), .D(_823_), .Q(_3637__46_) );
DFFPOSX1 DFFPOSX1_826 ( .CLK(clock_i_bF_buf68), .D(_824_), .Q(_3637__45_) );
DFFPOSX1 DFFPOSX1_827 ( .CLK(clock_i_bF_buf50), .D(_825_), .Q(_3637__44_) );
DFFPOSX1 DFFPOSX1_828 ( .CLK(clock_i_bF_buf68), .D(_826_), .Q(_3637__43_) );
DFFPOSX1 DFFPOSX1_829 ( .CLK(clock_i_bF_buf68), .D(_827_), .Q(_3637__42_) );
DFFPOSX1 DFFPOSX1_830 ( .CLK(clock_i_bF_buf50), .D(_828_), .Q(_3637__41_) );
DFFPOSX1 DFFPOSX1_831 ( .CLK(clock_i_bF_buf68), .D(_829_), .Q(_3637__40_) );
DFFPOSX1 DFFPOSX1_832 ( .CLK(clock_i_bF_buf88), .D(_830_), .Q(_3637__39_) );
DFFPOSX1 DFFPOSX1_833 ( .CLK(clock_i_bF_buf86), .D(_831_), .Q(_3637__38_) );
DFFPOSX1 DFFPOSX1_834 ( .CLK(clock_i_bF_buf47), .D(_832_), .Q(_3637__37_) );
DFFPOSX1 DFFPOSX1_835 ( .CLK(clock_i_bF_buf95), .D(_833_), .Q(_3637__36_) );
DFFPOSX1 DFFPOSX1_836 ( .CLK(clock_i_bF_buf52), .D(_834_), .Q(_3637__35_) );
DFFPOSX1 DFFPOSX1_837 ( .CLK(clock_i_bF_buf75), .D(_835_), .Q(_3637__34_) );
DFFPOSX1 DFFPOSX1_838 ( .CLK(clock_i_bF_buf75), .D(_836_), .Q(_3637__33_) );
DFFPOSX1 DFFPOSX1_839 ( .CLK(clock_i_bF_buf13), .D(_837_), .Q(_3637__32_) );
DFFPOSX1 DFFPOSX1_840 ( .CLK(clock_i_bF_buf13), .D(_838_), .Q(_3637__31_) );
DFFPOSX1 DFFPOSX1_841 ( .CLK(clock_i_bF_buf7), .D(_839_), .Q(_3637__30_) );
DFFPOSX1 DFFPOSX1_842 ( .CLK(clock_i_bF_buf74), .D(_840_), .Q(_3637__29_) );
DFFPOSX1 DFFPOSX1_843 ( .CLK(clock_i_bF_buf40), .D(_841_), .Q(_3637__28_) );
DFFPOSX1 DFFPOSX1_844 ( .CLK(clock_i_bF_buf40), .D(_842_), .Q(_3637__27_) );
DFFPOSX1 DFFPOSX1_845 ( .CLK(clock_i_bF_buf74), .D(_843_), .Q(_3637__26_) );
DFFPOSX1 DFFPOSX1_846 ( .CLK(clock_i_bF_buf74), .D(_844_), .Q(_3637__25_) );
DFFPOSX1 DFFPOSX1_847 ( .CLK(clock_i_bF_buf49), .D(_845_), .Q(_3637__24_) );
DFFPOSX1 DFFPOSX1_848 ( .CLK(clock_i_bF_buf49), .D(_846_), .Q(_3637__23_) );
DFFPOSX1 DFFPOSX1_849 ( .CLK(clock_i_bF_buf40), .D(_847_), .Q(_3637__22_) );
DFFPOSX1 DFFPOSX1_850 ( .CLK(clock_i_bF_buf17), .D(_848_), .Q(_3637__21_) );
DFFPOSX1 DFFPOSX1_851 ( .CLK(clock_i_bF_buf13), .D(_849_), .Q(_3637__20_) );
DFFPOSX1 DFFPOSX1_852 ( .CLK(clock_i_bF_buf34), .D(_850_), .Q(_3637__19_) );
DFFPOSX1 DFFPOSX1_853 ( .CLK(clock_i_bF_buf34), .D(_851_), .Q(_3637__18_) );
DFFPOSX1 DFFPOSX1_854 ( .CLK(clock_i_bF_buf66), .D(_852_), .Q(_3637__17_) );
DFFPOSX1 DFFPOSX1_855 ( .CLK(clock_i_bF_buf81), .D(_853_), .Q(_3637__16_) );
DFFPOSX1 DFFPOSX1_856 ( .CLK(clock_i_bF_buf81), .D(_854_), .Q(_3637__15_) );
DFFPOSX1 DFFPOSX1_857 ( .CLK(clock_i_bF_buf66), .D(_855_), .Q(_3637__14_) );
DFFPOSX1 DFFPOSX1_858 ( .CLK(clock_i_bF_buf17), .D(_856_), .Q(_3637__13_) );
DFFPOSX1 DFFPOSX1_859 ( .CLK(clock_i_bF_buf26), .D(_857_), .Q(_3637__12_) );
DFFPOSX1 DFFPOSX1_860 ( .CLK(clock_i_bF_buf26), .D(_858_), .Q(_3637__11_) );
DFFPOSX1 DFFPOSX1_861 ( .CLK(clock_i_bF_buf26), .D(_859_), .Q(_3637__10_) );
DFFPOSX1 DFFPOSX1_862 ( .CLK(clock_i_bF_buf82), .D(_860_), .Q(_3637__9_) );
DFFPOSX1 DFFPOSX1_863 ( .CLK(clock_i_bF_buf82), .D(_861_), .Q(_3637__8_) );
DFFPOSX1 DFFPOSX1_864 ( .CLK(clock_i_bF_buf82), .D(_862_), .Q(_3637__7_) );
DFFPOSX1 DFFPOSX1_865 ( .CLK(clock_i_bF_buf82), .D(_863_), .Q(_3637__6_) );
DFFPOSX1 DFFPOSX1_866 ( .CLK(clock_i_bF_buf66), .D(_864_), .Q(_3637__5_) );
DFFPOSX1 DFFPOSX1_867 ( .CLK(clock_i_bF_buf33), .D(_865_), .Q(_3637__4_) );
DFFPOSX1 DFFPOSX1_868 ( .CLK(clock_i_bF_buf33), .D(_866_), .Q(_3637__3_) );
DFFPOSX1 DFFPOSX1_869 ( .CLK(clock_i_bF_buf5), .D(_867_), .Q(_3637__2_) );
DFFPOSX1 DFFPOSX1_870 ( .CLK(clock_i_bF_buf5), .D(_868_), .Q(_3637__1_) );
DFFPOSX1 DFFPOSX1_871 ( .CLK(clock_i_bF_buf5), .D(_869_), .Q(_3637__0_) );
DFFPOSX1 DFFPOSX1_872 ( .CLK(clock_i_bF_buf95), .D(_870_), .Q(_3638__63_) );
DFFPOSX1 DFFPOSX1_873 ( .CLK(clock_i_bF_buf24), .D(_871_), .Q(_3638__62_) );
DFFPOSX1 DFFPOSX1_874 ( .CLK(clock_i_bF_buf28), .D(_872_), .Q(_3638__61_) );
DFFPOSX1 DFFPOSX1_875 ( .CLK(clock_i_bF_buf90), .D(_873_), .Q(_3638__60_) );
DFFPOSX1 DFFPOSX1_876 ( .CLK(clock_i_bF_buf1), .D(_874_), .Q(_3638__59_) );
DFFPOSX1 DFFPOSX1_877 ( .CLK(clock_i_bF_buf71), .D(_875_), .Q(_3638__58_) );
DFFPOSX1 DFFPOSX1_878 ( .CLK(clock_i_bF_buf71), .D(_876_), .Q(_3638__57_) );
DFFPOSX1 DFFPOSX1_879 ( .CLK(clock_i_bF_buf71), .D(_877_), .Q(_3638__56_) );
DFFPOSX1 DFFPOSX1_880 ( .CLK(clock_i_bF_buf90), .D(_878_), .Q(_3638__55_) );
DFFPOSX1 DFFPOSX1_881 ( .CLK(clock_i_bF_buf28), .D(_879_), .Q(_3638__54_) );
DFFPOSX1 DFFPOSX1_882 ( .CLK(clock_i_bF_buf30), .D(_880_), .Q(_3638__53_) );
DFFPOSX1 DFFPOSX1_883 ( .CLK(clock_i_bF_buf91), .D(_881_), .Q(_3638__52_) );
DFFPOSX1 DFFPOSX1_884 ( .CLK(clock_i_bF_buf91), .D(_882_), .Q(_3638__51_) );
DFFPOSX1 DFFPOSX1_885 ( .CLK(clock_i_bF_buf52), .D(_883_), .Q(_3638__50_) );
DFFPOSX1 DFFPOSX1_886 ( .CLK(clock_i_bF_buf97), .D(_884_), .Q(_3638__49_) );
DFFPOSX1 DFFPOSX1_887 ( .CLK(clock_i_bF_buf37), .D(_885_), .Q(_3638__48_) );
DFFPOSX1 DFFPOSX1_888 ( .CLK(clock_i_bF_buf79), .D(_886_), .Q(_3638__47_) );
DFFPOSX1 DFFPOSX1_889 ( .CLK(clock_i_bF_buf43), .D(_887_), .Q(_3638__46_) );
DFFPOSX1 DFFPOSX1_890 ( .CLK(clock_i_bF_buf79), .D(_888_), .Q(_3638__45_) );
DFFPOSX1 DFFPOSX1_891 ( .CLK(clock_i_bF_buf67), .D(_889_), .Q(_3638__44_) );
DFFPOSX1 DFFPOSX1_892 ( .CLK(clock_i_bF_buf68), .D(_890_), .Q(_3638__43_) );
DFFPOSX1 DFFPOSX1_893 ( .CLK(clock_i_bF_buf25), .D(_891_), .Q(_3638__42_) );
DFFPOSX1 DFFPOSX1_894 ( .CLK(clock_i_bF_buf19), .D(_892_), .Q(_3638__41_) );
DFFPOSX1 DFFPOSX1_895 ( .CLK(clock_i_bF_buf68), .D(_893_), .Q(_3638__40_) );
DFFPOSX1 DFFPOSX1_896 ( .CLK(clock_i_bF_buf42), .D(_894_), .Q(_3638__39_) );
DFFPOSX1 DFFPOSX1_897 ( .CLK(clock_i_bF_buf67), .D(_895_), .Q(_3638__38_) );
DFFPOSX1 DFFPOSX1_898 ( .CLK(clock_i_bF_buf47), .D(_896_), .Q(_3638__37_) );
DFFPOSX1 DFFPOSX1_899 ( .CLK(clock_i_bF_buf53), .D(_897_), .Q(_3638__36_) );
DFFPOSX1 DFFPOSX1_900 ( .CLK(clock_i_bF_buf47), .D(_898_), .Q(_3638__35_) );
DFFPOSX1 DFFPOSX1_901 ( .CLK(clock_i_bF_buf67), .D(_899_), .Q(_3638__34_) );
DFFPOSX1 DFFPOSX1_902 ( .CLK(clock_i_bF_buf75), .D(_900_), .Q(_3638__33_) );
DFFPOSX1 DFFPOSX1_903 ( .CLK(clock_i_bF_buf81), .D(_901_), .Q(_3638__32_) );
DFFPOSX1 DFFPOSX1_904 ( .CLK(clock_i_bF_buf34), .D(_902_), .Q(_3638__31_) );
DFFPOSX1 DFFPOSX1_905 ( .CLK(clock_i_bF_buf53), .D(_903_), .Q(_3638__30_) );
DFFPOSX1 DFFPOSX1_906 ( .CLK(clock_i_bF_buf13), .D(_904_), .Q(_3638__29_) );
DFFPOSX1 DFFPOSX1_907 ( .CLK(clock_i_bF_buf49), .D(_905_), .Q(_3638__28_) );
DFFPOSX1 DFFPOSX1_908 ( .CLK(clock_i_bF_buf40), .D(_906_), .Q(_3638__27_) );
DFFPOSX1 DFFPOSX1_909 ( .CLK(clock_i_bF_buf25), .D(_907_), .Q(_3638__26_) );
DFFPOSX1 DFFPOSX1_910 ( .CLK(clock_i_bF_buf74), .D(_908_), .Q(_3638__25_) );
DFFPOSX1 DFFPOSX1_911 ( .CLK(clock_i_bF_buf40), .D(_909_), .Q(_3638__24_) );
DFFPOSX1 DFFPOSX1_912 ( .CLK(clock_i_bF_buf49), .D(_910_), .Q(_3638__23_) );
DFFPOSX1 DFFPOSX1_913 ( .CLK(clock_i_bF_buf74), .D(_911_), .Q(_3638__22_) );
DFFPOSX1 DFFPOSX1_914 ( .CLK(clock_i_bF_buf17), .D(_912_), .Q(_3638__21_) );
DFFPOSX1 DFFPOSX1_915 ( .CLK(clock_i_bF_buf53), .D(_913_), .Q(_3638__20_) );
DFFPOSX1 DFFPOSX1_916 ( .CLK(clock_i_bF_buf34), .D(_914_), .Q(_3638__19_) );
DFFPOSX1 DFFPOSX1_917 ( .CLK(clock_i_bF_buf25), .D(_915_), .Q(_3638__18_) );
DFFPOSX1 DFFPOSX1_918 ( .CLK(clock_i_bF_buf34), .D(_916_), .Q(_3638__17_) );
DFFPOSX1 DFFPOSX1_919 ( .CLK(clock_i_bF_buf81), .D(_917_), .Q(_3638__16_) );
DFFPOSX1 DFFPOSX1_920 ( .CLK(clock_i_bF_buf81), .D(_918_), .Q(_3638__15_) );
DFFPOSX1 DFFPOSX1_921 ( .CLK(clock_i_bF_buf66), .D(_919_), .Q(_3638__14_) );
DFFPOSX1 DFFPOSX1_922 ( .CLK(clock_i_bF_buf17), .D(_920_), .Q(_3638__13_) );
DFFPOSX1 DFFPOSX1_923 ( .CLK(clock_i_bF_buf64), .D(_921_), .Q(_3638__12_) );
DFFPOSX1 DFFPOSX1_924 ( .CLK(clock_i_bF_buf33), .D(_922_), .Q(_3638__11_) );
DFFPOSX1 DFFPOSX1_925 ( .CLK(clock_i_bF_buf66), .D(_923_), .Q(_3638__10_) );
DFFPOSX1 DFFPOSX1_926 ( .CLK(clock_i_bF_buf26), .D(_924_), .Q(_3638__9_) );
DFFPOSX1 DFFPOSX1_927 ( .CLK(clock_i_bF_buf33), .D(_925_), .Q(_3638__8_) );
DFFPOSX1 DFFPOSX1_928 ( .CLK(clock_i_bF_buf65), .D(_926_), .Q(_3638__7_) );
DFFPOSX1 DFFPOSX1_929 ( .CLK(clock_i_bF_buf66), .D(_927_), .Q(_3638__6_) );
DFFPOSX1 DFFPOSX1_930 ( .CLK(clock_i_bF_buf74), .D(_928_), .Q(_3638__5_) );
DFFPOSX1 DFFPOSX1_931 ( .CLK(clock_i_bF_buf62), .D(_929_), .Q(_3638__4_) );
DFFPOSX1 DFFPOSX1_932 ( .CLK(clock_i_bF_buf5), .D(_930_), .Q(_3638__3_) );
DFFPOSX1 DFFPOSX1_933 ( .CLK(clock_i_bF_buf33), .D(_931_), .Q(_3638__2_) );
DFFPOSX1 DFFPOSX1_934 ( .CLK(clock_i_bF_buf72), .D(_932_), .Q(_3638__1_) );
DFFPOSX1 DFFPOSX1_935 ( .CLK(clock_i_bF_buf5), .D(_933_), .Q(_3638__0_) );
DFFPOSX1 DFFPOSX1_936 ( .CLK(clock_i_bF_buf45), .D(_934_), .Q(_3639__63_) );
DFFPOSX1 DFFPOSX1_937 ( .CLK(clock_i_bF_buf29), .D(_935_), .Q(_3639__62_) );
DFFPOSX1 DFFPOSX1_938 ( .CLK(clock_i_bF_buf11), .D(_936_), .Q(_3639__61_) );
DFFPOSX1 DFFPOSX1_939 ( .CLK(clock_i_bF_buf59), .D(_937_), .Q(_3639__60_) );
DFFPOSX1 DFFPOSX1_940 ( .CLK(clock_i_bF_buf18), .D(_938_), .Q(_3639__59_) );
DFFPOSX1 DFFPOSX1_941 ( .CLK(clock_i_bF_buf71), .D(_939_), .Q(_3639__58_) );
DFFPOSX1 DFFPOSX1_942 ( .CLK(clock_i_bF_buf4), .D(_940_), .Q(_3639__57_) );
DFFPOSX1 DFFPOSX1_943 ( .CLK(clock_i_bF_buf30), .D(_941_), .Q(_3639__56_) );
DFFPOSX1 DFFPOSX1_944 ( .CLK(clock_i_bF_buf71), .D(_942_), .Q(_3639__55_) );
DFFPOSX1 DFFPOSX1_945 ( .CLK(clock_i_bF_buf11), .D(_943_), .Q(_3639__54_) );
DFFPOSX1 DFFPOSX1_946 ( .CLK(clock_i_bF_buf30), .D(_944_), .Q(_3639__53_) );
DFFPOSX1 DFFPOSX1_947 ( .CLK(clock_i_bF_buf32), .D(_945_), .Q(_3639__52_) );
DFFPOSX1 DFFPOSX1_948 ( .CLK(clock_i_bF_buf73), .D(_946_), .Q(_3639__51_) );
DFFPOSX1 DFFPOSX1_949 ( .CLK(clock_i_bF_buf97), .D(_947_), .Q(_3639__50_) );
DFFPOSX1 DFFPOSX1_950 ( .CLK(clock_i_bF_buf32), .D(_948_), .Q(_3639__49_) );
DFFPOSX1 DFFPOSX1_951 ( .CLK(clock_i_bF_buf101), .D(_949_), .Q(_3639__48_) );
DFFPOSX1 DFFPOSX1_952 ( .CLK(clock_i_bF_buf79), .D(_950_), .Q(_3639__47_) );
DFFPOSX1 DFFPOSX1_953 ( .CLK(clock_i_bF_buf79), .D(_951_), .Q(_3639__46_) );
DFFPOSX1 DFFPOSX1_954 ( .CLK(clock_i_bF_buf86), .D(_952_), .Q(_3639__45_) );
DFFPOSX1 DFFPOSX1_955 ( .CLK(clock_i_bF_buf42), .D(_953_), .Q(_3639__44_) );
DFFPOSX1 DFFPOSX1_956 ( .CLK(clock_i_bF_buf19), .D(_954_), .Q(_3639__43_) );
DFFPOSX1 DFFPOSX1_957 ( .CLK(clock_i_bF_buf68), .D(_955_), .Q(_3639__42_) );
DFFPOSX1 DFFPOSX1_958 ( .CLK(clock_i_bF_buf68), .D(_956_), .Q(_3639__41_) );
DFFPOSX1 DFFPOSX1_959 ( .CLK(clock_i_bF_buf68), .D(_957_), .Q(_3639__40_) );
DFFPOSX1 DFFPOSX1_960 ( .CLK(clock_i_bF_buf67), .D(_958_), .Q(_3639__39_) );
DFFPOSX1 DFFPOSX1_961 ( .CLK(clock_i_bF_buf47), .D(_959_), .Q(_3639__38_) );
DFFPOSX1 DFFPOSX1_962 ( .CLK(clock_i_bF_buf47), .D(_960_), .Q(_3639__37_) );
DFFPOSX1 DFFPOSX1_963 ( .CLK(clock_i_bF_buf53), .D(_961_), .Q(_3639__36_) );
DFFPOSX1 DFFPOSX1_964 ( .CLK(clock_i_bF_buf75), .D(_962_), .Q(_3639__35_) );
DFFPOSX1 DFFPOSX1_965 ( .CLK(clock_i_bF_buf53), .D(_963_), .Q(_3639__34_) );
DFFPOSX1 DFFPOSX1_966 ( .CLK(clock_i_bF_buf75), .D(_964_), .Q(_3639__33_) );
DFFPOSX1 DFFPOSX1_967 ( .CLK(clock_i_bF_buf81), .D(_965_), .Q(_3639__32_) );
DFFPOSX1 DFFPOSX1_968 ( .CLK(clock_i_bF_buf13), .D(_966_), .Q(_3639__31_) );
DFFPOSX1 DFFPOSX1_969 ( .CLK(clock_i_bF_buf34), .D(_967_), .Q(_3639__30_) );
DFFPOSX1 DFFPOSX1_970 ( .CLK(clock_i_bF_buf17), .D(_968_), .Q(_3639__29_) );
DFFPOSX1 DFFPOSX1_971 ( .CLK(clock_i_bF_buf21), .D(_969_), .Q(_3639__28_) );
DFFPOSX1 DFFPOSX1_972 ( .CLK(clock_i_bF_buf17), .D(_970_), .Q(_3639__27_) );
DFFPOSX1 DFFPOSX1_973 ( .CLK(clock_i_bF_buf17), .D(_971_), .Q(_3639__26_) );
DFFPOSX1 DFFPOSX1_974 ( .CLK(clock_i_bF_buf74), .D(_972_), .Q(_3639__25_) );
DFFPOSX1 DFFPOSX1_975 ( .CLK(clock_i_bF_buf68), .D(_973_), .Q(_3639__24_) );
DFFPOSX1 DFFPOSX1_976 ( .CLK(clock_i_bF_buf26), .D(_974_), .Q(_3639__23_) );
DFFPOSX1 DFFPOSX1_977 ( .CLK(clock_i_bF_buf17), .D(_975_), .Q(_3639__22_) );
DFFPOSX1 DFFPOSX1_978 ( .CLK(clock_i_bF_buf17), .D(_976_), .Q(_3639__21_) );
DFFPOSX1 DFFPOSX1_979 ( .CLK(clock_i_bF_buf66), .D(_977_), .Q(_3639__20_) );
DFFPOSX1 DFFPOSX1_980 ( .CLK(clock_i_bF_buf34), .D(_978_), .Q(_3639__19_) );
DFFPOSX1 DFFPOSX1_981 ( .CLK(clock_i_bF_buf72), .D(_979_), .Q(_3639__18_) );
DFFPOSX1 DFFPOSX1_982 ( .CLK(clock_i_bF_buf34), .D(_980_), .Q(_3639__17_) );
DFFPOSX1 DFFPOSX1_983 ( .CLK(clock_i_bF_buf72), .D(_981_), .Q(_3639__16_) );
DFFPOSX1 DFFPOSX1_984 ( .CLK(clock_i_bF_buf72), .D(_982_), .Q(_3639__15_) );
DFFPOSX1 DFFPOSX1_985 ( .CLK(clock_i_bF_buf16), .D(_983_), .Q(_3639__14_) );
DFFPOSX1 DFFPOSX1_986 ( .CLK(clock_i_bF_buf21), .D(_984_), .Q(_3639__13_) );
DFFPOSX1 DFFPOSX1_987 ( .CLK(clock_i_bF_buf74), .D(_985_), .Q(_3639__12_) );
DFFPOSX1 DFFPOSX1_988 ( .CLK(clock_i_bF_buf17), .D(_986_), .Q(_3639__11_) );
DFFPOSX1 DFFPOSX1_989 ( .CLK(clock_i_bF_buf74), .D(_987_), .Q(_3639__10_) );
DFFPOSX1 DFFPOSX1_990 ( .CLK(clock_i_bF_buf82), .D(_988_), .Q(_3639__9_) );
DFFPOSX1 DFFPOSX1_991 ( .CLK(clock_i_bF_buf82), .D(_989_), .Q(_3639__8_) );
DFFPOSX1 DFFPOSX1_992 ( .CLK(clock_i_bF_buf82), .D(_990_), .Q(_3639__7_) );
DFFPOSX1 DFFPOSX1_993 ( .CLK(clock_i_bF_buf82), .D(_991_), .Q(_3639__6_) );
DFFPOSX1 DFFPOSX1_994 ( .CLK(clock_i_bF_buf66), .D(_992_), .Q(_3639__5_) );
DFFPOSX1 DFFPOSX1_995 ( .CLK(clock_i_bF_buf33), .D(_993_), .Q(_3639__4_) );
DFFPOSX1 DFFPOSX1_996 ( .CLK(clock_i_bF_buf62), .D(_994_), .Q(_3639__3_) );
DFFPOSX1 DFFPOSX1_997 ( .CLK(clock_i_bF_buf66), .D(_995_), .Q(_3639__2_) );
DFFPOSX1 DFFPOSX1_998 ( .CLK(clock_i_bF_buf72), .D(_996_), .Q(_3639__1_) );
DFFPOSX1 DFFPOSX1_999 ( .CLK(clock_i_bF_buf5), .D(_997_), .Q(_3639__0_) );
DFFPOSX1 DFFPOSX1_1000 ( .CLK(clock_i_bF_buf97), .D(_998_), .Q(_3648_) );
DFFPOSX1 DFFPOSX1_1001 ( .CLK(clock_i_bF_buf97), .D(_999_), .Q(_3649_) );
DFFPOSX1 DFFPOSX1_1002 ( .CLK(clock_i_bF_buf67), .D(_1000_), .Q(_3650_) );
DFFPOSX1 DFFPOSX1_1003 ( .CLK(clock_i_bF_buf25), .D(_1001_), .Q(_3651_) );
DFFPOSX1 DFFPOSX1_1004 ( .CLK(clock_i_bF_buf94), .D(_1002_), .Q(_3656__31_) );
DFFPOSX1 DFFPOSX1_1005 ( .CLK(clock_i_bF_buf37), .D(_1003_), .Q(_3656__30_) );
DFFPOSX1 DFFPOSX1_1006 ( .CLK(clock_i_bF_buf3), .D(_1004_), .Q(_3656__29_) );
DFFPOSX1 DFFPOSX1_1007 ( .CLK(clock_i_bF_buf99), .D(_1005_), .Q(_3656__28_) );
DFFPOSX1 DFFPOSX1_1008 ( .CLK(clock_i_bF_buf98), .D(_1006_), .Q(_3656__27_) );
DFFPOSX1 DFFPOSX1_1009 ( .CLK(clock_i_bF_buf44), .D(_1007_), .Q(_3656__26_) );
DFFPOSX1 DFFPOSX1_1010 ( .CLK(clock_i_bF_buf61), .D(_1008_), .Q(_3656__25_) );
DFFPOSX1 DFFPOSX1_1011 ( .CLK(clock_i_bF_buf9), .D(_1009_), .Q(_3656__24_) );
DFFPOSX1 DFFPOSX1_1012 ( .CLK(clock_i_bF_buf94), .D(_1010_), .Q(_3656__23_) );
DFFPOSX1 DFFPOSX1_1013 ( .CLK(clock_i_bF_buf45), .D(_1011_), .Q(_3656__22_) );
DFFPOSX1 DFFPOSX1_1014 ( .CLK(clock_i_bF_buf94), .D(_1012_), .Q(_3656__21_) );
DFFPOSX1 DFFPOSX1_1015 ( .CLK(clock_i_bF_buf38), .D(_1013_), .Q(_3656__20_) );
DFFPOSX1 DFFPOSX1_1016 ( .CLK(clock_i_bF_buf29), .D(_1014_), .Q(_3656__19_) );
DFFPOSX1 DFFPOSX1_1017 ( .CLK(clock_i_bF_buf99), .D(_1015_), .Q(_3656__18_) );
DFFPOSX1 DFFPOSX1_1018 ( .CLK(clock_i_bF_buf94), .D(_1016_), .Q(_3656__17_) );
DFFPOSX1 DFFPOSX1_1019 ( .CLK(clock_i_bF_buf45), .D(_1017_), .Q(_3656__16_) );
DFFPOSX1 DFFPOSX1_1020 ( .CLK(clock_i_bF_buf91), .D(_1018_), .Q(_3656__15_) );
DFFPOSX1 DFFPOSX1_1021 ( .CLK(clock_i_bF_buf7), .D(_1019_), .Q(_3656__14_) );
DFFPOSX1 DFFPOSX1_1022 ( .CLK(clock_i_bF_buf29), .D(_1020_), .Q(_3656__13_) );
DFFPOSX1 DFFPOSX1_1023 ( .CLK(clock_i_bF_buf57), .D(_1021_), .Q(_3656__12_) );
DFFPOSX1 DFFPOSX1_1024 ( .CLK(clock_i_bF_buf60), .D(_1022_), .Q(_3656__11_) );
DFFPOSX1 DFFPOSX1_1025 ( .CLK(clock_i_bF_buf38), .D(_1023_), .Q(_3656__10_) );
DFFPOSX1 DFFPOSX1_1026 ( .CLK(clock_i_bF_buf59), .D(_1024_), .Q(_3656__9_) );
DFFPOSX1 DFFPOSX1_1027 ( .CLK(clock_i_bF_buf70), .D(_1025_), .Q(_3656__8_) );
DFFPOSX1 DFFPOSX1_1028 ( .CLK(clock_i_bF_buf51), .D(_1026_), .Q(_3656__7_) );
DFFPOSX1 DFFPOSX1_1029 ( .CLK(clock_i_bF_buf50), .D(_1027_), .Q(_3656__6_) );
DFFPOSX1 DFFPOSX1_1030 ( .CLK(clock_i_bF_buf3), .D(_1028_), .Q(_3656__5_) );
DFFPOSX1 DFFPOSX1_1031 ( .CLK(clock_i_bF_buf86), .D(_1029_), .Q(_3656__4_) );
DFFPOSX1 DFFPOSX1_1032 ( .CLK(clock_i_bF_buf1), .D(_1030_), .Q(_3656__3_) );
BUFX2 BUFX2_1 ( .A(_3636__63_), .Y(addr1_o[63]) );
BUFX2 BUFX2_2 ( .A(_3636__62_), .Y(addr1_o[62]) );
BUFX2 BUFX2_3 ( .A(_3636__53_), .Y(addr1_o[53]) );
BUFX2 BUFX2_4 ( .A(_3636__52_), .Y(addr1_o[52]) );
BUFX2 BUFX2_5 ( .A(_3636__51_), .Y(addr1_o[51]) );
BUFX2 BUFX2_6 ( .A(_3636__50_), .Y(addr1_o[50]) );
BUFX2 BUFX2_7 ( .A(_3636__49_), .Y(addr1_o[49]) );
BUFX2 BUFX2_8 ( .A(_3636__48_), .Y(addr1_o[48]) );
BUFX2 BUFX2_9 ( .A(_3636__47_), .Y(addr1_o[47]) );
BUFX2 BUFX2_10 ( .A(_3636__46_), .Y(addr1_o[46]) );
BUFX2 BUFX2_11 ( .A(_3636__45_), .Y(addr1_o[45]) );
BUFX2 BUFX2_12 ( .A(_3636__44_), .Y(addr1_o[44]) );
BUFX2 BUFX2_13 ( .A(_3636__61_), .Y(addr1_o[61]) );
BUFX2 BUFX2_14 ( .A(_3636__43_), .Y(addr1_o[43]) );
BUFX2 BUFX2_15 ( .A(_3636__42_), .Y(addr1_o[42]) );
BUFX2 BUFX2_16 ( .A(_3636__41_), .Y(addr1_o[41]) );
BUFX2 BUFX2_17 ( .A(_3636__40_), .Y(addr1_o[40]) );
BUFX2 BUFX2_18 ( .A(_3636__39_), .Y(addr1_o[39]) );
BUFX2 BUFX2_19 ( .A(_3636__38_), .Y(addr1_o[38]) );
BUFX2 BUFX2_20 ( .A(_3636__37_), .Y(addr1_o[37]) );
BUFX2 BUFX2_21 ( .A(_3636__36_), .Y(addr1_o[36]) );
BUFX2 BUFX2_22 ( .A(_3636__35_), .Y(addr1_o[35]) );
BUFX2 BUFX2_23 ( .A(_3636__34_), .Y(addr1_o[34]) );
BUFX2 BUFX2_24 ( .A(_3636__60_), .Y(addr1_o[60]) );
BUFX2 BUFX2_25 ( .A(_3636__33_), .Y(addr1_o[33]) );
BUFX2 BUFX2_26 ( .A(_3636__32_), .Y(addr1_o[32]) );
BUFX2 BUFX2_27 ( .A(_3636__31_), .Y(addr1_o[31]) );
BUFX2 BUFX2_28 ( .A(_3636__30_), .Y(addr1_o[30]) );
BUFX2 BUFX2_29 ( .A(_3636__29_), .Y(addr1_o[29]) );
BUFX2 BUFX2_30 ( .A(_3636__28_), .Y(addr1_o[28]) );
BUFX2 BUFX2_31 ( .A(_3636__27_), .Y(addr1_o[27]) );
BUFX2 BUFX2_32 ( .A(_3636__26_), .Y(addr1_o[26]) );
BUFX2 BUFX2_33 ( .A(_3636__25_), .Y(addr1_o[25]) );
BUFX2 BUFX2_34 ( .A(_3636__24_), .Y(addr1_o[24]) );
BUFX2 BUFX2_35 ( .A(_3636__59_), .Y(addr1_o[59]) );
BUFX2 BUFX2_36 ( .A(_3636__23_), .Y(addr1_o[23]) );
BUFX2 BUFX2_37 ( .A(_3636__22_), .Y(addr1_o[22]) );
BUFX2 BUFX2_38 ( .A(_3636__21_), .Y(addr1_o[21]) );
BUFX2 BUFX2_39 ( .A(_3636__20_), .Y(addr1_o[20]) );
BUFX2 BUFX2_40 ( .A(_3636__19_), .Y(addr1_o[19]) );
BUFX2 BUFX2_41 ( .A(_3636__18_), .Y(addr1_o[18]) );
BUFX2 BUFX2_42 ( .A(_3636__17_), .Y(addr1_o[17]) );
BUFX2 BUFX2_43 ( .A(_3636__16_), .Y(addr1_o[16]) );
BUFX2 BUFX2_44 ( .A(_3636__15_), .Y(addr1_o[15]) );
BUFX2 BUFX2_45 ( .A(_3636__14_), .Y(addr1_o[14]) );
BUFX2 BUFX2_46 ( .A(_3636__58_), .Y(addr1_o[58]) );
BUFX2 BUFX2_47 ( .A(_3636__13_), .Y(addr1_o[13]) );
BUFX2 BUFX2_48 ( .A(_3636__12_), .Y(addr1_o[12]) );
BUFX2 BUFX2_49 ( .A(_3636__11_), .Y(addr1_o[11]) );
BUFX2 BUFX2_50 ( .A(_3636__10_), .Y(addr1_o[10]) );
BUFX2 BUFX2_51 ( .A(_3636__9_), .Y(addr1_o[9]) );
BUFX2 BUFX2_52 ( .A(_3636__8_), .Y(addr1_o[8]) );
BUFX2 BUFX2_53 ( .A(_3636__7_), .Y(addr1_o[7]) );
BUFX2 BUFX2_54 ( .A(_3636__6_), .Y(addr1_o[6]) );
BUFX2 BUFX2_55 ( .A(_3636__5_), .Y(addr1_o[5]) );
BUFX2 BUFX2_56 ( .A(_3636__4_), .Y(addr1_o[4]) );
BUFX2 BUFX2_57 ( .A(_3636__57_), .Y(addr1_o[57]) );
BUFX2 BUFX2_58 ( .A(_3636__3_), .Y(addr1_o[3]) );
BUFX2 BUFX2_59 ( .A(_3636__2_), .Y(addr1_o[2]) );
BUFX2 BUFX2_60 ( .A(_3636__1_), .Y(addr1_o[1]) );
BUFX2 BUFX2_61 ( .A(_3636__0_), .Y(addr1_o[0]) );
BUFX2 BUFX2_62 ( .A(_3636__56_), .Y(addr1_o[56]) );
BUFX2 BUFX2_63 ( .A(_3636__55_), .Y(addr1_o[55]) );
BUFX2 BUFX2_64 ( .A(_3636__54_), .Y(addr1_o[54]) );
BUFX2 BUFX2_65 ( .A(_3637__63_), .Y(addr2_o[63]) );
BUFX2 BUFX2_66 ( .A(_3637__62_), .Y(addr2_o[62]) );
BUFX2 BUFX2_67 ( .A(_3637__53_), .Y(addr2_o[53]) );
BUFX2 BUFX2_68 ( .A(_3637__52_), .Y(addr2_o[52]) );
BUFX2 BUFX2_69 ( .A(_3637__51_), .Y(addr2_o[51]) );
BUFX2 BUFX2_70 ( .A(_3637__50_), .Y(addr2_o[50]) );
BUFX2 BUFX2_71 ( .A(_3637__49_), .Y(addr2_o[49]) );
BUFX2 BUFX2_72 ( .A(_3637__48_), .Y(addr2_o[48]) );
BUFX2 BUFX2_73 ( .A(_3637__47_), .Y(addr2_o[47]) );
BUFX2 BUFX2_74 ( .A(_3637__46_), .Y(addr2_o[46]) );
BUFX2 BUFX2_75 ( .A(_3637__45_), .Y(addr2_o[45]) );
BUFX2 BUFX2_76 ( .A(_3637__44_), .Y(addr2_o[44]) );
BUFX2 BUFX2_77 ( .A(_3637__61_), .Y(addr2_o[61]) );
BUFX2 BUFX2_78 ( .A(_3637__43_), .Y(addr2_o[43]) );
BUFX2 BUFX2_79 ( .A(_3637__42_), .Y(addr2_o[42]) );
BUFX2 BUFX2_80 ( .A(_3637__41_), .Y(addr2_o[41]) );
BUFX2 BUFX2_81 ( .A(_3637__40_), .Y(addr2_o[40]) );
BUFX2 BUFX2_82 ( .A(_3637__39_), .Y(addr2_o[39]) );
BUFX2 BUFX2_83 ( .A(_3637__38_), .Y(addr2_o[38]) );
BUFX2 BUFX2_84 ( .A(_3637__37_), .Y(addr2_o[37]) );
BUFX2 BUFX2_85 ( .A(_3637__36_), .Y(addr2_o[36]) );
BUFX2 BUFX2_86 ( .A(_3637__35_), .Y(addr2_o[35]) );
BUFX2 BUFX2_87 ( .A(_3637__34_), .Y(addr2_o[34]) );
BUFX2 BUFX2_88 ( .A(_3637__60_), .Y(addr2_o[60]) );
BUFX2 BUFX2_89 ( .A(_3637__33_), .Y(addr2_o[33]) );
BUFX2 BUFX2_90 ( .A(_3637__32_), .Y(addr2_o[32]) );
BUFX2 BUFX2_91 ( .A(_3637__31_), .Y(addr2_o[31]) );
BUFX2 BUFX2_92 ( .A(_3637__30_), .Y(addr2_o[30]) );
BUFX2 BUFX2_93 ( .A(_3637__29_), .Y(addr2_o[29]) );
BUFX2 BUFX2_94 ( .A(_3637__28_), .Y(addr2_o[28]) );
BUFX2 BUFX2_95 ( .A(_3637__27_), .Y(addr2_o[27]) );
BUFX2 BUFX2_96 ( .A(_3637__26_), .Y(addr2_o[26]) );
BUFX2 BUFX2_97 ( .A(_3637__25_), .Y(addr2_o[25]) );
BUFX2 BUFX2_98 ( .A(_3637__24_), .Y(addr2_o[24]) );
BUFX2 BUFX2_99 ( .A(_3637__59_), .Y(addr2_o[59]) );
BUFX2 BUFX2_100 ( .A(_3637__23_), .Y(addr2_o[23]) );
BUFX2 BUFX2_101 ( .A(_3637__22_), .Y(addr2_o[22]) );
BUFX2 BUFX2_102 ( .A(_3637__21_), .Y(addr2_o[21]) );
BUFX2 BUFX2_103 ( .A(_3637__20_), .Y(addr2_o[20]) );
BUFX2 BUFX2_104 ( .A(_3637__19_), .Y(addr2_o[19]) );
BUFX2 BUFX2_105 ( .A(_3637__18_), .Y(addr2_o[18]) );
BUFX2 BUFX2_106 ( .A(_3637__17_), .Y(addr2_o[17]) );
BUFX2 BUFX2_107 ( .A(_3637__16_), .Y(addr2_o[16]) );
BUFX2 BUFX2_108 ( .A(_3637__15_), .Y(addr2_o[15]) );
BUFX2 BUFX2_109 ( .A(_3637__14_), .Y(addr2_o[14]) );
BUFX2 BUFX2_110 ( .A(_3637__58_), .Y(addr2_o[58]) );
BUFX2 BUFX2_111 ( .A(_3637__13_), .Y(addr2_o[13]) );
BUFX2 BUFX2_112 ( .A(_3637__12_), .Y(addr2_o[12]) );
BUFX2 BUFX2_113 ( .A(_3637__11_), .Y(addr2_o[11]) );
BUFX2 BUFX2_114 ( .A(_3637__10_), .Y(addr2_o[10]) );
BUFX2 BUFX2_115 ( .A(_3637__9_), .Y(addr2_o[9]) );
BUFX2 BUFX2_116 ( .A(_3637__8_), .Y(addr2_o[8]) );
BUFX2 BUFX2_117 ( .A(_3637__7_), .Y(addr2_o[7]) );
BUFX2 BUFX2_118 ( .A(_3637__6_), .Y(addr2_o[6]) );
BUFX2 BUFX2_119 ( .A(_3637__5_), .Y(addr2_o[5]) );
BUFX2 BUFX2_120 ( .A(_3637__4_), .Y(addr2_o[4]) );
BUFX2 BUFX2_121 ( .A(_3637__57_), .Y(addr2_o[57]) );
BUFX2 BUFX2_122 ( .A(_3637__3_), .Y(addr2_o[3]) );
BUFX2 BUFX2_123 ( .A(_3637__2_), .Y(addr2_o[2]) );
BUFX2 BUFX2_124 ( .A(_3637__1_), .Y(addr2_o[1]) );
BUFX2 BUFX2_125 ( .A(_3637__0_), .Y(addr2_o[0]) );
BUFX2 BUFX2_126 ( .A(_3637__56_), .Y(addr2_o[56]) );
BUFX2 BUFX2_127 ( .A(_3637__55_), .Y(addr2_o[55]) );
BUFX2 BUFX2_128 ( .A(_3637__54_), .Y(addr2_o[54]) );
BUFX2 BUFX2_129 ( .A(_3638__63_), .Y(addr3_o[63]) );
BUFX2 BUFX2_130 ( .A(_3638__62_), .Y(addr3_o[62]) );
BUFX2 BUFX2_131 ( .A(_3638__53_), .Y(addr3_o[53]) );
BUFX2 BUFX2_132 ( .A(_3638__52_), .Y(addr3_o[52]) );
BUFX2 BUFX2_133 ( .A(_3638__51_), .Y(addr3_o[51]) );
BUFX2 BUFX2_134 ( .A(_3638__50_), .Y(addr3_o[50]) );
BUFX2 BUFX2_135 ( .A(_3638__49_), .Y(addr3_o[49]) );
BUFX2 BUFX2_136 ( .A(_3638__48_), .Y(addr3_o[48]) );
BUFX2 BUFX2_137 ( .A(_3638__47_), .Y(addr3_o[47]) );
BUFX2 BUFX2_138 ( .A(_3638__46_), .Y(addr3_o[46]) );
BUFX2 BUFX2_139 ( .A(_3638__45_), .Y(addr3_o[45]) );
BUFX2 BUFX2_140 ( .A(_3638__44_), .Y(addr3_o[44]) );
BUFX2 BUFX2_141 ( .A(_3638__61_), .Y(addr3_o[61]) );
BUFX2 BUFX2_142 ( .A(_3638__43_), .Y(addr3_o[43]) );
BUFX2 BUFX2_143 ( .A(_3638__42_), .Y(addr3_o[42]) );
BUFX2 BUFX2_144 ( .A(_3638__41_), .Y(addr3_o[41]) );
BUFX2 BUFX2_145 ( .A(_3638__40_), .Y(addr3_o[40]) );
BUFX2 BUFX2_146 ( .A(_3638__39_), .Y(addr3_o[39]) );
BUFX2 BUFX2_147 ( .A(_3638__38_), .Y(addr3_o[38]) );
BUFX2 BUFX2_148 ( .A(_3638__37_), .Y(addr3_o[37]) );
BUFX2 BUFX2_149 ( .A(_3638__36_), .Y(addr3_o[36]) );
BUFX2 BUFX2_150 ( .A(_3638__35_), .Y(addr3_o[35]) );
BUFX2 BUFX2_151 ( .A(_3638__34_), .Y(addr3_o[34]) );
BUFX2 BUFX2_152 ( .A(_3638__60_), .Y(addr3_o[60]) );
BUFX2 BUFX2_153 ( .A(_3638__33_), .Y(addr3_o[33]) );
BUFX2 BUFX2_154 ( .A(_3638__32_), .Y(addr3_o[32]) );
BUFX2 BUFX2_155 ( .A(_3638__31_), .Y(addr3_o[31]) );
BUFX2 BUFX2_156 ( .A(_3638__30_), .Y(addr3_o[30]) );
BUFX2 BUFX2_157 ( .A(_3638__29_), .Y(addr3_o[29]) );
BUFX2 BUFX2_158 ( .A(_3638__28_), .Y(addr3_o[28]) );
BUFX2 BUFX2_159 ( .A(_3638__27_), .Y(addr3_o[27]) );
BUFX2 BUFX2_160 ( .A(_3638__26_), .Y(addr3_o[26]) );
BUFX2 BUFX2_161 ( .A(_3638__25_), .Y(addr3_o[25]) );
BUFX2 BUFX2_162 ( .A(_3638__24_), .Y(addr3_o[24]) );
BUFX2 BUFX2_163 ( .A(_3638__59_), .Y(addr3_o[59]) );
BUFX2 BUFX2_164 ( .A(_3638__23_), .Y(addr3_o[23]) );
BUFX2 BUFX2_165 ( .A(_3638__22_), .Y(addr3_o[22]) );
BUFX2 BUFX2_166 ( .A(_3638__21_), .Y(addr3_o[21]) );
BUFX2 BUFX2_167 ( .A(_3638__20_), .Y(addr3_o[20]) );
BUFX2 BUFX2_168 ( .A(_3638__19_), .Y(addr3_o[19]) );
BUFX2 BUFX2_169 ( .A(_3638__18_), .Y(addr3_o[18]) );
BUFX2 BUFX2_170 ( .A(_3638__17_), .Y(addr3_o[17]) );
BUFX2 BUFX2_171 ( .A(_3638__16_), .Y(addr3_o[16]) );
BUFX2 BUFX2_172 ( .A(_3638__15_), .Y(addr3_o[15]) );
BUFX2 BUFX2_173 ( .A(_3638__14_), .Y(addr3_o[14]) );
BUFX2 BUFX2_174 ( .A(_3638__58_), .Y(addr3_o[58]) );
BUFX2 BUFX2_175 ( .A(_3638__13_), .Y(addr3_o[13]) );
BUFX2 BUFX2_176 ( .A(_3638__12_), .Y(addr3_o[12]) );
BUFX2 BUFX2_177 ( .A(_3638__11_), .Y(addr3_o[11]) );
BUFX2 BUFX2_178 ( .A(_3638__10_), .Y(addr3_o[10]) );
BUFX2 BUFX2_179 ( .A(_3638__9_), .Y(addr3_o[9]) );
BUFX2 BUFX2_180 ( .A(_3638__8_), .Y(addr3_o[8]) );
BUFX2 BUFX2_181 ( .A(_3638__7_), .Y(addr3_o[7]) );
BUFX2 BUFX2_182 ( .A(_3638__6_), .Y(addr3_o[6]) );
BUFX2 BUFX2_183 ( .A(_3638__5_), .Y(addr3_o[5]) );
BUFX2 BUFX2_184 ( .A(_3638__4_), .Y(addr3_o[4]) );
BUFX2 BUFX2_185 ( .A(_3638__57_), .Y(addr3_o[57]) );
BUFX2 BUFX2_186 ( .A(_3638__3_), .Y(addr3_o[3]) );
BUFX2 BUFX2_187 ( .A(_3638__2_), .Y(addr3_o[2]) );
BUFX2 BUFX2_188 ( .A(_3638__1_), .Y(addr3_o[1]) );
BUFX2 BUFX2_189 ( .A(_3638__0_), .Y(addr3_o[0]) );
BUFX2 BUFX2_190 ( .A(_3638__56_), .Y(addr3_o[56]) );
BUFX2 BUFX2_191 ( .A(_3638__55_), .Y(addr3_o[55]) );
BUFX2 BUFX2_192 ( .A(_3638__54_), .Y(addr3_o[54]) );
BUFX2 BUFX2_193 ( .A(_3639__63_), .Y(addr4_o[63]) );
BUFX2 BUFX2_194 ( .A(_3639__62_), .Y(addr4_o[62]) );
BUFX2 BUFX2_195 ( .A(_3639__53_), .Y(addr4_o[53]) );
BUFX2 BUFX2_196 ( .A(_3639__52_), .Y(addr4_o[52]) );
BUFX2 BUFX2_197 ( .A(_3639__51_), .Y(addr4_o[51]) );
BUFX2 BUFX2_198 ( .A(_3639__50_), .Y(addr4_o[50]) );
BUFX2 BUFX2_199 ( .A(_3639__49_), .Y(addr4_o[49]) );
BUFX2 BUFX2_200 ( .A(_3639__48_), .Y(addr4_o[48]) );
BUFX2 BUFX2_201 ( .A(_3639__47_), .Y(addr4_o[47]) );
BUFX2 BUFX2_202 ( .A(_3639__46_), .Y(addr4_o[46]) );
BUFX2 BUFX2_203 ( .A(_3639__45_), .Y(addr4_o[45]) );
BUFX2 BUFX2_204 ( .A(_3639__44_), .Y(addr4_o[44]) );
BUFX2 BUFX2_205 ( .A(_3639__61_), .Y(addr4_o[61]) );
BUFX2 BUFX2_206 ( .A(_3639__43_), .Y(addr4_o[43]) );
BUFX2 BUFX2_207 ( .A(_3639__42_), .Y(addr4_o[42]) );
BUFX2 BUFX2_208 ( .A(_3639__41_), .Y(addr4_o[41]) );
BUFX2 BUFX2_209 ( .A(_3639__40_), .Y(addr4_o[40]) );
BUFX2 BUFX2_210 ( .A(_3639__39_), .Y(addr4_o[39]) );
BUFX2 BUFX2_211 ( .A(_3639__38_), .Y(addr4_o[38]) );
BUFX2 BUFX2_212 ( .A(_3639__37_), .Y(addr4_o[37]) );
BUFX2 BUFX2_213 ( .A(_3639__36_), .Y(addr4_o[36]) );
BUFX2 BUFX2_214 ( .A(_3639__35_), .Y(addr4_o[35]) );
BUFX2 BUFX2_215 ( .A(_3639__34_), .Y(addr4_o[34]) );
BUFX2 BUFX2_216 ( .A(_3639__60_), .Y(addr4_o[60]) );
BUFX2 BUFX2_217 ( .A(_3639__33_), .Y(addr4_o[33]) );
BUFX2 BUFX2_218 ( .A(_3639__32_), .Y(addr4_o[32]) );
BUFX2 BUFX2_219 ( .A(_3639__31_), .Y(addr4_o[31]) );
BUFX2 BUFX2_220 ( .A(_3639__30_), .Y(addr4_o[30]) );
BUFX2 BUFX2_221 ( .A(_3639__29_), .Y(addr4_o[29]) );
BUFX2 BUFX2_222 ( .A(_3639__28_), .Y(addr4_o[28]) );
BUFX2 BUFX2_223 ( .A(_3639__27_), .Y(addr4_o[27]) );
BUFX2 BUFX2_224 ( .A(_3639__26_), .Y(addr4_o[26]) );
BUFX2 BUFX2_225 ( .A(_3639__25_), .Y(addr4_o[25]) );
BUFX2 BUFX2_226 ( .A(_3639__24_), .Y(addr4_o[24]) );
BUFX2 BUFX2_227 ( .A(_3639__59_), .Y(addr4_o[59]) );
BUFX2 BUFX2_228 ( .A(_3639__23_), .Y(addr4_o[23]) );
BUFX2 BUFX2_229 ( .A(_3639__22_), .Y(addr4_o[22]) );
BUFX2 BUFX2_230 ( .A(_3639__21_), .Y(addr4_o[21]) );
BUFX2 BUFX2_231 ( .A(_3639__20_), .Y(addr4_o[20]) );
BUFX2 BUFX2_232 ( .A(_3639__19_), .Y(addr4_o[19]) );
BUFX2 BUFX2_233 ( .A(_3639__18_), .Y(addr4_o[18]) );
BUFX2 BUFX2_234 ( .A(_3639__17_), .Y(addr4_o[17]) );
BUFX2 BUFX2_235 ( .A(_3639__16_), .Y(addr4_o[16]) );
BUFX2 BUFX2_236 ( .A(_3639__15_), .Y(addr4_o[15]) );
BUFX2 BUFX2_237 ( .A(_3639__14_), .Y(addr4_o[14]) );
BUFX2 BUFX2_238 ( .A(_3639__58_), .Y(addr4_o[58]) );
BUFX2 BUFX2_239 ( .A(_3639__13_), .Y(addr4_o[13]) );
BUFX2 BUFX2_240 ( .A(_3639__12_), .Y(addr4_o[12]) );
BUFX2 BUFX2_241 ( .A(_3639__11_), .Y(addr4_o[11]) );
BUFX2 BUFX2_242 ( .A(_3639__10_), .Y(addr4_o[10]) );
BUFX2 BUFX2_243 ( .A(_3639__9_), .Y(addr4_o[9]) );
BUFX2 BUFX2_244 ( .A(_3639__8_), .Y(addr4_o[8]) );
BUFX2 BUFX2_245 ( .A(_3639__7_), .Y(addr4_o[7]) );
BUFX2 BUFX2_246 ( .A(_3639__6_), .Y(addr4_o[6]) );
BUFX2 BUFX2_247 ( .A(_3639__5_), .Y(addr4_o[5]) );
BUFX2 BUFX2_248 ( .A(_3639__4_), .Y(addr4_o[4]) );
BUFX2 BUFX2_249 ( .A(_3639__57_), .Y(addr4_o[57]) );
BUFX2 BUFX2_250 ( .A(_3639__3_), .Y(addr4_o[3]) );
BUFX2 BUFX2_251 ( .A(_3639__2_), .Y(addr4_o[2]) );
BUFX2 BUFX2_252 ( .A(_3639__1_), .Y(addr4_o[1]) );
BUFX2 BUFX2_253 ( .A(_3639__0_), .Y(addr4_o[0]) );
BUFX2 BUFX2_254 ( .A(_3639__56_), .Y(addr4_o[56]) );
BUFX2 BUFX2_255 ( .A(_3639__55_), .Y(addr4_o[55]) );
BUFX2 BUFX2_256 ( .A(_3639__54_), .Y(addr4_o[54]) );
BUFX2 BUFX2_257 ( .A(_3640_), .Y(enable1_o) );
BUFX2 BUFX2_258 ( .A(_3641_), .Y(enable2_o) );
BUFX2 BUFX2_259 ( .A(_3642_), .Y(enable3_o) );
BUFX2 BUFX2_260 ( .A(_3643_), .Y(enable4_o) );
BUFX2 BUFX2_261 ( .A(_3644__31_), .Y(instr1_o[31]) );
BUFX2 BUFX2_262 ( .A(_3644__30_), .Y(instr1_o[30]) );
BUFX2 BUFX2_263 ( .A(_3644__21_), .Y(instr1_o[21]) );
BUFX2 BUFX2_264 ( .A(_3644__20_), .Y(instr1_o[20]) );
BUFX2 BUFX2_265 ( .A(_3644__19_), .Y(instr1_o[19]) );
BUFX2 BUFX2_266 ( .A(_3644__18_), .Y(instr1_o[18]) );
BUFX2 BUFX2_267 ( .A(_3644__17_), .Y(instr1_o[17]) );
BUFX2 BUFX2_268 ( .A(_3644__16_), .Y(instr1_o[16]) );
BUFX2 BUFX2_269 ( .A(_3644__15_), .Y(instr1_o[15]) );
BUFX2 BUFX2_270 ( .A(_3644__14_), .Y(instr1_o[14]) );
BUFX2 BUFX2_271 ( .A(_3644__13_), .Y(instr1_o[13]) );
BUFX2 BUFX2_272 ( .A(_3644__12_), .Y(instr1_o[12]) );
BUFX2 BUFX2_273 ( .A(_3644__29_), .Y(instr1_o[29]) );
BUFX2 BUFX2_274 ( .A(_3644__11_), .Y(instr1_o[11]) );
BUFX2 BUFX2_275 ( .A(_3644__10_), .Y(instr1_o[10]) );
BUFX2 BUFX2_276 ( .A(_3644__9_), .Y(instr1_o[9]) );
BUFX2 BUFX2_277 ( .A(_3644__8_), .Y(instr1_o[8]) );
BUFX2 BUFX2_278 ( .A(_3644__7_), .Y(instr1_o[7]) );
BUFX2 BUFX2_279 ( .A(_3644__6_), .Y(instr1_o[6]) );
BUFX2 BUFX2_280 ( .A(_3644__5_), .Y(instr1_o[5]) );
BUFX2 BUFX2_281 ( .A(_3644__4_), .Y(instr1_o[4]) );
BUFX2 BUFX2_282 ( .A(_3644__3_), .Y(instr1_o[3]) );
BUFX2 BUFX2_283 ( .A(_3644__2_), .Y(instr1_o[2]) );
BUFX2 BUFX2_284 ( .A(_3644__28_), .Y(instr1_o[28]) );
BUFX2 BUFX2_285 ( .A(_3644__1_), .Y(instr1_o[1]) );
BUFX2 BUFX2_286 ( .A(_3644__0_), .Y(instr1_o[0]) );
BUFX2 BUFX2_287 ( .A(_3644__27_), .Y(instr1_o[27]) );
BUFX2 BUFX2_288 ( .A(_3644__26_), .Y(instr1_o[26]) );
BUFX2 BUFX2_289 ( .A(_3644__25_), .Y(instr1_o[25]) );
BUFX2 BUFX2_290 ( .A(_3644__24_), .Y(instr1_o[24]) );
BUFX2 BUFX2_291 ( .A(_3644__23_), .Y(instr1_o[23]) );
BUFX2 BUFX2_292 ( .A(_3644__22_), .Y(instr1_o[22]) );
BUFX2 BUFX2_293 ( .A(_3645__31_), .Y(instr2_o[31]) );
BUFX2 BUFX2_294 ( .A(_3645__30_), .Y(instr2_o[30]) );
BUFX2 BUFX2_295 ( .A(_3645__21_), .Y(instr2_o[21]) );
BUFX2 BUFX2_296 ( .A(_3645__20_), .Y(instr2_o[20]) );
BUFX2 BUFX2_297 ( .A(_3645__19_), .Y(instr2_o[19]) );
BUFX2 BUFX2_298 ( .A(_3645__18_), .Y(instr2_o[18]) );
BUFX2 BUFX2_299 ( .A(_3645__17_), .Y(instr2_o[17]) );
BUFX2 BUFX2_300 ( .A(_3645__16_), .Y(instr2_o[16]) );
BUFX2 BUFX2_301 ( .A(_3645__15_), .Y(instr2_o[15]) );
BUFX2 BUFX2_302 ( .A(_3645__14_), .Y(instr2_o[14]) );
BUFX2 BUFX2_303 ( .A(_3645__13_), .Y(instr2_o[13]) );
BUFX2 BUFX2_304 ( .A(_3645__12_), .Y(instr2_o[12]) );
BUFX2 BUFX2_305 ( .A(_3645__29_), .Y(instr2_o[29]) );
BUFX2 BUFX2_306 ( .A(_3645__11_), .Y(instr2_o[11]) );
BUFX2 BUFX2_307 ( .A(_3645__10_), .Y(instr2_o[10]) );
BUFX2 BUFX2_308 ( .A(_3645__9_), .Y(instr2_o[9]) );
BUFX2 BUFX2_309 ( .A(_3645__8_), .Y(instr2_o[8]) );
BUFX2 BUFX2_310 ( .A(_3645__7_), .Y(instr2_o[7]) );
BUFX2 BUFX2_311 ( .A(_3645__6_), .Y(instr2_o[6]) );
BUFX2 BUFX2_312 ( .A(_3645__5_), .Y(instr2_o[5]) );
BUFX2 BUFX2_313 ( .A(_3645__4_), .Y(instr2_o[4]) );
BUFX2 BUFX2_314 ( .A(_3645__3_), .Y(instr2_o[3]) );
BUFX2 BUFX2_315 ( .A(_3645__2_), .Y(instr2_o[2]) );
BUFX2 BUFX2_316 ( .A(_3645__28_), .Y(instr2_o[28]) );
BUFX2 BUFX2_317 ( .A(_3645__1_), .Y(instr2_o[1]) );
BUFX2 BUFX2_318 ( .A(_3645__0_), .Y(instr2_o[0]) );
BUFX2 BUFX2_319 ( .A(_3645__27_), .Y(instr2_o[27]) );
BUFX2 BUFX2_320 ( .A(_3645__26_), .Y(instr2_o[26]) );
BUFX2 BUFX2_321 ( .A(_3645__25_), .Y(instr2_o[25]) );
BUFX2 BUFX2_322 ( .A(_3645__24_), .Y(instr2_o[24]) );
BUFX2 BUFX2_323 ( .A(_3645__23_), .Y(instr2_o[23]) );
BUFX2 BUFX2_324 ( .A(_3645__22_), .Y(instr2_o[22]) );
BUFX2 BUFX2_325 ( .A(_3646__31_), .Y(instr3_o[31]) );
BUFX2 BUFX2_326 ( .A(_3646__30_), .Y(instr3_o[30]) );
BUFX2 BUFX2_327 ( .A(_3646__21_), .Y(instr3_o[21]) );
BUFX2 BUFX2_328 ( .A(_3646__20_), .Y(instr3_o[20]) );
BUFX2 BUFX2_329 ( .A(_3646__19_), .Y(instr3_o[19]) );
BUFX2 BUFX2_330 ( .A(_3646__18_), .Y(instr3_o[18]) );
BUFX2 BUFX2_331 ( .A(_3646__17_), .Y(instr3_o[17]) );
BUFX2 BUFX2_332 ( .A(_3646__16_), .Y(instr3_o[16]) );
BUFX2 BUFX2_333 ( .A(_3646__15_), .Y(instr3_o[15]) );
BUFX2 BUFX2_334 ( .A(_3646__14_), .Y(instr3_o[14]) );
BUFX2 BUFX2_335 ( .A(_3646__13_), .Y(instr3_o[13]) );
BUFX2 BUFX2_336 ( .A(_3646__12_), .Y(instr3_o[12]) );
BUFX2 BUFX2_337 ( .A(_3646__29_), .Y(instr3_o[29]) );
BUFX2 BUFX2_338 ( .A(_3646__11_), .Y(instr3_o[11]) );
BUFX2 BUFX2_339 ( .A(_3646__10_), .Y(instr3_o[10]) );
BUFX2 BUFX2_340 ( .A(_3646__9_), .Y(instr3_o[9]) );
BUFX2 BUFX2_341 ( .A(_3646__8_), .Y(instr3_o[8]) );
BUFX2 BUFX2_342 ( .A(_3646__7_), .Y(instr3_o[7]) );
BUFX2 BUFX2_343 ( .A(_3646__6_), .Y(instr3_o[6]) );
BUFX2 BUFX2_344 ( .A(_3646__5_), .Y(instr3_o[5]) );
BUFX2 BUFX2_345 ( .A(_3646__4_), .Y(instr3_o[4]) );
BUFX2 BUFX2_346 ( .A(_3646__3_), .Y(instr3_o[3]) );
BUFX2 BUFX2_347 ( .A(_3646__2_), .Y(instr3_o[2]) );
BUFX2 BUFX2_348 ( .A(_3646__28_), .Y(instr3_o[28]) );
BUFX2 BUFX2_349 ( .A(_3646__1_), .Y(instr3_o[1]) );
BUFX2 BUFX2_350 ( .A(_3646__0_), .Y(instr3_o[0]) );
BUFX2 BUFX2_351 ( .A(_3646__27_), .Y(instr3_o[27]) );
BUFX2 BUFX2_352 ( .A(_3646__26_), .Y(instr3_o[26]) );
BUFX2 BUFX2_353 ( .A(_3646__25_), .Y(instr3_o[25]) );
BUFX2 BUFX2_354 ( .A(_3646__24_), .Y(instr3_o[24]) );
BUFX2 BUFX2_355 ( .A(_3646__23_), .Y(instr3_o[23]) );
BUFX2 BUFX2_356 ( .A(_3646__22_), .Y(instr3_o[22]) );
BUFX2 BUFX2_357 ( .A(_3647__31_), .Y(instr4_o[31]) );
BUFX2 BUFX2_358 ( .A(_3647__30_), .Y(instr4_o[30]) );
BUFX2 BUFX2_359 ( .A(_3647__21_), .Y(instr4_o[21]) );
BUFX2 BUFX2_360 ( .A(_3647__20_), .Y(instr4_o[20]) );
BUFX2 BUFX2_361 ( .A(_3647__19_), .Y(instr4_o[19]) );
BUFX2 BUFX2_362 ( .A(_3647__18_), .Y(instr4_o[18]) );
BUFX2 BUFX2_363 ( .A(_3647__17_), .Y(instr4_o[17]) );
BUFX2 BUFX2_364 ( .A(_3647__16_), .Y(instr4_o[16]) );
BUFX2 BUFX2_365 ( .A(_3647__15_), .Y(instr4_o[15]) );
BUFX2 BUFX2_366 ( .A(_3647__14_), .Y(instr4_o[14]) );
BUFX2 BUFX2_367 ( .A(_3647__13_), .Y(instr4_o[13]) );
BUFX2 BUFX2_368 ( .A(_3647__12_), .Y(instr4_o[12]) );
BUFX2 BUFX2_369 ( .A(_3647__29_), .Y(instr4_o[29]) );
BUFX2 BUFX2_370 ( .A(_3647__11_), .Y(instr4_o[11]) );
BUFX2 BUFX2_371 ( .A(_3647__10_), .Y(instr4_o[10]) );
BUFX2 BUFX2_372 ( .A(_3647__9_), .Y(instr4_o[9]) );
BUFX2 BUFX2_373 ( .A(_3647__8_), .Y(instr4_o[8]) );
BUFX2 BUFX2_374 ( .A(_3647__7_), .Y(instr4_o[7]) );
BUFX2 BUFX2_375 ( .A(_3647__6_), .Y(instr4_o[6]) );
BUFX2 BUFX2_376 ( .A(_3647__5_), .Y(instr4_o[5]) );
BUFX2 BUFX2_377 ( .A(_3647__4_), .Y(instr4_o[4]) );
BUFX2 BUFX2_378 ( .A(_3647__3_), .Y(instr4_o[3]) );
BUFX2 BUFX2_379 ( .A(_3647__2_), .Y(instr4_o[2]) );
BUFX2 BUFX2_380 ( .A(_3647__28_), .Y(instr4_o[28]) );
BUFX2 BUFX2_381 ( .A(_3647__1_), .Y(instr4_o[1]) );
BUFX2 BUFX2_382 ( .A(_3647__0_), .Y(instr4_o[0]) );
BUFX2 BUFX2_383 ( .A(_3647__27_), .Y(instr4_o[27]) );
BUFX2 BUFX2_384 ( .A(_3647__26_), .Y(instr4_o[26]) );
BUFX2 BUFX2_385 ( .A(_3647__25_), .Y(instr4_o[25]) );
BUFX2 BUFX2_386 ( .A(_3647__24_), .Y(instr4_o[24]) );
BUFX2 BUFX2_387 ( .A(_3647__23_), .Y(instr4_o[23]) );
BUFX2 BUFX2_388 ( .A(_3647__22_), .Y(instr4_o[22]) );
BUFX2 BUFX2_389 ( .A(_3648_), .Y(is64b1_o) );
BUFX2 BUFX2_390 ( .A(_3649_), .Y(is64b2_o) );
BUFX2 BUFX2_391 ( .A(_3650_), .Y(is64b3_o) );
BUFX2 BUFX2_392 ( .A(_3651_), .Y(is64b4_o) );
BUFX2 BUFX2_393 ( .A(_3652__63_), .Y(majID1_o[63]) );
BUFX2 BUFX2_394 ( .A(_3652__62_), .Y(majID1_o[62]) );
BUFX2 BUFX2_395 ( .A(_3652__53_), .Y(majID1_o[53]) );
BUFX2 BUFX2_396 ( .A(_3652__52_), .Y(majID1_o[52]) );
BUFX2 BUFX2_397 ( .A(_3652__51_), .Y(majID1_o[51]) );
BUFX2 BUFX2_398 ( .A(_3652__50_), .Y(majID1_o[50]) );
BUFX2 BUFX2_399 ( .A(_3652__49_), .Y(majID1_o[49]) );
BUFX2 BUFX2_400 ( .A(_3652__48_), .Y(majID1_o[48]) );
BUFX2 BUFX2_401 ( .A(_3652__47_), .Y(majID1_o[47]) );
BUFX2 BUFX2_402 ( .A(_3652__46_), .Y(majID1_o[46]) );
BUFX2 BUFX2_403 ( .A(_3652__45_), .Y(majID1_o[45]) );
BUFX2 BUFX2_404 ( .A(_3652__44_), .Y(majID1_o[44]) );
BUFX2 BUFX2_405 ( .A(_3652__61_), .Y(majID1_o[61]) );
BUFX2 BUFX2_406 ( .A(_3652__43_), .Y(majID1_o[43]) );
BUFX2 BUFX2_407 ( .A(_3652__42_), .Y(majID1_o[42]) );
BUFX2 BUFX2_408 ( .A(_3652__41_), .Y(majID1_o[41]) );
BUFX2 BUFX2_409 ( .A(_3652__40_), .Y(majID1_o[40]) );
BUFX2 BUFX2_410 ( .A(_3652__39_), .Y(majID1_o[39]) );
BUFX2 BUFX2_411 ( .A(_3652__38_), .Y(majID1_o[38]) );
BUFX2 BUFX2_412 ( .A(_3652__37_), .Y(majID1_o[37]) );
BUFX2 BUFX2_413 ( .A(_3652__36_), .Y(majID1_o[36]) );
BUFX2 BUFX2_414 ( .A(_3652__35_), .Y(majID1_o[35]) );
BUFX2 BUFX2_415 ( .A(_3652__34_), .Y(majID1_o[34]) );
BUFX2 BUFX2_416 ( .A(_3652__60_), .Y(majID1_o[60]) );
BUFX2 BUFX2_417 ( .A(_3652__33_), .Y(majID1_o[33]) );
BUFX2 BUFX2_418 ( .A(_3652__32_), .Y(majID1_o[32]) );
BUFX2 BUFX2_419 ( .A(_3652__31_), .Y(majID1_o[31]) );
BUFX2 BUFX2_420 ( .A(_3652__30_), .Y(majID1_o[30]) );
BUFX2 BUFX2_421 ( .A(_3652__29_), .Y(majID1_o[29]) );
BUFX2 BUFX2_422 ( .A(_3652__28_), .Y(majID1_o[28]) );
BUFX2 BUFX2_423 ( .A(_3652__27_), .Y(majID1_o[27]) );
BUFX2 BUFX2_424 ( .A(_3652__26_), .Y(majID1_o[26]) );
BUFX2 BUFX2_425 ( .A(_3652__25_), .Y(majID1_o[25]) );
BUFX2 BUFX2_426 ( .A(_3652__24_), .Y(majID1_o[24]) );
BUFX2 BUFX2_427 ( .A(_3652__59_), .Y(majID1_o[59]) );
BUFX2 BUFX2_428 ( .A(_3652__23_), .Y(majID1_o[23]) );
BUFX2 BUFX2_429 ( .A(_3652__22_), .Y(majID1_o[22]) );
BUFX2 BUFX2_430 ( .A(_3652__21_), .Y(majID1_o[21]) );
BUFX2 BUFX2_431 ( .A(_3652__20_), .Y(majID1_o[20]) );
BUFX2 BUFX2_432 ( .A(_3652__19_), .Y(majID1_o[19]) );
BUFX2 BUFX2_433 ( .A(_3652__18_), .Y(majID1_o[18]) );
BUFX2 BUFX2_434 ( .A(_3652__17_), .Y(majID1_o[17]) );
BUFX2 BUFX2_435 ( .A(_3652__16_), .Y(majID1_o[16]) );
BUFX2 BUFX2_436 ( .A(_3652__15_), .Y(majID1_o[15]) );
BUFX2 BUFX2_437 ( .A(_3652__14_), .Y(majID1_o[14]) );
BUFX2 BUFX2_438 ( .A(_3652__58_), .Y(majID1_o[58]) );
BUFX2 BUFX2_439 ( .A(_3652__13_), .Y(majID1_o[13]) );
BUFX2 BUFX2_440 ( .A(_3652__12_), .Y(majID1_o[12]) );
BUFX2 BUFX2_441 ( .A(_3652__11_), .Y(majID1_o[11]) );
BUFX2 BUFX2_442 ( .A(_3652__10_), .Y(majID1_o[10]) );
BUFX2 BUFX2_443 ( .A(_3652__9_), .Y(majID1_o[9]) );
BUFX2 BUFX2_444 ( .A(_3652__8_), .Y(majID1_o[8]) );
BUFX2 BUFX2_445 ( .A(_3652__7_), .Y(majID1_o[7]) );
BUFX2 BUFX2_446 ( .A(_3652__6_), .Y(majID1_o[6]) );
BUFX2 BUFX2_447 ( .A(_3652__5_), .Y(majID1_o[5]) );
BUFX2 BUFX2_448 ( .A(_3652__4_), .Y(majID1_o[4]) );
BUFX2 BUFX2_449 ( .A(_3652__57_), .Y(majID1_o[57]) );
BUFX2 BUFX2_450 ( .A(_3652__3_), .Y(majID1_o[3]) );
BUFX2 BUFX2_451 ( .A(_3652__2_), .Y(majID1_o[2]) );
BUFX2 BUFX2_452 ( .A(_3652__1_), .Y(majID1_o[1]) );
BUFX2 BUFX2_453 ( .A(_3652__0_), .Y(majID1_o[0]) );
BUFX2 BUFX2_454 ( .A(_3652__56_), .Y(majID1_o[56]) );
BUFX2 BUFX2_455 ( .A(_3652__55_), .Y(majID1_o[55]) );
BUFX2 BUFX2_456 ( .A(_3652__54_), .Y(majID1_o[54]) );
BUFX2 BUFX2_457 ( .A(_3653__63_), .Y(majID2_o[63]) );
BUFX2 BUFX2_458 ( .A(_3653__62_), .Y(majID2_o[62]) );
BUFX2 BUFX2_459 ( .A(_3653__53_), .Y(majID2_o[53]) );
BUFX2 BUFX2_460 ( .A(_3653__52_), .Y(majID2_o[52]) );
BUFX2 BUFX2_461 ( .A(_3653__51_), .Y(majID2_o[51]) );
BUFX2 BUFX2_462 ( .A(_3653__50_), .Y(majID2_o[50]) );
BUFX2 BUFX2_463 ( .A(_3653__49_), .Y(majID2_o[49]) );
BUFX2 BUFX2_464 ( .A(_3653__48_), .Y(majID2_o[48]) );
BUFX2 BUFX2_465 ( .A(_3653__47_), .Y(majID2_o[47]) );
BUFX2 BUFX2_466 ( .A(_3653__46_), .Y(majID2_o[46]) );
BUFX2 BUFX2_467 ( .A(_3653__45_), .Y(majID2_o[45]) );
BUFX2 BUFX2_468 ( .A(_3653__44_), .Y(majID2_o[44]) );
BUFX2 BUFX2_469 ( .A(_3653__61_), .Y(majID2_o[61]) );
BUFX2 BUFX2_470 ( .A(_3653__43_), .Y(majID2_o[43]) );
BUFX2 BUFX2_471 ( .A(_3653__42_), .Y(majID2_o[42]) );
BUFX2 BUFX2_472 ( .A(_3653__41_), .Y(majID2_o[41]) );
BUFX2 BUFX2_473 ( .A(_3653__40_), .Y(majID2_o[40]) );
BUFX2 BUFX2_474 ( .A(_3653__39_), .Y(majID2_o[39]) );
BUFX2 BUFX2_475 ( .A(_3653__38_), .Y(majID2_o[38]) );
BUFX2 BUFX2_476 ( .A(_3653__37_), .Y(majID2_o[37]) );
BUFX2 BUFX2_477 ( .A(_3653__36_), .Y(majID2_o[36]) );
BUFX2 BUFX2_478 ( .A(_3653__35_), .Y(majID2_o[35]) );
BUFX2 BUFX2_479 ( .A(_3653__34_), .Y(majID2_o[34]) );
BUFX2 BUFX2_480 ( .A(_3653__60_), .Y(majID2_o[60]) );
BUFX2 BUFX2_481 ( .A(_3653__33_), .Y(majID2_o[33]) );
BUFX2 BUFX2_482 ( .A(_3653__32_), .Y(majID2_o[32]) );
BUFX2 BUFX2_483 ( .A(_3653__31_), .Y(majID2_o[31]) );
BUFX2 BUFX2_484 ( .A(_3653__30_), .Y(majID2_o[30]) );
BUFX2 BUFX2_485 ( .A(_3653__29_), .Y(majID2_o[29]) );
BUFX2 BUFX2_486 ( .A(_3653__28_), .Y(majID2_o[28]) );
BUFX2 BUFX2_487 ( .A(_3653__27_), .Y(majID2_o[27]) );
BUFX2 BUFX2_488 ( .A(_3653__26_), .Y(majID2_o[26]) );
BUFX2 BUFX2_489 ( .A(_3653__25_), .Y(majID2_o[25]) );
BUFX2 BUFX2_490 ( .A(_3653__24_), .Y(majID2_o[24]) );
BUFX2 BUFX2_491 ( .A(_3653__59_), .Y(majID2_o[59]) );
BUFX2 BUFX2_492 ( .A(_3653__23_), .Y(majID2_o[23]) );
BUFX2 BUFX2_493 ( .A(_3653__22_), .Y(majID2_o[22]) );
BUFX2 BUFX2_494 ( .A(_3653__21_), .Y(majID2_o[21]) );
BUFX2 BUFX2_495 ( .A(_3653__20_), .Y(majID2_o[20]) );
BUFX2 BUFX2_496 ( .A(_3653__19_), .Y(majID2_o[19]) );
BUFX2 BUFX2_497 ( .A(_3653__18_), .Y(majID2_o[18]) );
BUFX2 BUFX2_498 ( .A(_3653__17_), .Y(majID2_o[17]) );
BUFX2 BUFX2_499 ( .A(_3653__16_), .Y(majID2_o[16]) );
BUFX2 BUFX2_500 ( .A(_3653__15_), .Y(majID2_o[15]) );
BUFX2 BUFX2_501 ( .A(_3653__14_), .Y(majID2_o[14]) );
BUFX2 BUFX2_502 ( .A(_3653__58_), .Y(majID2_o[58]) );
BUFX2 BUFX2_503 ( .A(_3653__13_), .Y(majID2_o[13]) );
BUFX2 BUFX2_504 ( .A(_3653__12_), .Y(majID2_o[12]) );
BUFX2 BUFX2_505 ( .A(_3653__11_), .Y(majID2_o[11]) );
BUFX2 BUFX2_506 ( .A(_3653__10_), .Y(majID2_o[10]) );
BUFX2 BUFX2_507 ( .A(_3653__9_), .Y(majID2_o[9]) );
BUFX2 BUFX2_508 ( .A(_3653__8_), .Y(majID2_o[8]) );
BUFX2 BUFX2_509 ( .A(_3653__7_), .Y(majID2_o[7]) );
BUFX2 BUFX2_510 ( .A(_3653__6_), .Y(majID2_o[6]) );
BUFX2 BUFX2_511 ( .A(_3653__5_), .Y(majID2_o[5]) );
BUFX2 BUFX2_512 ( .A(_3653__4_), .Y(majID2_o[4]) );
BUFX2 BUFX2_513 ( .A(_3653__57_), .Y(majID2_o[57]) );
BUFX2 BUFX2_514 ( .A(_3653__3_), .Y(majID2_o[3]) );
BUFX2 BUFX2_515 ( .A(_3653__2_), .Y(majID2_o[2]) );
BUFX2 BUFX2_516 ( .A(_3653__1_), .Y(majID2_o[1]) );
BUFX2 BUFX2_517 ( .A(_3653__0_), .Y(majID2_o[0]) );
BUFX2 BUFX2_518 ( .A(_3653__56_), .Y(majID2_o[56]) );
BUFX2 BUFX2_519 ( .A(_3653__55_), .Y(majID2_o[55]) );
BUFX2 BUFX2_520 ( .A(_3653__54_), .Y(majID2_o[54]) );
BUFX2 BUFX2_521 ( .A(_3654__63_), .Y(majID3_o[63]) );
BUFX2 BUFX2_522 ( .A(_3654__62_), .Y(majID3_o[62]) );
BUFX2 BUFX2_523 ( .A(_3654__53_), .Y(majID3_o[53]) );
BUFX2 BUFX2_524 ( .A(_3654__52_), .Y(majID3_o[52]) );
BUFX2 BUFX2_525 ( .A(_3654__51_), .Y(majID3_o[51]) );
BUFX2 BUFX2_526 ( .A(_3654__50_), .Y(majID3_o[50]) );
BUFX2 BUFX2_527 ( .A(_3654__49_), .Y(majID3_o[49]) );
BUFX2 BUFX2_528 ( .A(_3654__48_), .Y(majID3_o[48]) );
BUFX2 BUFX2_529 ( .A(_3654__47_), .Y(majID3_o[47]) );
BUFX2 BUFX2_530 ( .A(_3654__46_), .Y(majID3_o[46]) );
BUFX2 BUFX2_531 ( .A(_3654__45_), .Y(majID3_o[45]) );
BUFX2 BUFX2_532 ( .A(_3654__44_), .Y(majID3_o[44]) );
BUFX2 BUFX2_533 ( .A(_3654__61_), .Y(majID3_o[61]) );
BUFX2 BUFX2_534 ( .A(_3654__43_), .Y(majID3_o[43]) );
BUFX2 BUFX2_535 ( .A(_3654__42_), .Y(majID3_o[42]) );
BUFX2 BUFX2_536 ( .A(_3654__41_), .Y(majID3_o[41]) );
BUFX2 BUFX2_537 ( .A(_3654__40_), .Y(majID3_o[40]) );
BUFX2 BUFX2_538 ( .A(_3654__39_), .Y(majID3_o[39]) );
BUFX2 BUFX2_539 ( .A(_3654__38_), .Y(majID3_o[38]) );
BUFX2 BUFX2_540 ( .A(_3654__37_), .Y(majID3_o[37]) );
BUFX2 BUFX2_541 ( .A(_3654__36_), .Y(majID3_o[36]) );
BUFX2 BUFX2_542 ( .A(_3654__35_), .Y(majID3_o[35]) );
BUFX2 BUFX2_543 ( .A(_3654__34_), .Y(majID3_o[34]) );
BUFX2 BUFX2_544 ( .A(_3654__60_), .Y(majID3_o[60]) );
BUFX2 BUFX2_545 ( .A(_3654__33_), .Y(majID3_o[33]) );
BUFX2 BUFX2_546 ( .A(_3654__32_), .Y(majID3_o[32]) );
BUFX2 BUFX2_547 ( .A(_3654__31_), .Y(majID3_o[31]) );
BUFX2 BUFX2_548 ( .A(_3654__30_), .Y(majID3_o[30]) );
BUFX2 BUFX2_549 ( .A(_3654__29_), .Y(majID3_o[29]) );
BUFX2 BUFX2_550 ( .A(_3654__28_), .Y(majID3_o[28]) );
BUFX2 BUFX2_551 ( .A(_3654__27_), .Y(majID3_o[27]) );
BUFX2 BUFX2_552 ( .A(_3654__26_), .Y(majID3_o[26]) );
BUFX2 BUFX2_553 ( .A(_3654__25_), .Y(majID3_o[25]) );
BUFX2 BUFX2_554 ( .A(_3654__24_), .Y(majID3_o[24]) );
BUFX2 BUFX2_555 ( .A(_3654__59_), .Y(majID3_o[59]) );
BUFX2 BUFX2_556 ( .A(_3654__23_), .Y(majID3_o[23]) );
BUFX2 BUFX2_557 ( .A(_3654__22_), .Y(majID3_o[22]) );
BUFX2 BUFX2_558 ( .A(_3654__21_), .Y(majID3_o[21]) );
BUFX2 BUFX2_559 ( .A(_3654__20_), .Y(majID3_o[20]) );
BUFX2 BUFX2_560 ( .A(_3654__19_), .Y(majID3_o[19]) );
BUFX2 BUFX2_561 ( .A(_3654__18_), .Y(majID3_o[18]) );
BUFX2 BUFX2_562 ( .A(_3654__17_), .Y(majID3_o[17]) );
BUFX2 BUFX2_563 ( .A(_3654__16_), .Y(majID3_o[16]) );
BUFX2 BUFX2_564 ( .A(_3654__15_), .Y(majID3_o[15]) );
BUFX2 BUFX2_565 ( .A(_3654__14_), .Y(majID3_o[14]) );
BUFX2 BUFX2_566 ( .A(_3654__58_), .Y(majID3_o[58]) );
BUFX2 BUFX2_567 ( .A(_3654__13_), .Y(majID3_o[13]) );
BUFX2 BUFX2_568 ( .A(_3654__12_), .Y(majID3_o[12]) );
BUFX2 BUFX2_569 ( .A(_3654__11_), .Y(majID3_o[11]) );
BUFX2 BUFX2_570 ( .A(_3654__10_), .Y(majID3_o[10]) );
BUFX2 BUFX2_571 ( .A(_3654__9_), .Y(majID3_o[9]) );
BUFX2 BUFX2_572 ( .A(_3654__8_), .Y(majID3_o[8]) );
BUFX2 BUFX2_573 ( .A(_3654__7_), .Y(majID3_o[7]) );
BUFX2 BUFX2_574 ( .A(_3654__6_), .Y(majID3_o[6]) );
BUFX2 BUFX2_575 ( .A(_3654__5_), .Y(majID3_o[5]) );
BUFX2 BUFX2_576 ( .A(_3654__4_), .Y(majID3_o[4]) );
BUFX2 BUFX2_577 ( .A(_3654__57_), .Y(majID3_o[57]) );
BUFX2 BUFX2_578 ( .A(_3654__3_), .Y(majID3_o[3]) );
BUFX2 BUFX2_579 ( .A(_3654__2_), .Y(majID3_o[2]) );
BUFX2 BUFX2_580 ( .A(_3654__1_), .Y(majID3_o[1]) );
BUFX2 BUFX2_581 ( .A(_3654__0_), .Y(majID3_o[0]) );
BUFX2 BUFX2_582 ( .A(_3654__56_), .Y(majID3_o[56]) );
BUFX2 BUFX2_583 ( .A(_3654__55_), .Y(majID3_o[55]) );
BUFX2 BUFX2_584 ( .A(_3654__54_), .Y(majID3_o[54]) );
BUFX2 BUFX2_585 ( .A(_3655__63_), .Y(majID4_o[63]) );
BUFX2 BUFX2_586 ( .A(_3655__62_), .Y(majID4_o[62]) );
BUFX2 BUFX2_587 ( .A(_3655__53_), .Y(majID4_o[53]) );
BUFX2 BUFX2_588 ( .A(_3655__52_), .Y(majID4_o[52]) );
BUFX2 BUFX2_589 ( .A(_3655__51_), .Y(majID4_o[51]) );
BUFX2 BUFX2_590 ( .A(_3655__50_), .Y(majID4_o[50]) );
BUFX2 BUFX2_591 ( .A(_3655__49_), .Y(majID4_o[49]) );
BUFX2 BUFX2_592 ( .A(_3655__48_), .Y(majID4_o[48]) );
BUFX2 BUFX2_593 ( .A(_3655__47_), .Y(majID4_o[47]) );
BUFX2 BUFX2_594 ( .A(_3655__46_), .Y(majID4_o[46]) );
BUFX2 BUFX2_595 ( .A(_3655__45_), .Y(majID4_o[45]) );
BUFX2 BUFX2_596 ( .A(_3655__44_), .Y(majID4_o[44]) );
BUFX2 BUFX2_597 ( .A(_3655__61_), .Y(majID4_o[61]) );
BUFX2 BUFX2_598 ( .A(_3655__43_), .Y(majID4_o[43]) );
BUFX2 BUFX2_599 ( .A(_3655__42_), .Y(majID4_o[42]) );
BUFX2 BUFX2_600 ( .A(_3655__41_), .Y(majID4_o[41]) );
BUFX2 BUFX2_601 ( .A(_3655__40_), .Y(majID4_o[40]) );
BUFX2 BUFX2_602 ( .A(_3655__39_), .Y(majID4_o[39]) );
BUFX2 BUFX2_603 ( .A(_3655__38_), .Y(majID4_o[38]) );
BUFX2 BUFX2_604 ( .A(_3655__37_), .Y(majID4_o[37]) );
BUFX2 BUFX2_605 ( .A(_3655__36_), .Y(majID4_o[36]) );
BUFX2 BUFX2_606 ( .A(_3655__35_), .Y(majID4_o[35]) );
BUFX2 BUFX2_607 ( .A(_3655__34_), .Y(majID4_o[34]) );
BUFX2 BUFX2_608 ( .A(_3655__60_), .Y(majID4_o[60]) );
BUFX2 BUFX2_609 ( .A(_3655__33_), .Y(majID4_o[33]) );
BUFX2 BUFX2_610 ( .A(_3655__32_), .Y(majID4_o[32]) );
BUFX2 BUFX2_611 ( .A(_3655__31_), .Y(majID4_o[31]) );
BUFX2 BUFX2_612 ( .A(_3655__30_), .Y(majID4_o[30]) );
BUFX2 BUFX2_613 ( .A(_3655__29_), .Y(majID4_o[29]) );
BUFX2 BUFX2_614 ( .A(_3655__28_), .Y(majID4_o[28]) );
BUFX2 BUFX2_615 ( .A(_3655__27_), .Y(majID4_o[27]) );
BUFX2 BUFX2_616 ( .A(_3655__26_), .Y(majID4_o[26]) );
BUFX2 BUFX2_617 ( .A(_3655__25_), .Y(majID4_o[25]) );
BUFX2 BUFX2_618 ( .A(_3655__24_), .Y(majID4_o[24]) );
BUFX2 BUFX2_619 ( .A(_3655__59_), .Y(majID4_o[59]) );
BUFX2 BUFX2_620 ( .A(_3655__23_), .Y(majID4_o[23]) );
BUFX2 BUFX2_621 ( .A(_3655__22_), .Y(majID4_o[22]) );
BUFX2 BUFX2_622 ( .A(_3655__21_), .Y(majID4_o[21]) );
BUFX2 BUFX2_623 ( .A(_3655__20_), .Y(majID4_o[20]) );
BUFX2 BUFX2_624 ( .A(_3655__19_), .Y(majID4_o[19]) );
BUFX2 BUFX2_625 ( .A(_3655__18_), .Y(majID4_o[18]) );
BUFX2 BUFX2_626 ( .A(_3655__17_), .Y(majID4_o[17]) );
BUFX2 BUFX2_627 ( .A(_3655__16_), .Y(majID4_o[16]) );
BUFX2 BUFX2_628 ( .A(_3655__15_), .Y(majID4_o[15]) );
BUFX2 BUFX2_629 ( .A(_3655__14_), .Y(majID4_o[14]) );
BUFX2 BUFX2_630 ( .A(_3655__58_), .Y(majID4_o[58]) );
BUFX2 BUFX2_631 ( .A(_3655__13_), .Y(majID4_o[13]) );
BUFX2 BUFX2_632 ( .A(_3655__12_), .Y(majID4_o[12]) );
BUFX2 BUFX2_633 ( .A(_3655__11_), .Y(majID4_o[11]) );
BUFX2 BUFX2_634 ( .A(_3655__10_), .Y(majID4_o[10]) );
BUFX2 BUFX2_635 ( .A(_3655__9_), .Y(majID4_o[9]) );
BUFX2 BUFX2_636 ( .A(_3655__8_), .Y(majID4_o[8]) );
BUFX2 BUFX2_637 ( .A(_3655__7_), .Y(majID4_o[7]) );
BUFX2 BUFX2_638 ( .A(_3655__6_), .Y(majID4_o[6]) );
BUFX2 BUFX2_639 ( .A(_3655__5_), .Y(majID4_o[5]) );
BUFX2 BUFX2_640 ( .A(_3655__4_), .Y(majID4_o[4]) );
BUFX2 BUFX2_641 ( .A(_3655__57_), .Y(majID4_o[57]) );
BUFX2 BUFX2_642 ( .A(_3655__3_), .Y(majID4_o[3]) );
BUFX2 BUFX2_643 ( .A(_3655__2_), .Y(majID4_o[2]) );
BUFX2 BUFX2_644 ( .A(_3655__1_), .Y(majID4_o[1]) );
BUFX2 BUFX2_645 ( .A(_3655__0_), .Y(majID4_o[0]) );
BUFX2 BUFX2_646 ( .A(_3655__56_), .Y(majID4_o[56]) );
BUFX2 BUFX2_647 ( .A(_3655__55_), .Y(majID4_o[55]) );
BUFX2 BUFX2_648 ( .A(_3655__54_), .Y(majID4_o[54]) );
BUFX2 BUFX2_649 ( .A(_3656__31_), .Y(pid1_o[31]) );
BUFX2 BUFX2_650 ( .A(_3656__30_), .Y(pid1_o[30]) );
BUFX2 BUFX2_651 ( .A(_3656__21_), .Y(pid1_o[21]) );
BUFX2 BUFX2_652 ( .A(_3656__20_), .Y(pid1_o[20]) );
BUFX2 BUFX2_653 ( .A(_3656__19_), .Y(pid1_o[19]) );
BUFX2 BUFX2_654 ( .A(_3656__18_), .Y(pid1_o[18]) );
BUFX2 BUFX2_655 ( .A(_3656__17_), .Y(pid1_o[17]) );
BUFX2 BUFX2_656 ( .A(_3656__16_), .Y(pid1_o[16]) );
BUFX2 BUFX2_657 ( .A(_3656__15_), .Y(pid1_o[15]) );
BUFX2 BUFX2_658 ( .A(_3656__14_), .Y(pid1_o[14]) );
BUFX2 BUFX2_659 ( .A(_3656__13_), .Y(pid1_o[13]) );
BUFX2 BUFX2_660 ( .A(_3656__12_), .Y(pid1_o[12]) );
BUFX2 BUFX2_661 ( .A(_3656__29_), .Y(pid1_o[29]) );
BUFX2 BUFX2_662 ( .A(_3656__11_), .Y(pid1_o[11]) );
BUFX2 BUFX2_663 ( .A(_3656__10_), .Y(pid1_o[10]) );
BUFX2 BUFX2_664 ( .A(_3656__9_), .Y(pid1_o[9]) );
BUFX2 BUFX2_665 ( .A(_3656__8_), .Y(pid1_o[8]) );
BUFX2 BUFX2_666 ( .A(_3656__7_), .Y(pid1_o[7]) );
BUFX2 BUFX2_667 ( .A(_3656__6_), .Y(pid1_o[6]) );
BUFX2 BUFX2_668 ( .A(_3656__5_), .Y(pid1_o[5]) );
BUFX2 BUFX2_669 ( .A(_3656__4_), .Y(pid1_o[4]) );
BUFX2 BUFX2_670 ( .A(_3656__3_), .Y(pid1_o[3]) );
BUFX2 BUFX2_671 ( .A(_3656__2_), .Y(pid1_o[2]) );
BUFX2 BUFX2_672 ( .A(_3656__28_), .Y(pid1_o[28]) );
BUFX2 BUFX2_673 ( .A(_3656__1_), .Y(pid1_o[1]) );
BUFX2 BUFX2_674 ( .A(_3656__0_), .Y(pid1_o[0]) );
BUFX2 BUFX2_675 ( .A(_3656__27_), .Y(pid1_o[27]) );
BUFX2 BUFX2_676 ( .A(_3656__26_), .Y(pid1_o[26]) );
BUFX2 BUFX2_677 ( .A(_3656__25_), .Y(pid1_o[25]) );
BUFX2 BUFX2_678 ( .A(_3656__24_), .Y(pid1_o[24]) );
BUFX2 BUFX2_679 ( .A(_3656__23_), .Y(pid1_o[23]) );
BUFX2 BUFX2_680 ( .A(_3656__22_), .Y(pid1_o[22]) );
BUFX2 BUFX2_681 ( .A(_3657__31_), .Y(pid2_o[31]) );
BUFX2 BUFX2_682 ( .A(_3657__30_), .Y(pid2_o[30]) );
BUFX2 BUFX2_683 ( .A(_3657__21_), .Y(pid2_o[21]) );
BUFX2 BUFX2_684 ( .A(_3657__20_), .Y(pid2_o[20]) );
BUFX2 BUFX2_685 ( .A(_3657__19_), .Y(pid2_o[19]) );
BUFX2 BUFX2_686 ( .A(_3657__18_), .Y(pid2_o[18]) );
BUFX2 BUFX2_687 ( .A(_3657__17_), .Y(pid2_o[17]) );
BUFX2 BUFX2_688 ( .A(_3657__16_), .Y(pid2_o[16]) );
BUFX2 BUFX2_689 ( .A(_3657__15_), .Y(pid2_o[15]) );
BUFX2 BUFX2_690 ( .A(_3657__14_), .Y(pid2_o[14]) );
BUFX2 BUFX2_691 ( .A(_3657__13_), .Y(pid2_o[13]) );
BUFX2 BUFX2_692 ( .A(_3657__12_), .Y(pid2_o[12]) );
BUFX2 BUFX2_693 ( .A(_3657__29_), .Y(pid2_o[29]) );
BUFX2 BUFX2_694 ( .A(_3657__11_), .Y(pid2_o[11]) );
BUFX2 BUFX2_695 ( .A(_3657__10_), .Y(pid2_o[10]) );
BUFX2 BUFX2_696 ( .A(_3657__9_), .Y(pid2_o[9]) );
BUFX2 BUFX2_697 ( .A(_3657__8_), .Y(pid2_o[8]) );
BUFX2 BUFX2_698 ( .A(_3657__7_), .Y(pid2_o[7]) );
BUFX2 BUFX2_699 ( .A(_3657__6_), .Y(pid2_o[6]) );
BUFX2 BUFX2_700 ( .A(_3657__5_), .Y(pid2_o[5]) );
BUFX2 BUFX2_701 ( .A(_3657__4_), .Y(pid2_o[4]) );
BUFX2 BUFX2_702 ( .A(_3657__3_), .Y(pid2_o[3]) );
BUFX2 BUFX2_703 ( .A(_3657__2_), .Y(pid2_o[2]) );
BUFX2 BUFX2_704 ( .A(_3657__28_), .Y(pid2_o[28]) );
BUFX2 BUFX2_705 ( .A(_3657__1_), .Y(pid2_o[1]) );
BUFX2 BUFX2_706 ( .A(_3657__0_), .Y(pid2_o[0]) );
BUFX2 BUFX2_707 ( .A(_3657__27_), .Y(pid2_o[27]) );
BUFX2 BUFX2_708 ( .A(_3657__26_), .Y(pid2_o[26]) );
BUFX2 BUFX2_709 ( .A(_3657__25_), .Y(pid2_o[25]) );
BUFX2 BUFX2_710 ( .A(_3657__24_), .Y(pid2_o[24]) );
BUFX2 BUFX2_711 ( .A(_3657__23_), .Y(pid2_o[23]) );
BUFX2 BUFX2_712 ( .A(_3657__22_), .Y(pid2_o[22]) );
BUFX2 BUFX2_713 ( .A(_3658__31_), .Y(pid3_o[31]) );
BUFX2 BUFX2_714 ( .A(_3658__30_), .Y(pid3_o[30]) );
BUFX2 BUFX2_715 ( .A(_3658__21_), .Y(pid3_o[21]) );
BUFX2 BUFX2_716 ( .A(_3658__20_), .Y(pid3_o[20]) );
BUFX2 BUFX2_717 ( .A(_3658__19_), .Y(pid3_o[19]) );
BUFX2 BUFX2_718 ( .A(_3658__18_), .Y(pid3_o[18]) );
BUFX2 BUFX2_719 ( .A(_3658__17_), .Y(pid3_o[17]) );
BUFX2 BUFX2_720 ( .A(_3658__16_), .Y(pid3_o[16]) );
BUFX2 BUFX2_721 ( .A(_3658__15_), .Y(pid3_o[15]) );
BUFX2 BUFX2_722 ( .A(_3658__14_), .Y(pid3_o[14]) );
BUFX2 BUFX2_723 ( .A(_3658__13_), .Y(pid3_o[13]) );
BUFX2 BUFX2_724 ( .A(_3658__12_), .Y(pid3_o[12]) );
BUFX2 BUFX2_725 ( .A(_3658__29_), .Y(pid3_o[29]) );
BUFX2 BUFX2_726 ( .A(_3658__11_), .Y(pid3_o[11]) );
BUFX2 BUFX2_727 ( .A(_3658__10_), .Y(pid3_o[10]) );
BUFX2 BUFX2_728 ( .A(_3658__9_), .Y(pid3_o[9]) );
BUFX2 BUFX2_729 ( .A(_3658__8_), .Y(pid3_o[8]) );
BUFX2 BUFX2_730 ( .A(_3658__7_), .Y(pid3_o[7]) );
BUFX2 BUFX2_731 ( .A(_3658__6_), .Y(pid3_o[6]) );
BUFX2 BUFX2_732 ( .A(_3658__5_), .Y(pid3_o[5]) );
BUFX2 BUFX2_733 ( .A(_3658__4_), .Y(pid3_o[4]) );
BUFX2 BUFX2_734 ( .A(_3658__3_), .Y(pid3_o[3]) );
BUFX2 BUFX2_735 ( .A(_3658__2_), .Y(pid3_o[2]) );
BUFX2 BUFX2_736 ( .A(_3658__28_), .Y(pid3_o[28]) );
BUFX2 BUFX2_737 ( .A(_3658__1_), .Y(pid3_o[1]) );
BUFX2 BUFX2_738 ( .A(_3658__0_), .Y(pid3_o[0]) );
BUFX2 BUFX2_739 ( .A(_3658__27_), .Y(pid3_o[27]) );
BUFX2 BUFX2_740 ( .A(_3658__26_), .Y(pid3_o[26]) );
BUFX2 BUFX2_741 ( .A(_3658__25_), .Y(pid3_o[25]) );
BUFX2 BUFX2_742 ( .A(_3658__24_), .Y(pid3_o[24]) );
BUFX2 BUFX2_743 ( .A(_3658__23_), .Y(pid3_o[23]) );
BUFX2 BUFX2_744 ( .A(_3658__22_), .Y(pid3_o[22]) );
BUFX2 BUFX2_745 ( .A(_3659__31_), .Y(pid4_o[31]) );
BUFX2 BUFX2_746 ( .A(_3659__30_), .Y(pid4_o[30]) );
BUFX2 BUFX2_747 ( .A(_3659__21_), .Y(pid4_o[21]) );
BUFX2 BUFX2_748 ( .A(_3659__20_), .Y(pid4_o[20]) );
BUFX2 BUFX2_749 ( .A(_3659__19_), .Y(pid4_o[19]) );
BUFX2 BUFX2_750 ( .A(_3659__18_), .Y(pid4_o[18]) );
BUFX2 BUFX2_751 ( .A(_3659__17_), .Y(pid4_o[17]) );
BUFX2 BUFX2_752 ( .A(_3659__16_), .Y(pid4_o[16]) );
BUFX2 BUFX2_753 ( .A(_3659__15_), .Y(pid4_o[15]) );
BUFX2 BUFX2_754 ( .A(_3659__14_), .Y(pid4_o[14]) );
BUFX2 BUFX2_755 ( .A(_3659__13_), .Y(pid4_o[13]) );
BUFX2 BUFX2_756 ( .A(_3659__12_), .Y(pid4_o[12]) );
BUFX2 BUFX2_757 ( .A(_3659__29_), .Y(pid4_o[29]) );
BUFX2 BUFX2_758 ( .A(_3659__11_), .Y(pid4_o[11]) );
BUFX2 BUFX2_759 ( .A(_3659__10_), .Y(pid4_o[10]) );
BUFX2 BUFX2_760 ( .A(_3659__9_), .Y(pid4_o[9]) );
BUFX2 BUFX2_761 ( .A(_3659__8_), .Y(pid4_o[8]) );
BUFX2 BUFX2_762 ( .A(_3659__7_), .Y(pid4_o[7]) );
BUFX2 BUFX2_763 ( .A(_3659__6_), .Y(pid4_o[6]) );
BUFX2 BUFX2_764 ( .A(_3659__5_), .Y(pid4_o[5]) );
BUFX2 BUFX2_765 ( .A(_3659__4_), .Y(pid4_o[4]) );
BUFX2 BUFX2_766 ( .A(_3659__3_), .Y(pid4_o[3]) );
BUFX2 BUFX2_767 ( .A(_3659__2_), .Y(pid4_o[2]) );
BUFX2 BUFX2_768 ( .A(_3659__28_), .Y(pid4_o[28]) );
BUFX2 BUFX2_769 ( .A(_3659__1_), .Y(pid4_o[1]) );
BUFX2 BUFX2_770 ( .A(_3659__0_), .Y(pid4_o[0]) );
BUFX2 BUFX2_771 ( .A(_3659__27_), .Y(pid4_o[27]) );
BUFX2 BUFX2_772 ( .A(_3659__26_), .Y(pid4_o[26]) );
BUFX2 BUFX2_773 ( .A(_3659__25_), .Y(pid4_o[25]) );
BUFX2 BUFX2_774 ( .A(_3659__24_), .Y(pid4_o[24]) );
BUFX2 BUFX2_775 ( .A(_3659__23_), .Y(pid4_o[23]) );
BUFX2 BUFX2_776 ( .A(_3659__22_), .Y(pid4_o[22]) );
BUFX2 BUFX2_777 ( .A(_3660__63_), .Y(tid1_o[63]) );
BUFX2 BUFX2_778 ( .A(_3660__62_), .Y(tid1_o[62]) );
BUFX2 BUFX2_779 ( .A(_3660__53_), .Y(tid1_o[53]) );
BUFX2 BUFX2_780 ( .A(_3660__52_), .Y(tid1_o[52]) );
BUFX2 BUFX2_781 ( .A(_3660__51_), .Y(tid1_o[51]) );
BUFX2 BUFX2_782 ( .A(_3660__50_), .Y(tid1_o[50]) );
BUFX2 BUFX2_783 ( .A(_3660__49_), .Y(tid1_o[49]) );
BUFX2 BUFX2_784 ( .A(_3660__48_), .Y(tid1_o[48]) );
BUFX2 BUFX2_785 ( .A(_3660__47_), .Y(tid1_o[47]) );
BUFX2 BUFX2_786 ( .A(_3660__46_), .Y(tid1_o[46]) );
BUFX2 BUFX2_787 ( .A(_3660__45_), .Y(tid1_o[45]) );
BUFX2 BUFX2_788 ( .A(_3660__44_), .Y(tid1_o[44]) );
BUFX2 BUFX2_789 ( .A(_3660__61_), .Y(tid1_o[61]) );
BUFX2 BUFX2_790 ( .A(_3660__43_), .Y(tid1_o[43]) );
BUFX2 BUFX2_791 ( .A(_3660__42_), .Y(tid1_o[42]) );
BUFX2 BUFX2_792 ( .A(_3660__41_), .Y(tid1_o[41]) );
BUFX2 BUFX2_793 ( .A(_3660__40_), .Y(tid1_o[40]) );
BUFX2 BUFX2_794 ( .A(_3660__39_), .Y(tid1_o[39]) );
BUFX2 BUFX2_795 ( .A(_3660__38_), .Y(tid1_o[38]) );
BUFX2 BUFX2_796 ( .A(_3660__37_), .Y(tid1_o[37]) );
BUFX2 BUFX2_797 ( .A(_3660__36_), .Y(tid1_o[36]) );
BUFX2 BUFX2_798 ( .A(_3660__35_), .Y(tid1_o[35]) );
BUFX2 BUFX2_799 ( .A(_3660__34_), .Y(tid1_o[34]) );
BUFX2 BUFX2_800 ( .A(_3660__60_), .Y(tid1_o[60]) );
BUFX2 BUFX2_801 ( .A(_3660__33_), .Y(tid1_o[33]) );
BUFX2 BUFX2_802 ( .A(_3660__32_), .Y(tid1_o[32]) );
BUFX2 BUFX2_803 ( .A(_3660__31_), .Y(tid1_o[31]) );
BUFX2 BUFX2_804 ( .A(_3660__30_), .Y(tid1_o[30]) );
BUFX2 BUFX2_805 ( .A(_3660__29_), .Y(tid1_o[29]) );
BUFX2 BUFX2_806 ( .A(_3660__28_), .Y(tid1_o[28]) );
BUFX2 BUFX2_807 ( .A(_3660__27_), .Y(tid1_o[27]) );
BUFX2 BUFX2_808 ( .A(_3660__26_), .Y(tid1_o[26]) );
BUFX2 BUFX2_809 ( .A(_3660__25_), .Y(tid1_o[25]) );
BUFX2 BUFX2_810 ( .A(_3660__24_), .Y(tid1_o[24]) );
BUFX2 BUFX2_811 ( .A(_3660__59_), .Y(tid1_o[59]) );
BUFX2 BUFX2_812 ( .A(_3660__23_), .Y(tid1_o[23]) );
BUFX2 BUFX2_813 ( .A(_3660__22_), .Y(tid1_o[22]) );
BUFX2 BUFX2_814 ( .A(_3660__21_), .Y(tid1_o[21]) );
BUFX2 BUFX2_815 ( .A(_3660__20_), .Y(tid1_o[20]) );
BUFX2 BUFX2_816 ( .A(_3660__19_), .Y(tid1_o[19]) );
BUFX2 BUFX2_817 ( .A(_3660__18_), .Y(tid1_o[18]) );
BUFX2 BUFX2_818 ( .A(_3660__17_), .Y(tid1_o[17]) );
BUFX2 BUFX2_819 ( .A(_3660__16_), .Y(tid1_o[16]) );
BUFX2 BUFX2_820 ( .A(_3660__15_), .Y(tid1_o[15]) );
BUFX2 BUFX2_821 ( .A(_3660__14_), .Y(tid1_o[14]) );
BUFX2 BUFX2_822 ( .A(_3660__58_), .Y(tid1_o[58]) );
BUFX2 BUFX2_823 ( .A(_3660__13_), .Y(tid1_o[13]) );
BUFX2 BUFX2_824 ( .A(_3660__12_), .Y(tid1_o[12]) );
BUFX2 BUFX2_825 ( .A(_3660__11_), .Y(tid1_o[11]) );
BUFX2 BUFX2_826 ( .A(_3660__10_), .Y(tid1_o[10]) );
BUFX2 BUFX2_827 ( .A(_3660__9_), .Y(tid1_o[9]) );
BUFX2 BUFX2_828 ( .A(_3660__8_), .Y(tid1_o[8]) );
BUFX2 BUFX2_829 ( .A(_3660__7_), .Y(tid1_o[7]) );
BUFX2 BUFX2_830 ( .A(_3660__6_), .Y(tid1_o[6]) );
BUFX2 BUFX2_831 ( .A(_3660__5_), .Y(tid1_o[5]) );
BUFX2 BUFX2_832 ( .A(_3660__4_), .Y(tid1_o[4]) );
BUFX2 BUFX2_833 ( .A(_3660__57_), .Y(tid1_o[57]) );
BUFX2 BUFX2_834 ( .A(_3660__3_), .Y(tid1_o[3]) );
BUFX2 BUFX2_835 ( .A(_3660__2_), .Y(tid1_o[2]) );
BUFX2 BUFX2_836 ( .A(_3660__1_), .Y(tid1_o[1]) );
BUFX2 BUFX2_837 ( .A(_3660__0_), .Y(tid1_o[0]) );
BUFX2 BUFX2_838 ( .A(_3660__56_), .Y(tid1_o[56]) );
BUFX2 BUFX2_839 ( .A(_3660__55_), .Y(tid1_o[55]) );
BUFX2 BUFX2_840 ( .A(_3660__54_), .Y(tid1_o[54]) );
BUFX2 BUFX2_841 ( .A(_3661__63_), .Y(tid2_o[63]) );
BUFX2 BUFX2_842 ( .A(_3661__62_), .Y(tid2_o[62]) );
BUFX2 BUFX2_843 ( .A(_3661__53_), .Y(tid2_o[53]) );
BUFX2 BUFX2_844 ( .A(_3661__52_), .Y(tid2_o[52]) );
BUFX2 BUFX2_845 ( .A(_3661__51_), .Y(tid2_o[51]) );
BUFX2 BUFX2_846 ( .A(_3661__50_), .Y(tid2_o[50]) );
BUFX2 BUFX2_847 ( .A(_3661__49_), .Y(tid2_o[49]) );
BUFX2 BUFX2_848 ( .A(_3661__48_), .Y(tid2_o[48]) );
BUFX2 BUFX2_849 ( .A(_3661__47_), .Y(tid2_o[47]) );
BUFX2 BUFX2_850 ( .A(_3661__46_), .Y(tid2_o[46]) );
BUFX2 BUFX2_851 ( .A(_3661__45_), .Y(tid2_o[45]) );
BUFX2 BUFX2_852 ( .A(_3661__44_), .Y(tid2_o[44]) );
BUFX2 BUFX2_853 ( .A(_3661__61_), .Y(tid2_o[61]) );
BUFX2 BUFX2_854 ( .A(_3661__43_), .Y(tid2_o[43]) );
BUFX2 BUFX2_855 ( .A(_3661__42_), .Y(tid2_o[42]) );
BUFX2 BUFX2_856 ( .A(_3661__41_), .Y(tid2_o[41]) );
BUFX2 BUFX2_857 ( .A(_3661__40_), .Y(tid2_o[40]) );
BUFX2 BUFX2_858 ( .A(_3661__39_), .Y(tid2_o[39]) );
BUFX2 BUFX2_859 ( .A(_3661__38_), .Y(tid2_o[38]) );
BUFX2 BUFX2_860 ( .A(_3661__37_), .Y(tid2_o[37]) );
BUFX2 BUFX2_861 ( .A(_3661__36_), .Y(tid2_o[36]) );
BUFX2 BUFX2_862 ( .A(_3661__35_), .Y(tid2_o[35]) );
BUFX2 BUFX2_863 ( .A(_3661__34_), .Y(tid2_o[34]) );
BUFX2 BUFX2_864 ( .A(_3661__60_), .Y(tid2_o[60]) );
BUFX2 BUFX2_865 ( .A(_3661__33_), .Y(tid2_o[33]) );
BUFX2 BUFX2_866 ( .A(_3661__32_), .Y(tid2_o[32]) );
BUFX2 BUFX2_867 ( .A(_3661__31_), .Y(tid2_o[31]) );
BUFX2 BUFX2_868 ( .A(_3661__30_), .Y(tid2_o[30]) );
BUFX2 BUFX2_869 ( .A(_3661__29_), .Y(tid2_o[29]) );
BUFX2 BUFX2_870 ( .A(_3661__28_), .Y(tid2_o[28]) );
BUFX2 BUFX2_871 ( .A(_3661__27_), .Y(tid2_o[27]) );
BUFX2 BUFX2_872 ( .A(_3661__26_), .Y(tid2_o[26]) );
BUFX2 BUFX2_873 ( .A(_3661__25_), .Y(tid2_o[25]) );
BUFX2 BUFX2_874 ( .A(_3661__24_), .Y(tid2_o[24]) );
BUFX2 BUFX2_875 ( .A(_3661__59_), .Y(tid2_o[59]) );
BUFX2 BUFX2_876 ( .A(_3661__23_), .Y(tid2_o[23]) );
BUFX2 BUFX2_877 ( .A(_3661__22_), .Y(tid2_o[22]) );
BUFX2 BUFX2_878 ( .A(_3661__21_), .Y(tid2_o[21]) );
BUFX2 BUFX2_879 ( .A(_3661__20_), .Y(tid2_o[20]) );
BUFX2 BUFX2_880 ( .A(_3661__19_), .Y(tid2_o[19]) );
BUFX2 BUFX2_881 ( .A(_3661__18_), .Y(tid2_o[18]) );
BUFX2 BUFX2_882 ( .A(_3661__17_), .Y(tid2_o[17]) );
BUFX2 BUFX2_883 ( .A(_3661__16_), .Y(tid2_o[16]) );
BUFX2 BUFX2_884 ( .A(_3661__15_), .Y(tid2_o[15]) );
BUFX2 BUFX2_885 ( .A(_3661__14_), .Y(tid2_o[14]) );
BUFX2 BUFX2_886 ( .A(_3661__58_), .Y(tid2_o[58]) );
BUFX2 BUFX2_887 ( .A(_3661__13_), .Y(tid2_o[13]) );
BUFX2 BUFX2_888 ( .A(_3661__12_), .Y(tid2_o[12]) );
BUFX2 BUFX2_889 ( .A(_3661__11_), .Y(tid2_o[11]) );
BUFX2 BUFX2_890 ( .A(_3661__10_), .Y(tid2_o[10]) );
BUFX2 BUFX2_891 ( .A(_3661__9_), .Y(tid2_o[9]) );
BUFX2 BUFX2_892 ( .A(_3661__8_), .Y(tid2_o[8]) );
BUFX2 BUFX2_893 ( .A(_3661__7_), .Y(tid2_o[7]) );
BUFX2 BUFX2_894 ( .A(_3661__6_), .Y(tid2_o[6]) );
BUFX2 BUFX2_895 ( .A(_3661__5_), .Y(tid2_o[5]) );
BUFX2 BUFX2_896 ( .A(_3661__4_), .Y(tid2_o[4]) );
BUFX2 BUFX2_897 ( .A(_3661__57_), .Y(tid2_o[57]) );
BUFX2 BUFX2_898 ( .A(_3661__3_), .Y(tid2_o[3]) );
BUFX2 BUFX2_899 ( .A(_3661__2_), .Y(tid2_o[2]) );
BUFX2 BUFX2_900 ( .A(_3661__1_), .Y(tid2_o[1]) );
BUFX2 BUFX2_901 ( .A(_3661__0_), .Y(tid2_o[0]) );
BUFX2 BUFX2_902 ( .A(_3661__56_), .Y(tid2_o[56]) );
BUFX2 BUFX2_903 ( .A(_3661__55_), .Y(tid2_o[55]) );
BUFX2 BUFX2_904 ( .A(_3661__54_), .Y(tid2_o[54]) );
BUFX2 BUFX2_905 ( .A(_3662__63_), .Y(tid3_o[63]) );
BUFX2 BUFX2_906 ( .A(_3662__62_), .Y(tid3_o[62]) );
BUFX2 BUFX2_907 ( .A(_3662__53_), .Y(tid3_o[53]) );
BUFX2 BUFX2_908 ( .A(_3662__52_), .Y(tid3_o[52]) );
BUFX2 BUFX2_909 ( .A(_3662__51_), .Y(tid3_o[51]) );
BUFX2 BUFX2_910 ( .A(_3662__50_), .Y(tid3_o[50]) );
BUFX2 BUFX2_911 ( .A(_3662__49_), .Y(tid3_o[49]) );
BUFX2 BUFX2_912 ( .A(_3662__48_), .Y(tid3_o[48]) );
BUFX2 BUFX2_913 ( .A(_3662__47_), .Y(tid3_o[47]) );
BUFX2 BUFX2_914 ( .A(_3662__46_), .Y(tid3_o[46]) );
BUFX2 BUFX2_915 ( .A(_3662__45_), .Y(tid3_o[45]) );
BUFX2 BUFX2_916 ( .A(_3662__44_), .Y(tid3_o[44]) );
BUFX2 BUFX2_917 ( .A(_3662__61_), .Y(tid3_o[61]) );
BUFX2 BUFX2_918 ( .A(_3662__43_), .Y(tid3_o[43]) );
BUFX2 BUFX2_919 ( .A(_3662__42_), .Y(tid3_o[42]) );
BUFX2 BUFX2_920 ( .A(_3662__41_), .Y(tid3_o[41]) );
BUFX2 BUFX2_921 ( .A(_3662__40_), .Y(tid3_o[40]) );
BUFX2 BUFX2_922 ( .A(_3662__39_), .Y(tid3_o[39]) );
BUFX2 BUFX2_923 ( .A(_3662__38_), .Y(tid3_o[38]) );
BUFX2 BUFX2_924 ( .A(_3662__37_), .Y(tid3_o[37]) );
BUFX2 BUFX2_925 ( .A(_3662__36_), .Y(tid3_o[36]) );
BUFX2 BUFX2_926 ( .A(_3662__35_), .Y(tid3_o[35]) );
BUFX2 BUFX2_927 ( .A(_3662__34_), .Y(tid3_o[34]) );
BUFX2 BUFX2_928 ( .A(_3662__60_), .Y(tid3_o[60]) );
BUFX2 BUFX2_929 ( .A(_3662__33_), .Y(tid3_o[33]) );
BUFX2 BUFX2_930 ( .A(_3662__32_), .Y(tid3_o[32]) );
BUFX2 BUFX2_931 ( .A(_3662__31_), .Y(tid3_o[31]) );
BUFX2 BUFX2_932 ( .A(_3662__30_), .Y(tid3_o[30]) );
BUFX2 BUFX2_933 ( .A(_3662__29_), .Y(tid3_o[29]) );
BUFX2 BUFX2_934 ( .A(_3662__28_), .Y(tid3_o[28]) );
BUFX2 BUFX2_935 ( .A(_3662__27_), .Y(tid3_o[27]) );
BUFX2 BUFX2_936 ( .A(_3662__26_), .Y(tid3_o[26]) );
BUFX2 BUFX2_937 ( .A(_3662__25_), .Y(tid3_o[25]) );
BUFX2 BUFX2_938 ( .A(_3662__24_), .Y(tid3_o[24]) );
BUFX2 BUFX2_939 ( .A(_3662__59_), .Y(tid3_o[59]) );
BUFX2 BUFX2_940 ( .A(_3662__23_), .Y(tid3_o[23]) );
BUFX2 BUFX2_941 ( .A(_3662__22_), .Y(tid3_o[22]) );
BUFX2 BUFX2_942 ( .A(_3662__21_), .Y(tid3_o[21]) );
BUFX2 BUFX2_943 ( .A(_3662__20_), .Y(tid3_o[20]) );
BUFX2 BUFX2_944 ( .A(_3662__19_), .Y(tid3_o[19]) );
BUFX2 BUFX2_945 ( .A(_3662__18_), .Y(tid3_o[18]) );
BUFX2 BUFX2_946 ( .A(_3662__17_), .Y(tid3_o[17]) );
BUFX2 BUFX2_947 ( .A(_3662__16_), .Y(tid3_o[16]) );
BUFX2 BUFX2_948 ( .A(_3662__15_), .Y(tid3_o[15]) );
BUFX2 BUFX2_949 ( .A(_3662__14_), .Y(tid3_o[14]) );
BUFX2 BUFX2_950 ( .A(_3662__58_), .Y(tid3_o[58]) );
BUFX2 BUFX2_951 ( .A(_3662__13_), .Y(tid3_o[13]) );
BUFX2 BUFX2_952 ( .A(_3662__12_), .Y(tid3_o[12]) );
BUFX2 BUFX2_953 ( .A(_3662__11_), .Y(tid3_o[11]) );
BUFX2 BUFX2_954 ( .A(_3662__10_), .Y(tid3_o[10]) );
BUFX2 BUFX2_955 ( .A(_3662__9_), .Y(tid3_o[9]) );
BUFX2 BUFX2_956 ( .A(_3662__8_), .Y(tid3_o[8]) );
BUFX2 BUFX2_957 ( .A(_3662__7_), .Y(tid3_o[7]) );
BUFX2 BUFX2_958 ( .A(_3662__6_), .Y(tid3_o[6]) );
BUFX2 BUFX2_959 ( .A(_3662__5_), .Y(tid3_o[5]) );
BUFX2 BUFX2_960 ( .A(_3662__4_), .Y(tid3_o[4]) );
BUFX2 BUFX2_961 ( .A(_3662__57_), .Y(tid3_o[57]) );
BUFX2 BUFX2_962 ( .A(_3662__3_), .Y(tid3_o[3]) );
BUFX2 BUFX2_963 ( .A(_3662__2_), .Y(tid3_o[2]) );
BUFX2 BUFX2_964 ( .A(_3662__1_), .Y(tid3_o[1]) );
BUFX2 BUFX2_965 ( .A(_3662__0_), .Y(tid3_o[0]) );
BUFX2 BUFX2_966 ( .A(_3662__56_), .Y(tid3_o[56]) );
BUFX2 BUFX2_967 ( .A(_3662__55_), .Y(tid3_o[55]) );
BUFX2 BUFX2_968 ( .A(_3662__54_), .Y(tid3_o[54]) );
BUFX2 BUFX2_969 ( .A(_3663__63_), .Y(tid4_o[63]) );
BUFX2 BUFX2_970 ( .A(_3663__62_), .Y(tid4_o[62]) );
BUFX2 BUFX2_971 ( .A(_3663__53_), .Y(tid4_o[53]) );
BUFX2 BUFX2_972 ( .A(_3663__52_), .Y(tid4_o[52]) );
BUFX2 BUFX2_973 ( .A(_3663__51_), .Y(tid4_o[51]) );
BUFX2 BUFX2_974 ( .A(_3663__50_), .Y(tid4_o[50]) );
BUFX2 BUFX2_975 ( .A(_3663__49_), .Y(tid4_o[49]) );
BUFX2 BUFX2_976 ( .A(_3663__48_), .Y(tid4_o[48]) );
BUFX2 BUFX2_977 ( .A(_3663__47_), .Y(tid4_o[47]) );
BUFX2 BUFX2_978 ( .A(_3663__46_), .Y(tid4_o[46]) );
BUFX2 BUFX2_979 ( .A(_3663__45_), .Y(tid4_o[45]) );
BUFX2 BUFX2_980 ( .A(_3663__44_), .Y(tid4_o[44]) );
BUFX2 BUFX2_981 ( .A(_3663__61_), .Y(tid4_o[61]) );
BUFX2 BUFX2_982 ( .A(_3663__43_), .Y(tid4_o[43]) );
BUFX2 BUFX2_983 ( .A(_3663__42_), .Y(tid4_o[42]) );
BUFX2 BUFX2_984 ( .A(_3663__41_), .Y(tid4_o[41]) );
BUFX2 BUFX2_985 ( .A(_3663__40_), .Y(tid4_o[40]) );
BUFX2 BUFX2_986 ( .A(_3663__39_), .Y(tid4_o[39]) );
BUFX2 BUFX2_987 ( .A(_3663__38_), .Y(tid4_o[38]) );
BUFX2 BUFX2_988 ( .A(_3663__37_), .Y(tid4_o[37]) );
BUFX2 BUFX2_989 ( .A(_3663__36_), .Y(tid4_o[36]) );
BUFX2 BUFX2_990 ( .A(_3663__35_), .Y(tid4_o[35]) );
BUFX2 BUFX2_991 ( .A(_3663__34_), .Y(tid4_o[34]) );
BUFX2 BUFX2_992 ( .A(_3663__60_), .Y(tid4_o[60]) );
BUFX2 BUFX2_993 ( .A(_3663__33_), .Y(tid4_o[33]) );
BUFX2 BUFX2_994 ( .A(_3663__32_), .Y(tid4_o[32]) );
BUFX2 BUFX2_995 ( .A(_3663__31_), .Y(tid4_o[31]) );
BUFX2 BUFX2_996 ( .A(_3663__30_), .Y(tid4_o[30]) );
BUFX2 BUFX2_997 ( .A(_3663__29_), .Y(tid4_o[29]) );
BUFX2 BUFX2_998 ( .A(_3663__28_), .Y(tid4_o[28]) );
BUFX2 BUFX2_999 ( .A(_3663__27_), .Y(tid4_o[27]) );
BUFX2 BUFX2_1000 ( .A(_3663__26_), .Y(tid4_o[26]) );
BUFX2 BUFX2_1001 ( .A(_3663__25_), .Y(tid4_o[25]) );
BUFX2 BUFX2_1002 ( .A(_3663__24_), .Y(tid4_o[24]) );
BUFX2 BUFX2_1003 ( .A(_3663__59_), .Y(tid4_o[59]) );
BUFX2 BUFX2_1004 ( .A(_3663__23_), .Y(tid4_o[23]) );
BUFX2 BUFX2_1005 ( .A(_3663__22_), .Y(tid4_o[22]) );
BUFX2 BUFX2_1006 ( .A(_3663__21_), .Y(tid4_o[21]) );
BUFX2 BUFX2_1007 ( .A(_3663__20_), .Y(tid4_o[20]) );
BUFX2 BUFX2_1008 ( .A(_3663__19_), .Y(tid4_o[19]) );
BUFX2 BUFX2_1009 ( .A(_3663__18_), .Y(tid4_o[18]) );
BUFX2 BUFX2_1010 ( .A(_3663__17_), .Y(tid4_o[17]) );
BUFX2 BUFX2_1011 ( .A(_3663__16_), .Y(tid4_o[16]) );
BUFX2 BUFX2_1012 ( .A(_3663__15_), .Y(tid4_o[15]) );
BUFX2 BUFX2_1013 ( .A(_3663__14_), .Y(tid4_o[14]) );
BUFX2 BUFX2_1014 ( .A(_3663__58_), .Y(tid4_o[58]) );
BUFX2 BUFX2_1015 ( .A(_3663__13_), .Y(tid4_o[13]) );
BUFX2 BUFX2_1016 ( .A(_3663__12_), .Y(tid4_o[12]) );
BUFX2 BUFX2_1017 ( .A(_3663__11_), .Y(tid4_o[11]) );
BUFX2 BUFX2_1018 ( .A(_3663__10_), .Y(tid4_o[10]) );
BUFX2 BUFX2_1019 ( .A(_3663__9_), .Y(tid4_o[9]) );
BUFX2 BUFX2_1020 ( .A(_3663__8_), .Y(tid4_o[8]) );
BUFX2 BUFX2_1021 ( .A(_3663__7_), .Y(tid4_o[7]) );
BUFX2 BUFX2_1022 ( .A(_3663__6_), .Y(tid4_o[6]) );
BUFX2 BUFX2_1023 ( .A(_3663__5_), .Y(tid4_o[5]) );
BUFX2 BUFX2_1024 ( .A(_3663__4_), .Y(tid4_o[4]) );
BUFX2 BUFX2_1025 ( .A(_3663__57_), .Y(tid4_o[57]) );
BUFX2 BUFX2_1026 ( .A(_3663__3_), .Y(tid4_o[3]) );
BUFX2 BUFX2_1027 ( .A(_3663__2_), .Y(tid4_o[2]) );
BUFX2 BUFX2_1028 ( .A(_3663__1_), .Y(tid4_o[1]) );
BUFX2 BUFX2_1029 ( .A(_3663__0_), .Y(tid4_o[0]) );
BUFX2 BUFX2_1030 ( .A(_3663__56_), .Y(tid4_o[56]) );
BUFX2 BUFX2_1031 ( .A(_3663__55_), .Y(tid4_o[55]) );
BUFX2 BUFX2_1032 ( .A(_3663__54_), .Y(tid4_o[54]) );
FILL FILL_0_INVX1_103 ( );
FILL FILL_1_INVX1_103 ( );
FILL FILL_0_NAND2X1_368 ( );
FILL FILL_0_OAI21X1_902 ( );
FILL FILL_1_OAI21X1_902 ( );
FILL FILL_0_NAND2X1_396 ( );
FILL FILL_0_DFFPOSX1_674 ( );
FILL FILL_1_DFFPOSX1_674 ( );
FILL FILL_2_DFFPOSX1_674 ( );
FILL FILL_3_DFFPOSX1_674 ( );
FILL FILL_4_DFFPOSX1_674 ( );
FILL FILL_5_DFFPOSX1_674 ( );
FILL FILL_6_DFFPOSX1_674 ( );
FILL FILL_0_BUFX2_312 ( );
FILL FILL_1_BUFX2_312 ( );
FILL FILL_0_NAND2X1_369 ( );
FILL FILL_0_INVX1_86 ( );
FILL FILL_0_BUFX2_324 ( );
FILL FILL_0_OAI21X1_885 ( );
FILL FILL_1_OAI21X1_885 ( );
FILL FILL_0_NAND2X1_379 ( );
FILL FILL_1_NAND2X1_379 ( );
FILL FILL_0_NAND2X1_348 ( );
FILL FILL_1_NAND2X1_348 ( );
FILL FILL_0_BUFX2_286 ( );
FILL FILL_1_BUFX2_286 ( );
FILL FILL_0_DFFPOSX1_657 ( );
FILL FILL_1_DFFPOSX1_657 ( );
FILL FILL_2_DFFPOSX1_657 ( );
FILL FILL_3_DFFPOSX1_657 ( );
FILL FILL_4_DFFPOSX1_657 ( );
FILL FILL_5_DFFPOSX1_657 ( );
FILL FILL_6_DFFPOSX1_657 ( );
FILL FILL_0_BUFX2_263 ( );
FILL FILL_1_BUFX2_263 ( );
FILL FILL_0_NAND2X1_342 ( );
FILL FILL_0_BUFX2_287 ( );
FILL FILL_0_DFFPOSX1_620 ( );
FILL FILL_1_DFFPOSX1_620 ( );
FILL FILL_2_DFFPOSX1_620 ( );
FILL FILL_3_DFFPOSX1_620 ( );
FILL FILL_4_DFFPOSX1_620 ( );
FILL FILL_5_DFFPOSX1_620 ( );
FILL FILL_6_DFFPOSX1_620 ( );
FILL FILL_0_INVX1_49 ( );
FILL FILL_0_OAI21X1_848 ( );
FILL FILL_1_OAI21X1_848 ( );
FILL FILL_2_OAI21X1_848 ( );
FILL FILL_0_BUFX2_846 ( );
FILL FILL_0_BUFX2_309 ( );
FILL FILL_1_BUFX2_309 ( );
FILL FILL_0_NAND2X1_353 ( );
FILL FILL_1_NAND2X1_353 ( );
FILL FILL_0_NAND2X1_359 ( );
FILL FILL_1_NAND2X1_359 ( );
FILL FILL_0_BUFX2_268 ( );
FILL FILL_1_BUFX2_268 ( );
FILL FILL_0_BUFX2_275 ( );
FILL FILL_1_BUFX2_275 ( );
FILL FILL_0_BUFX2_527 ( );
FILL FILL_0_OAI21X1_865 ( );
FILL FILL_1_OAI21X1_865 ( );
FILL FILL_0_INVX1_66 ( );
FILL FILL_0_INVX2_136 ( );
FILL FILL_0_DFFPOSX1_637 ( );
FILL FILL_1_DFFPOSX1_637 ( );
FILL FILL_2_DFFPOSX1_637 ( );
FILL FILL_3_DFFPOSX1_637 ( );
FILL FILL_4_DFFPOSX1_637 ( );
FILL FILL_5_DFFPOSX1_637 ( );
FILL FILL_6_DFFPOSX1_637 ( );
FILL FILL_0_BUFX2_302 ( );
FILL FILL_1_BUFX2_302 ( );
FILL FILL_0_BUFX2_282 ( );
FILL FILL_0_NAND2X1_366 ( );
FILL FILL_1_NAND2X1_366 ( );
FILL FILL_0_INVX1_73 ( );
FILL FILL_0_OAI21X1_872 ( );
FILL FILL_1_OAI21X1_872 ( );
FILL FILL_0_DFFPOSX1_644 ( );
FILL FILL_1_DFFPOSX1_644 ( );
FILL FILL_2_DFFPOSX1_644 ( );
FILL FILL_3_DFFPOSX1_644 ( );
FILL FILL_4_DFFPOSX1_644 ( );
FILL FILL_5_DFFPOSX1_644 ( );
FILL FILL_6_DFFPOSX1_644 ( );
FILL FILL_0_BUFX2_257 ( );
FILL FILL_1_BUFX2_257 ( );
FILL FILL_0_DFFPOSX1_612 ( );
FILL FILL_1_DFFPOSX1_612 ( );
FILL FILL_2_DFFPOSX1_612 ( );
FILL FILL_3_DFFPOSX1_612 ( );
FILL FILL_4_DFFPOSX1_612 ( );
FILL FILL_5_DFFPOSX1_612 ( );
FILL FILL_0_NAND2X1_347 ( );
FILL FILL_1_NAND2X1_347 ( );
FILL FILL_0_BUFX2_292 ( );
FILL FILL_1_BUFX2_292 ( );
FILL FILL_0_DFFPOSX1_625 ( );
FILL FILL_1_DFFPOSX1_625 ( );
FILL FILL_2_DFFPOSX1_625 ( );
FILL FILL_3_DFFPOSX1_625 ( );
FILL FILL_4_DFFPOSX1_625 ( );
FILL FILL_5_DFFPOSX1_625 ( );
FILL FILL_0_OAI21X1_853 ( );
FILL FILL_1_OAI21X1_853 ( );
FILL FILL_0_INVX1_54 ( );
FILL FILL_0_BUFX2_462 ( );
FILL FILL_0_BUFX2_519 ( );
FILL FILL_0_BUFX2_705 ( );
FILL FILL_1_BUFX2_705 ( );
FILL FILL_0_BUFX2_523 ( );
FILL FILL_1_BUFX2_523 ( );
FILL FILL_0_BUFX2_590 ( );
FILL FILL_1_BUFX2_590 ( );
FILL FILL_0_BUFX2_400 ( );
FILL FILL_1_BUFX2_400 ( );
FILL FILL_0_BUFX2_464 ( );
FILL FILL_0_BUFX2_395 ( );
FILL FILL_1_BUFX2_395 ( );
FILL FILL_0_BUFX2_591 ( );
FILL FILL_1_BUFX2_591 ( );
FILL FILL_0_BUFX2_526 ( );
FILL FILL_1_BUFX2_526 ( );
FILL FILL_0_BUFX2_461 ( );
FILL FILL_1_BUFX2_461 ( );
FILL FILL_0_DFFPOSX1_432 ( );
FILL FILL_1_DFFPOSX1_432 ( );
FILL FILL_2_DFFPOSX1_432 ( );
FILL FILL_3_DFFPOSX1_432 ( );
FILL FILL_4_DFFPOSX1_432 ( );
FILL FILL_5_DFFPOSX1_432 ( );
FILL FILL_6_DFFPOSX1_432 ( );
FILL FILL_0_NAND2X1_160 ( );
FILL FILL_0_OAI21X1_419 ( );
FILL FILL_1_OAI21X1_419 ( );
FILL FILL_0_BUFX2_456 ( );
FILL FILL_0_BUFX2_313 ( );
FILL FILL_0_NAND2X1_397 ( );
FILL FILL_1_NAND2X1_397 ( );
FILL FILL_0_NAND2X1_154 ( );
FILL FILL_0_BUFX2_520 ( );
FILL FILL_1_BUFX2_520 ( );
FILL FILL_0_BUFX2_647 ( );
FILL FILL_1_BUFX2_647 ( );
FILL FILL_0_BUFX2_128 ( );
FILL FILL_1_BUFX2_128 ( );
FILL FILL_0_BUFX2_648 ( );
FILL FILL_1_BUFX2_648 ( );
FILL FILL_0_BUFX2_506 ( );
FILL FILL_0_BUFX2_463 ( );
FILL FILL_1_BUFX2_463 ( );
FILL FILL_0_NAND2X1_344 ( );
FILL FILL_0_DFFPOSX1_434 ( );
FILL FILL_1_DFFPOSX1_434 ( );
FILL FILL_2_DFFPOSX1_434 ( );
FILL FILL_3_DFFPOSX1_434 ( );
FILL FILL_4_DFFPOSX1_434 ( );
FILL FILL_5_DFFPOSX1_434 ( );
FILL FILL_6_DFFPOSX1_434 ( );
FILL FILL_0_BUFX2_284 ( );
FILL FILL_1_BUFX2_284 ( );
FILL FILL_0_BUFX2_548 ( );
FILL FILL_1_BUFX2_548 ( );
FILL FILL_0_BUFX2_346 ( );
FILL FILL_1_BUFX2_346 ( );
FILL FILL_0_NAND2X1_341 ( );
FILL FILL_1_NAND2X1_341 ( );
FILL FILL_0_BUFX2_917 ( );
FILL FILL_0_OAI21X1_847 ( );
FILL FILL_1_OAI21X1_847 ( );
FILL FILL_0_BUFX2_789 ( );
FILL FILL_0_INVX1_48 ( );
FILL FILL_0_BUFX2_1023 ( );
FILL FILL_0_BUFX2_289 ( );
FILL FILL_1_BUFX2_289 ( );
FILL FILL_0_DFFPOSX1_619 ( );
FILL FILL_1_DFFPOSX1_619 ( );
FILL FILL_2_DFFPOSX1_619 ( );
FILL FILL_3_DFFPOSX1_619 ( );
FILL FILL_4_DFFPOSX1_619 ( );
FILL FILL_5_DFFPOSX1_619 ( );
FILL FILL_0_BUFX2_673 ( );
FILL FILL_1_BUFX2_673 ( );
FILL FILL_0_BUFX2_556 ( );
FILL FILL_1_BUFX2_556 ( );
FILL FILL_0_BUFX2_360 ( );
FILL FILL_0_BUFX2_769 ( );
FILL FILL_1_BUFX2_769 ( );
FILL FILL_0_BUFX2_505 ( );
FILL FILL_1_BUFX2_505 ( );
FILL FILL_0_BUFX2_421 ( );
FILL FILL_1_BUFX2_421 ( );
FILL FILL_0_BUFX2_625 ( );
FILL FILL_0_BUFX2_422 ( );
FILL FILL_1_BUFX2_422 ( );
FILL FILL_0_BUFX2_451 ( );
FILL FILL_0_BUFX2_645 ( );
FILL FILL_1_BUFX2_645 ( );
FILL FILL_0_BUFX2_484 ( );
FILL FILL_1_BUFX2_484 ( );
FILL FILL_0_BUFX2_853 ( );
FILL FILL_1_BUFX2_853 ( );
FILL FILL_0_BUFX2_409 ( );
FILL FILL_1_BUFX2_409 ( );
FILL FILL_0_BUFX2_407 ( );
FILL FILL_0_BUFX2_854 ( );
FILL FILL_0_BUFX2_483 ( );
FILL FILL_1_BUFX2_483 ( );
FILL FILL_0_BUFX2_472 ( );
FILL FILL_0_BUFX2_981 ( );
FILL FILL_1_BUFX2_981 ( );
FILL FILL_0_BUFX2_473 ( );
FILL FILL_1_BUFX2_473 ( );
FILL FILL_0_BUFX2_601 ( );
FILL FILL_1_BUFX2_601 ( );
FILL FILL_0_BUFX2_537 ( );
FILL FILL_0_BUFX2_992 ( );
FILL FILL_0_BUFX2_692 ( );
FILL FILL_1_BUFX2_692 ( );
FILL FILL_0_BUFX2_535 ( );
FILL FILL_1_BUFX2_535 ( );
FILL FILL_0_DFFPOSX1_23 ( );
FILL FILL_1_DFFPOSX1_23 ( );
FILL FILL_2_DFFPOSX1_23 ( );
FILL FILL_3_DFFPOSX1_23 ( );
FILL FILL_4_DFFPOSX1_23 ( );
FILL FILL_5_DFFPOSX1_23 ( );
FILL FILL_0_BUFX2_478 ( );
FILL FILL_1_BUFX2_478 ( );
FILL FILL_0_BUFX2_831 ( );
FILL FILL_0_BUFX2_470 ( );
FILL FILL_1_BUFX2_470 ( );
FILL FILL_0_BUFX2_538 ( );
FILL FILL_1_BUFX2_538 ( );
FILL FILL_0_BUFX2_408 ( );
FILL FILL_1_BUFX2_408 ( );
FILL FILL_0_BUFX2_476 ( );
FILL FILL_1_BUFX2_476 ( );
FILL FILL_0_BUFX2_790 ( );
FILL FILL_1_BUFX2_790 ( );
FILL FILL_0_BUFX2_414 ( );
FILL FILL_1_BUFX2_414 ( );
FILL FILL_0_BUFX2_825 ( );
FILL FILL_1_BUFX2_825 ( );
FILL FILL_0_DFFPOSX1_152 ( );
FILL FILL_1_DFFPOSX1_152 ( );
FILL FILL_2_DFFPOSX1_152 ( );
FILL FILL_3_DFFPOSX1_152 ( );
FILL FILL_4_DFFPOSX1_152 ( );
FILL FILL_5_DFFPOSX1_152 ( );
FILL FILL_6_DFFPOSX1_152 ( );
FILL FILL_0_INVX2_198 ( );
FILL FILL_0_BUFX2_895 ( );
FILL FILL_1_BUFX2_895 ( );
FILL FILL_0_NAND2X1_66 ( );
FILL FILL_1_NAND2X1_66 ( );
FILL FILL_0_INVX2_144 ( );
FILL FILL_0_BUFX2_418 ( );
FILL FILL_1_BUFX2_418 ( );
FILL FILL_0_NAND2X1_48 ( );
FILL FILL_1_NAND2X1_48 ( );
FILL FILL_0_NAND2X1_60 ( );
FILL FILL_1_NAND2X1_60 ( );
FILL FILL_0_NAND2X1_709 ( );
FILL FILL_1_NAND2X1_709 ( );
FILL FILL_0_BUFX2_889 ( );
FILL FILL_1_BUFX2_889 ( );
FILL FILL_0_BUFX2_701 ( );
FILL FILL_0_BUFX2_940 ( );
FILL FILL_0_BUFX2_876 ( );
FILL FILL_1_BUFX2_876 ( );
FILL FILL_0_BUFX2_334 ( );
FILL FILL_0_BUFX2_206 ( );
FILL FILL_1_BUFX2_206 ( );
FILL FILL_0_BUFX2_942 ( );
FILL FILL_1_BUFX2_942 ( );
FILL FILL_0_BUFX2_959 ( );
FILL FILL_1_BUFX2_959 ( );
FILL FILL_0_BUFX2_341 ( );
FILL FILL_1_BUFX2_341 ( );
FILL FILL_0_BUFX2_14 ( );
FILL FILL_0_INVX1_87 ( );
FILL FILL_0_BUFX2_898 ( );
FILL FILL_0_BUFX2_295 ( );
FILL FILL_0_DFFPOSX1_678 ( );
FILL FILL_1_DFFPOSX1_678 ( );
FILL FILL_2_DFFPOSX1_678 ( );
FILL FILL_3_DFFPOSX1_678 ( );
FILL FILL_4_DFFPOSX1_678 ( );
FILL FILL_5_DFFPOSX1_678 ( );
FILL FILL_0_BUFX2_80 ( );
FILL FILL_1_BUFX2_80 ( );
FILL FILL_0_BUFX2_81 ( );
FILL FILL_1_BUFX2_81 ( );
FILL FILL_0_BUFX2_698 ( );
FILL FILL_0_BUFX2_834 ( );
FILL FILL_1_BUFX2_834 ( );
FILL FILL_0_BUFX2_317 ( );
FILL FILL_1_BUFX2_317 ( );
FILL FILL_0_NAND2X1_389 ( );
FILL FILL_0_OAI21X1_895 ( );
FILL FILL_1_OAI21X1_895 ( );
FILL FILL_0_INVX1_96 ( );
FILL FILL_0_BUFX2_896 ( );
FILL FILL_0_BUFX2_1024 ( );
FILL FILL_1_BUFX2_1024 ( );
FILL FILL_0_BUFX2_304 ( );
FILL FILL_1_BUFX2_304 ( );
FILL FILL_0_BUFX2_970 ( );
FILL FILL_1_BUFX2_970 ( );
FILL FILL_0_BUFX2_843 ( );
FILL FILL_1_BUFX2_843 ( );
FILL FILL_0_BUFX2_666 ( );
FILL FILL_1_BUFX2_666 ( );
FILL FILL_0_BUFX2_842 ( );
FILL FILL_1_BUFX2_842 ( );
FILL FILL_0_BUFX2_832 ( );
FILL FILL_1_BUFX2_832 ( );
FILL FILL_0_BUFX2_718 ( );
FILL FILL_1_BUFX2_718 ( );
FILL FILL_0_BUFX2_686 ( );
FILL FILL_1_BUFX2_686 ( );
FILL FILL_0_BUFX2_162 ( );
FILL FILL_1_BUFX2_162 ( );
FILL FILL_0_BUFX2_95 ( );
FILL FILL_0_BUFX2_384 ( );
FILL FILL_0_BUFX2_37 ( );
FILL FILL_1_BUFX2_37 ( );
FILL FILL_0_INVX1_146 ( );
FILL FILL_0_BUFX2_799 ( );
FILL FILL_1_BUFX2_799 ( );
FILL FILL_0_BUFX2_94 ( );
FILL FILL_1_BUFX2_94 ( );
FILL FILL_0_BUFX2_314 ( );
FILL FILL_1_BUFX2_314 ( );
FILL FILL_0_BUFX2_814 ( );
FILL FILL_1_BUFX2_814 ( );
FILL FILL_0_BUFX2_33 ( );
FILL FILL_0_BUFX2_221 ( );
FILL FILL_1_BUFX2_221 ( );
FILL FILL_0_BUFX2_225 ( );
FILL FILL_0_BUFX2_30 ( );
FILL FILL_0_INVX1_106 ( );
FILL FILL_0_BUFX2_36 ( );
FILL FILL_1_BUFX2_36 ( );
FILL FILL_0_BUFX2_165 ( );
FILL FILL_0_BUFX2_98 ( );
FILL FILL_0_BUFX2_315 ( );
FILL FILL_1_BUFX2_315 ( );
FILL FILL_0_DFFPOSX1_618 ( );
FILL FILL_1_DFFPOSX1_618 ( );
FILL FILL_2_DFFPOSX1_618 ( );
FILL FILL_3_DFFPOSX1_618 ( );
FILL FILL_4_DFFPOSX1_618 ( );
FILL FILL_5_DFFPOSX1_618 ( );
FILL FILL_6_DFFPOSX1_618 ( );
FILL FILL_0_OAI21X1_846 ( );
FILL FILL_1_OAI21X1_846 ( );
FILL FILL_0_INVX1_47 ( );
FILL FILL_0_NAND2X1_340 ( );
FILL FILL_1_NAND2X1_340 ( );
FILL FILL_0_BUFX2_368 ( );
FILL FILL_0_BUFX2_307 ( );
FILL FILL_1_BUFX2_307 ( );
FILL FILL_0_BUFX2_273 ( );
FILL FILL_1_BUFX2_273 ( );
FILL FILL_0_DFFPOSX1_719 ( );
FILL FILL_1_DFFPOSX1_719 ( );
FILL FILL_2_DFFPOSX1_719 ( );
FILL FILL_3_DFFPOSX1_719 ( );
FILL FILL_4_DFFPOSX1_719 ( );
FILL FILL_5_DFFPOSX1_719 ( );
FILL FILL_0_BUFX2_370 ( );
FILL FILL_1_BUFX2_370 ( );
FILL FILL_0_BUFX2_363 ( );
FILL FILL_0_BUFX2_386 ( );
FILL FILL_0_BUFX2_112 ( );
FILL FILL_1_BUFX2_112 ( );
FILL FILL_0_INVX1_72 ( );
FILL FILL_0_OAI21X1_871 ( );
FILL FILL_1_OAI21X1_871 ( );
FILL FILL_0_DFFPOSX1_643 ( );
FILL FILL_1_DFFPOSX1_643 ( );
FILL FILL_2_DFFPOSX1_643 ( );
FILL FILL_3_DFFPOSX1_643 ( );
FILL FILL_4_DFFPOSX1_643 ( );
FILL FILL_5_DFFPOSX1_643 ( );
FILL FILL_0_NAND2X1_350 ( );
FILL FILL_0_BUFX2_990 ( );
FILL FILL_1_BUFX2_990 ( );
FILL FILL_0_NAND2X1_365 ( );
FILL FILL_1_NAND2X1_365 ( );
FILL FILL_0_BUFX2_822 ( );
FILL FILL_1_BUFX2_822 ( );
FILL FILL_0_BUFX2_778 ( );
FILL FILL_1_BUFX2_778 ( );
FILL FILL_0_BUFX2_281 ( );
FILL FILL_1_BUFX2_281 ( );
FILL FILL_0_BUFX2_54 ( );
FILL FILL_1_BUFX2_54 ( );
FILL FILL_0_BUFX2_265 ( );
FILL FILL_1_BUFX2_265 ( );
FILL FILL_0_NAND2X1_363 ( );
FILL FILL_0_BUFX2_311 ( );
FILL FILL_0_BUFX2_279 ( );
FILL FILL_1_BUFX2_279 ( );
FILL FILL_0_NAND2X1_338 ( );
FILL FILL_1_NAND2X1_338 ( );
FILL FILL_0_OAI21X1_844 ( );
FILL FILL_1_OAI21X1_844 ( );
FILL FILL_0_INVX1_45 ( );
FILL FILL_0_DFFPOSX1_616 ( );
FILL FILL_1_DFFPOSX1_616 ( );
FILL FILL_2_DFFPOSX1_616 ( );
FILL FILL_3_DFFPOSX1_616 ( );
FILL FILL_4_DFFPOSX1_616 ( );
FILL FILL_5_DFFPOSX1_616 ( );
FILL FILL_6_DFFPOSX1_616 ( );
FILL FILL_0_OAI21X1_863 ( );
FILL FILL_1_OAI21X1_863 ( );
FILL FILL_0_BUFX2_300 ( );
FILL FILL_0_BUFX2_276 ( );
FILL FILL_1_BUFX2_276 ( );
FILL FILL_0_INVX1_64 ( );
FILL FILL_1_INVX1_64 ( );
FILL FILL_0_NAND2X1_357 ( );
FILL FILL_0_BUFX2_261 ( );
FILL FILL_0_BUFX2_272 ( );
FILL FILL_0_BUFX2_290 ( );
FILL FILL_0_BUFX2_376 ( );
FILL FILL_0_NAND2X1_360 ( );
FILL FILL_1_NAND2X1_360 ( );
FILL FILL_0_INVX1_88 ( );
FILL FILL_0_BUFX2_296 ( );
FILL FILL_1_BUFX2_296 ( );
FILL FILL_0_OAI21X1_887 ( );
FILL FILL_1_OAI21X1_887 ( );
FILL FILL_2_OAI21X1_887 ( );
FILL FILL_0_NAND2X1_381 ( );
FILL FILL_0_DFFPOSX1_659 ( );
FILL FILL_1_DFFPOSX1_659 ( );
FILL FILL_2_DFFPOSX1_659 ( );
FILL FILL_3_DFFPOSX1_659 ( );
FILL FILL_4_DFFPOSX1_659 ( );
FILL FILL_5_DFFPOSX1_659 ( );
FILL FILL_6_DFFPOSX1_659 ( );
FILL FILL_0_INVX1_122 ( );
FILL FILL_0_OAI21X1_875 ( );
FILL FILL_1_OAI21X1_875 ( );
FILL FILL_0_INVX1_76 ( );
FILL FILL_0_DFFPOSX1_647 ( );
FILL FILL_1_DFFPOSX1_647 ( );
FILL FILL_2_DFFPOSX1_647 ( );
FILL FILL_3_DFFPOSX1_647 ( );
FILL FILL_4_DFFPOSX1_647 ( );
FILL FILL_5_DFFPOSX1_647 ( );
FILL FILL_0_OAI21X1_854 ( );
FILL FILL_1_OAI21X1_854 ( );
FILL FILL_0_INVX1_136 ( );
FILL FILL_0_INVX2_154 ( );
FILL FILL_0_INVX1_55 ( );
FILL FILL_0_DFFPOSX1_626 ( );
FILL FILL_1_DFFPOSX1_626 ( );
FILL FILL_2_DFFPOSX1_626 ( );
FILL FILL_3_DFFPOSX1_626 ( );
FILL FILL_4_DFFPOSX1_626 ( );
FILL FILL_5_DFFPOSX1_626 ( );
FILL FILL_0_INVX1_100 ( );
FILL FILL_0_BUFX4_232 ( );
FILL FILL_1_BUFX4_232 ( );
FILL FILL_0_OAI21X1_899 ( );
FILL FILL_1_OAI21X1_899 ( );
FILL FILL_0_NAND2X1_393 ( );
FILL FILL_1_NAND2X1_393 ( );
FILL FILL_0_DFFPOSX1_671 ( );
FILL FILL_1_DFFPOSX1_671 ( );
FILL FILL_2_DFFPOSX1_671 ( );
FILL FILL_3_DFFPOSX1_671 ( );
FILL FILL_4_DFFPOSX1_671 ( );
FILL FILL_5_DFFPOSX1_671 ( );
FILL FILL_0_BUFX2_438 ( );
FILL FILL_0_OAI21X1_859 ( );
FILL FILL_1_OAI21X1_859 ( );
FILL FILL_0_INVX1_60 ( );
FILL FILL_0_DFFPOSX1_631 ( );
FILL FILL_1_DFFPOSX1_631 ( );
FILL FILL_2_DFFPOSX1_631 ( );
FILL FILL_3_DFFPOSX1_631 ( );
FILL FILL_4_DFFPOSX1_631 ( );
FILL FILL_5_DFFPOSX1_631 ( );
FILL FILL_6_DFFPOSX1_631 ( );
FILL FILL_0_BUFX2_513 ( );
FILL FILL_1_BUFX2_513 ( );
FILL FILL_0_BUFX2_458 ( );
FILL FILL_1_BUFX2_458 ( );
FILL FILL_0_BUFX2_491 ( );
FILL FILL_1_BUFX2_491 ( );
FILL FILL_0_INVX1_94 ( );
FILL FILL_0_BUFX4_262 ( );
FILL FILL_1_BUFX4_262 ( );
FILL FILL_0_OAI21X1_893 ( );
FILL FILL_1_OAI21X1_893 ( );
FILL FILL_0_NAND2X1_387 ( );
FILL FILL_1_NAND2X1_387 ( );
FILL FILL_0_DFFPOSX1_665 ( );
FILL FILL_1_DFFPOSX1_665 ( );
FILL FILL_2_DFFPOSX1_665 ( );
FILL FILL_3_DFFPOSX1_665 ( );
FILL FILL_4_DFFPOSX1_665 ( );
FILL FILL_5_DFFPOSX1_665 ( );
FILL FILL_0_OAI21X1_1644 ( );
FILL FILL_1_OAI21X1_1644 ( );
FILL FILL_2_OAI21X1_1644 ( );
FILL FILL_0_NAND2X1_712 ( );
FILL FILL_0_DFFPOSX1_34 ( );
FILL FILL_1_DFFPOSX1_34 ( );
FILL FILL_2_DFFPOSX1_34 ( );
FILL FILL_3_DFFPOSX1_34 ( );
FILL FILL_4_DFFPOSX1_34 ( );
FILL FILL_5_DFFPOSX1_34 ( );
FILL FILL_0_DFFPOSX1_433 ( );
FILL FILL_1_DFFPOSX1_433 ( );
FILL FILL_2_DFFPOSX1_433 ( );
FILL FILL_3_DFFPOSX1_433 ( );
FILL FILL_4_DFFPOSX1_433 ( );
FILL FILL_5_DFFPOSX1_433 ( );
FILL FILL_0_OAI21X1_420 ( );
FILL FILL_1_OAI21X1_420 ( );
FILL FILL_2_OAI21X1_420 ( );
FILL FILL_0_NAND2X1_161 ( );
FILL FILL_0_BUFX2_459 ( );
FILL FILL_0_BUFX2_436 ( );
FILL FILL_0_INVX1_104 ( );
FILL FILL_0_OAI21X1_903 ( );
FILL FILL_1_OAI21X1_903 ( );
FILL FILL_0_DFFPOSX1_675 ( );
FILL FILL_1_DFFPOSX1_675 ( );
FILL FILL_2_DFFPOSX1_675 ( );
FILL FILL_3_DFFPOSX1_675 ( );
FILL FILL_4_DFFPOSX1_675 ( );
FILL FILL_5_DFFPOSX1_675 ( );
FILL FILL_0_OAI21X1_412 ( );
FILL FILL_1_OAI21X1_412 ( );
FILL FILL_2_OAI21X1_412 ( );
FILL FILL_0_DFFPOSX1_429 ( );
FILL FILL_1_DFFPOSX1_429 ( );
FILL FILL_2_DFFPOSX1_429 ( );
FILL FILL_3_DFFPOSX1_429 ( );
FILL FILL_4_DFFPOSX1_429 ( );
FILL FILL_5_DFFPOSX1_429 ( );
FILL FILL_6_DFFPOSX1_429 ( );
FILL FILL_0_OAI21X1_421 ( );
FILL FILL_1_OAI21X1_421 ( );
FILL FILL_0_NAND2X1_163 ( );
FILL FILL_1_NAND2X1_163 ( );
FILL FILL_0_DFFPOSX1_365 ( );
FILL FILL_1_DFFPOSX1_365 ( );
FILL FILL_2_DFFPOSX1_365 ( );
FILL FILL_3_DFFPOSX1_365 ( );
FILL FILL_4_DFFPOSX1_365 ( );
FILL FILL_5_DFFPOSX1_365 ( );
FILL FILL_0_BUFX2_499 ( );
FILL FILL_1_BUFX2_499 ( );
FILL FILL_0_BUFX2_455 ( );
FILL FILL_1_BUFX2_455 ( );
FILL FILL_0_BUFX2_402 ( );
FILL FILL_0_BUFX2_629 ( );
FILL FILL_1_BUFX2_629 ( );
FILL FILL_0_BUFX2_444 ( );
FILL FILL_1_BUFX2_444 ( );
FILL FILL_0_INVX2_115 ( );
FILL FILL_0_INVX1_137 ( );
FILL FILL_0_OAI21X1_965 ( );
FILL FILL_1_OAI21X1_965 ( );
FILL FILL_0_DFFPOSX1_708 ( );
FILL FILL_1_DFFPOSX1_708 ( );
FILL FILL_2_DFFPOSX1_708 ( );
FILL FILL_3_DFFPOSX1_708 ( );
FILL FILL_4_DFFPOSX1_708 ( );
FILL FILL_5_DFFPOSX1_708 ( );
FILL FILL_0_OAI21X1_850 ( );
FILL FILL_1_OAI21X1_850 ( );
FILL FILL_0_INVX1_51 ( );
FILL FILL_1_INVX1_51 ( );
FILL FILL_0_OAI21X1_1611 ( );
FILL FILL_1_OAI21X1_1611 ( );
FILL FILL_0_NAND2X1_680 ( );
FILL FILL_0_INVX2_2 ( );
FILL FILL_0_DFFPOSX1_2 ( );
FILL FILL_1_DFFPOSX1_2 ( );
FILL FILL_2_DFFPOSX1_2 ( );
FILL FILL_3_DFFPOSX1_2 ( );
FILL FILL_4_DFFPOSX1_2 ( );
FILL FILL_5_DFFPOSX1_2 ( );
FILL FILL_0_INVX1_152 ( );
FILL FILL_0_INVX2_166 ( );
FILL FILL_0_DFFPOSX1_166 ( );
FILL FILL_1_DFFPOSX1_166 ( );
FILL FILL_2_DFFPOSX1_166 ( );
FILL FILL_3_DFFPOSX1_166 ( );
FILL FILL_4_DFFPOSX1_166 ( );
FILL FILL_5_DFFPOSX1_166 ( );
FILL FILL_0_NAND2X1_10 ( );
FILL FILL_1_NAND2X1_10 ( );
FILL FILL_0_DFFPOSX1_443 ( );
FILL FILL_1_DFFPOSX1_443 ( );
FILL FILL_2_DFFPOSX1_443 ( );
FILL FILL_3_DFFPOSX1_443 ( );
FILL FILL_4_DFFPOSX1_443 ( );
FILL FILL_5_DFFPOSX1_443 ( );
FILL FILL_0_OAI21X1_1633 ( );
FILL FILL_1_OAI21X1_1633 ( );
FILL FILL_0_NAND2X1_701 ( );
FILL FILL_0_OAI21X1_28 ( );
FILL FILL_1_OAI21X1_28 ( );
FILL FILL_2_OAI21X1_28 ( );
FILL FILL_0_NAND2X1_28 ( );
FILL FILL_0_DFFPOSX1_184 ( );
FILL FILL_1_DFFPOSX1_184 ( );
FILL FILL_2_DFFPOSX1_184 ( );
FILL FILL_3_DFFPOSX1_184 ( );
FILL FILL_4_DFFPOSX1_184 ( );
FILL FILL_5_DFFPOSX1_184 ( );
FILL FILL_0_BUFX2_406 ( );
FILL FILL_1_BUFX2_406 ( );
FILL FILL_0_OAI21X1_1794 ( );
FILL FILL_1_OAI21X1_1794 ( );
FILL FILL_0_NAND2X1_735 ( );
FILL FILL_1_NAND2X1_735 ( );
FILL FILL_0_DFFPOSX1_120 ( );
FILL FILL_1_DFFPOSX1_120 ( );
FILL FILL_2_DFFPOSX1_120 ( );
FILL FILL_3_DFFPOSX1_120 ( );
FILL FILL_4_DFFPOSX1_120 ( );
FILL FILL_5_DFFPOSX1_120 ( );
FILL FILL_6_DFFPOSX1_120 ( );
FILL FILL_0_NAND2X1_2 ( );
FILL FILL_1_NAND2X1_2 ( );
FILL FILL_0_DFFPOSX1_222 ( );
FILL FILL_1_DFFPOSX1_222 ( );
FILL FILL_2_DFFPOSX1_222 ( );
FILL FILL_3_DFFPOSX1_222 ( );
FILL FILL_4_DFFPOSX1_222 ( );
FILL FILL_5_DFFPOSX1_222 ( );
FILL FILL_0_OAI21X1_66 ( );
FILL FILL_1_OAI21X1_66 ( );
FILL FILL_0_DFFPOSX1_216 ( );
FILL FILL_1_DFFPOSX1_216 ( );
FILL FILL_2_DFFPOSX1_216 ( );
FILL FILL_3_DFFPOSX1_216 ( );
FILL FILL_4_DFFPOSX1_216 ( );
FILL FILL_5_DFFPOSX1_216 ( );
FILL FILL_0_NAND2X1_767 ( );
FILL FILL_1_NAND2X1_767 ( );
FILL FILL_0_INVX2_186 ( );
FILL FILL_0_OAI21X1_60 ( );
FILL FILL_1_OAI21X1_60 ( );
FILL FILL_0_OAI21X1_1826 ( );
FILL FILL_1_OAI21X1_1826 ( );
FILL FILL_0_DFFPOSX1_204 ( );
FILL FILL_1_DFFPOSX1_204 ( );
FILL FILL_2_DFFPOSX1_204 ( );
FILL FILL_3_DFFPOSX1_204 ( );
FILL FILL_4_DFFPOSX1_204 ( );
FILL FILL_5_DFFPOSX1_204 ( );
FILL FILL_6_DFFPOSX1_204 ( );
FILL FILL_0_BUFX2_357 ( );
FILL FILL_1_BUFX2_357 ( );
FILL FILL_0_OAI21X1_48 ( );
FILL FILL_1_OAI21X1_48 ( );
FILL FILL_0_OAI21X1_955 ( );
FILL FILL_1_OAI21X1_955 ( );
FILL FILL_0_INVX1_132 ( );
FILL FILL_0_DFFPOSX1_703 ( );
FILL FILL_1_DFFPOSX1_703 ( );
FILL FILL_2_DFFPOSX1_703 ( );
FILL FILL_3_DFFPOSX1_703 ( );
FILL FILL_4_DFFPOSX1_703 ( );
FILL FILL_5_DFFPOSX1_703 ( );
FILL FILL_0_INVX1_126 ( );
FILL FILL_0_BUFX2_76 ( );
FILL FILL_1_BUFX2_76 ( );
FILL FILL_0_NAND2X1_380 ( );
FILL FILL_1_NAND2X1_380 ( );
FILL FILL_0_OAI21X1_886 ( );
FILL FILL_1_OAI21X1_886 ( );
FILL FILL_0_INVX2_141 ( );
FILL FILL_0_INVX1_118 ( );
FILL FILL_0_OAI21X1_927 ( );
FILL FILL_1_OAI21X1_927 ( );
FILL FILL_0_BUFX2_356 ( );
FILL FILL_1_BUFX2_356 ( );
FILL FILL_0_INVX1_107 ( );
FILL FILL_0_OAI21X1_906 ( );
FILL FILL_1_OAI21X1_906 ( );
FILL FILL_0_NAND2X1_400 ( );
FILL FILL_1_NAND2X1_400 ( );
FILL FILL_0_DFFPOSX1_223 ( );
FILL FILL_1_DFFPOSX1_223 ( );
FILL FILL_2_DFFPOSX1_223 ( );
FILL FILL_3_DFFPOSX1_223 ( );
FILL FILL_4_DFFPOSX1_223 ( );
FILL FILL_5_DFFPOSX1_223 ( );
FILL FILL_0_DFFPOSX1_667 ( );
FILL FILL_1_DFFPOSX1_667 ( );
FILL FILL_2_DFFPOSX1_667 ( );
FILL FILL_3_DFFPOSX1_667 ( );
FILL FILL_4_DFFPOSX1_667 ( );
FILL FILL_5_DFFPOSX1_667 ( );
FILL FILL_0_INVX2_120 ( );
FILL FILL_0_OAI21X1_67 ( );
FILL FILL_1_OAI21X1_67 ( );
FILL FILL_2_OAI21X1_67 ( );
FILL FILL_0_NAND2X1_67 ( );
FILL FILL_0_BUFX2_391 ( );
FILL FILL_0_DFFPOSX1_129 ( );
FILL FILL_1_DFFPOSX1_129 ( );
FILL FILL_2_DFFPOSX1_129 ( );
FILL FILL_3_DFFPOSX1_129 ( );
FILL FILL_4_DFFPOSX1_129 ( );
FILL FILL_5_DFFPOSX1_129 ( );
FILL FILL_0_DFFPOSX1_844 ( );
FILL FILL_1_DFFPOSX1_844 ( );
FILL FILL_2_DFFPOSX1_844 ( );
FILL FILL_3_DFFPOSX1_844 ( );
FILL FILL_4_DFFPOSX1_844 ( );
FILL FILL_5_DFFPOSX1_844 ( );
FILL FILL_0_NAND2X1_537 ( );
FILL FILL_0_INVX2_3 ( );
FILL FILL_0_DFFPOSX1_847 ( );
FILL FILL_1_DFFPOSX1_847 ( );
FILL FILL_2_DFFPOSX1_847 ( );
FILL FILL_3_DFFPOSX1_847 ( );
FILL FILL_4_DFFPOSX1_847 ( );
FILL FILL_5_DFFPOSX1_847 ( );
FILL FILL_0_BUFX2_97 ( );
FILL FILL_1_BUFX2_97 ( );
FILL FILL_0_INVX2_188 ( );
FILL FILL_0_NAND2X1_398 ( );
FILL FILL_1_NAND2X1_398 ( );
FILL FILL_0_OAI21X1_904 ( );
FILL FILL_1_OAI21X1_904 ( );
FILL FILL_0_INVX1_105 ( );
FILL FILL_0_DFFPOSX1_677 ( );
FILL FILL_1_DFFPOSX1_677 ( );
FILL FILL_2_DFFPOSX1_677 ( );
FILL FILL_3_DFFPOSX1_677 ( );
FILL FILL_4_DFFPOSX1_677 ( );
FILL FILL_5_DFFPOSX1_677 ( );
FILL FILL_0_NAND2X1_399 ( );
FILL FILL_1_NAND2X1_399 ( );
FILL FILL_0_OAI21X1_905 ( );
FILL FILL_1_OAI21X1_905 ( );
FILL FILL_0_INVX2_175 ( );
FILL FILL_0_BUFX2_158 ( );
FILL FILL_1_BUFX2_158 ( );
FILL FILL_0_INVX1_98 ( );
FILL FILL_0_OAI21X1_897 ( );
FILL FILL_1_OAI21X1_897 ( );
FILL FILL_0_NAND2X1_391 ( );
FILL FILL_1_NAND2X1_391 ( );
FILL FILL_0_DFFPOSX1_726 ( );
FILL FILL_1_DFFPOSX1_726 ( );
FILL FILL_2_DFFPOSX1_726 ( );
FILL FILL_3_DFFPOSX1_726 ( );
FILL FILL_4_DFFPOSX1_726 ( );
FILL FILL_5_DFFPOSX1_726 ( );
FILL FILL_6_DFFPOSX1_726 ( );
FILL FILL_0_OAI21X1_1001 ( );
FILL FILL_1_OAI21X1_1001 ( );
FILL FILL_2_OAI21X1_1001 ( );
FILL FILL_0_INVX1_155 ( );
FILL FILL_0_BUFX4_261 ( );
FILL FILL_1_BUFX4_261 ( );
FILL FILL_2_BUFX4_261 ( );
FILL FILL_0_BUFX4_264 ( );
FILL FILL_1_BUFX4_264 ( );
FILL FILL_0_DFFPOSX1_628 ( );
FILL FILL_1_DFFPOSX1_628 ( );
FILL FILL_2_DFFPOSX1_628 ( );
FILL FILL_3_DFFPOSX1_628 ( );
FILL FILL_4_DFFPOSX1_628 ( );
FILL FILL_5_DFFPOSX1_628 ( );
FILL FILL_0_BUFX2_798 ( );
FILL FILL_1_BUFX2_798 ( );
FILL FILL_0_INVX1_161 ( );
FILL FILL_0_BUFX2_1014 ( );
FILL FILL_1_BUFX2_1014 ( );
FILL FILL_0_OAI21X1_856 ( );
FILL FILL_1_OAI21X1_856 ( );
FILL FILL_0_INVX1_57 ( );
FILL FILL_0_OAI21X1_987 ( );
FILL FILL_1_OAI21X1_987 ( );
FILL FILL_0_INVX1_148 ( );
FILL FILL_0_DFFPOSX1_641 ( );
FILL FILL_1_DFFPOSX1_641 ( );
FILL FILL_2_DFFPOSX1_641 ( );
FILL FILL_3_DFFPOSX1_641 ( );
FILL FILL_4_DFFPOSX1_641 ( );
FILL FILL_5_DFFPOSX1_641 ( );
FILL FILL_0_INVX1_70 ( );
FILL FILL_0_OAI21X1_869 ( );
FILL FILL_1_OAI21X1_869 ( );
FILL FILL_0_DFFPOSX1_673 ( );
FILL FILL_1_DFFPOSX1_673 ( );
FILL FILL_2_DFFPOSX1_673 ( );
FILL FILL_3_DFFPOSX1_673 ( );
FILL FILL_4_DFFPOSX1_673 ( );
FILL FILL_5_DFFPOSX1_673 ( );
FILL FILL_0_NAND2X1_395 ( );
FILL FILL_0_OAI21X1_901 ( );
FILL FILL_1_OAI21X1_901 ( );
FILL FILL_0_INVX2_174 ( );
FILL FILL_0_INVX1_102 ( );
FILL FILL_0_DFFPOSX1_663 ( );
FILL FILL_1_DFFPOSX1_663 ( );
FILL FILL_2_DFFPOSX1_663 ( );
FILL FILL_3_DFFPOSX1_663 ( );
FILL FILL_4_DFFPOSX1_663 ( );
FILL FILL_5_DFFPOSX1_663 ( );
FILL FILL_6_DFFPOSX1_663 ( );
FILL FILL_0_DFFPOSX1_635 ( );
FILL FILL_1_DFFPOSX1_635 ( );
FILL FILL_2_DFFPOSX1_635 ( );
FILL FILL_3_DFFPOSX1_635 ( );
FILL FILL_4_DFFPOSX1_635 ( );
FILL FILL_5_DFFPOSX1_635 ( );
FILL FILL_6_DFFPOSX1_635 ( );
FILL FILL_0_INVX2_7 ( );
FILL FILL_0_NAND2X1_385 ( );
FILL FILL_1_NAND2X1_385 ( );
FILL FILL_0_OAI21X1_891 ( );
FILL FILL_1_OAI21X1_891 ( );
FILL FILL_0_INVX1_92 ( );
FILL FILL_0_DFFPOSX1_638 ( );
FILL FILL_1_DFFPOSX1_638 ( );
FILL FILL_2_DFFPOSX1_638 ( );
FILL FILL_3_DFFPOSX1_638 ( );
FILL FILL_4_DFFPOSX1_638 ( );
FILL FILL_5_DFFPOSX1_638 ( );
FILL FILL_0_INVX1_67 ( );
FILL FILL_0_OAI21X1_866 ( );
FILL FILL_1_OAI21X1_866 ( );
FILL FILL_0_DFFPOSX1_629 ( );
FILL FILL_1_DFFPOSX1_629 ( );
FILL FILL_2_DFFPOSX1_629 ( );
FILL FILL_3_DFFPOSX1_629 ( );
FILL FILL_4_DFFPOSX1_629 ( );
FILL FILL_5_DFFPOSX1_629 ( );
FILL FILL_6_DFFPOSX1_629 ( );
FILL FILL_0_INVX1_58 ( );
FILL FILL_0_OAI21X1_857 ( );
FILL FILL_1_OAI21X1_857 ( );
FILL FILL_0_INVX1_167 ( );
FILL FILL_0_BUFX2_949 ( );
FILL FILL_1_BUFX2_949 ( );
FILL FILL_0_INVX2_187 ( );
FILL FILL_0_BUFX2_285 ( );
FILL FILL_0_NAND2X1_339 ( );
FILL FILL_1_NAND2X1_339 ( );
FILL FILL_0_OAI21X1_874 ( );
FILL FILL_1_OAI21X1_874 ( );
FILL FILL_2_OAI21X1_874 ( );
FILL FILL_0_INVX1_75 ( );
FILL FILL_0_BUFX2_344 ( );
FILL FILL_1_BUFX2_344 ( );
FILL FILL_0_BUFX2_330 ( );
FILL FILL_1_BUFX2_330 ( );
FILL FILL_0_OAI21X1_934 ( );
FILL FILL_1_OAI21X1_934 ( );
FILL FILL_0_OAI21X1_935 ( );
FILL FILL_1_OAI21X1_935 ( );
FILL FILL_0_DFFPOSX1_693 ( );
FILL FILL_1_DFFPOSX1_693 ( );
FILL FILL_2_DFFPOSX1_693 ( );
FILL FILL_3_DFFPOSX1_693 ( );
FILL FILL_4_DFFPOSX1_693 ( );
FILL FILL_5_DFFPOSX1_693 ( );
FILL FILL_0_BUFX4_268 ( );
FILL FILL_1_BUFX4_268 ( );
FILL FILL_0_DFFPOSX1_707 ( );
FILL FILL_1_DFFPOSX1_707 ( );
FILL FILL_2_DFFPOSX1_707 ( );
FILL FILL_3_DFFPOSX1_707 ( );
FILL FILL_4_DFFPOSX1_707 ( );
FILL FILL_5_DFFPOSX1_707 ( );
FILL FILL_6_DFFPOSX1_707 ( );
FILL FILL_0_OAI21X1_963 ( );
FILL FILL_1_OAI21X1_963 ( );
FILL FILL_0_OAI21X1_962 ( );
FILL FILL_1_OAI21X1_962 ( );
FILL FILL_0_BUFX2_903 ( );
FILL FILL_1_BUFX2_903 ( );
FILL FILL_0_BUFX2_345 ( );
FILL FILL_0_OAI21X1_16 ( );
FILL FILL_1_OAI21X1_16 ( );
FILL FILL_0_NAND2X1_16 ( );
FILL FILL_0_DFFPOSX1_172 ( );
FILL FILL_1_DFFPOSX1_172 ( );
FILL FILL_2_DFFPOSX1_172 ( );
FILL FILL_3_DFFPOSX1_172 ( );
FILL FILL_4_DFFPOSX1_172 ( );
FILL FILL_5_DFFPOSX1_172 ( );
FILL FILL_6_DFFPOSX1_172 ( );
FILL FILL_0_BUFX2_457 ( );
FILL FILL_1_BUFX2_457 ( );
FILL FILL_0_NAND2X1_136 ( );
FILL FILL_0_OAI21X1_392 ( );
FILL FILL_1_OAI21X1_392 ( );
FILL FILL_0_BUFX4_237 ( );
FILL FILL_1_BUFX4_237 ( );
FILL FILL_0_DFFPOSX1_420 ( );
FILL FILL_1_DFFPOSX1_420 ( );
FILL FILL_2_DFFPOSX1_420 ( );
FILL FILL_3_DFFPOSX1_420 ( );
FILL FILL_4_DFFPOSX1_420 ( );
FILL FILL_5_DFFPOSX1_420 ( );
FILL FILL_0_NAND2X1_148 ( );
FILL FILL_1_NAND2X1_148 ( );
FILL FILL_0_BUFX2_401 ( );
FILL FILL_1_BUFX2_401 ( );
FILL FILL_0_BUFX2_518 ( );
FILL FILL_1_BUFX2_518 ( );
FILL FILL_0_DFFPOSX1_427 ( );
FILL FILL_1_DFFPOSX1_427 ( );
FILL FILL_2_DFFPOSX1_427 ( );
FILL FILL_3_DFFPOSX1_427 ( );
FILL FILL_4_DFFPOSX1_427 ( );
FILL FILL_5_DFFPOSX1_427 ( );
FILL FILL_6_DFFPOSX1_427 ( );
FILL FILL_0_OAI21X1_409 ( );
FILL FILL_1_OAI21X1_409 ( );
FILL FILL_0_NAND2X1_152 ( );
FILL FILL_0_BUFX2_497 ( );
FILL FILL_1_BUFX2_497 ( );
FILL FILL_0_NAND2X1_227 ( );
FILL FILL_0_BUFX2_737 ( );
FILL FILL_0_BUFX2_460 ( );
FILL FILL_1_BUFX2_460 ( );
FILL FILL_0_DFFPOSX1_431 ( );
FILL FILL_1_DFFPOSX1_431 ( );
FILL FILL_2_DFFPOSX1_431 ( );
FILL FILL_3_DFFPOSX1_431 ( );
FILL FILL_4_DFFPOSX1_431 ( );
FILL FILL_5_DFFPOSX1_431 ( );
FILL FILL_0_NAND2X1_158 ( );
FILL FILL_0_OAI21X1_416 ( );
FILL FILL_1_OAI21X1_416 ( );
FILL FILL_2_OAI21X1_416 ( );
FILL FILL_0_BUFX4_225 ( );
FILL FILL_1_BUFX4_225 ( );
FILL FILL_0_BUFX2_587 ( );
FILL FILL_1_BUFX2_587 ( );
FILL FILL_0_DFFPOSX1_430 ( );
FILL FILL_1_DFFPOSX1_430 ( );
FILL FILL_2_DFFPOSX1_430 ( );
FILL FILL_3_DFFPOSX1_430 ( );
FILL FILL_4_DFFPOSX1_430 ( );
FILL FILL_5_DFFPOSX1_430 ( );
FILL FILL_0_NAND2X1_156 ( );
FILL FILL_0_OAI21X1_415 ( );
FILL FILL_1_OAI21X1_415 ( );
FILL FILL_0_NAND2X1_153 ( );
FILL FILL_1_NAND2X1_153 ( );
FILL FILL_0_XNOR2X1_1 ( );
FILL FILL_1_XNOR2X1_1 ( );
FILL FILL_2_XNOR2X1_1 ( );
FILL FILL_3_XNOR2X1_1 ( );
FILL FILL_0_BUFX2_498 ( );
FILL FILL_0_NAND2X1_164 ( );
FILL FILL_1_NAND2X1_164 ( );
FILL FILL_0_BUFX2_867 ( );
FILL FILL_0_BUFX4_215 ( );
FILL FILL_1_BUFX4_215 ( );
FILL FILL_2_BUFX4_215 ( );
FILL FILL_0_NAND2X1_40 ( );
FILL FILL_1_NAND2X1_40 ( );
FILL FILL_0_BUFX2_399 ( );
FILL FILL_0_BUFX2_443 ( );
FILL FILL_0_BUFX2_586 ( );
FILL FILL_0_OAI21X1_337 ( );
FILL FILL_1_OAI21X1_337 ( );
FILL FILL_0_NAND2X1_81 ( );
FILL FILL_1_NAND2X1_81 ( );
FILL FILL_0_DFFPOSX1_364 ( );
FILL FILL_1_DFFPOSX1_364 ( );
FILL FILL_2_DFFPOSX1_364 ( );
FILL FILL_3_DFFPOSX1_364 ( );
FILL FILL_4_DFFPOSX1_364 ( );
FILL FILL_5_DFFPOSX1_364 ( );
FILL FILL_6_DFFPOSX1_364 ( );
FILL FILL_0_BUFX2_514 ( );
FILL FILL_0_INVX2_148 ( );
FILL FILL_0_BUFX2_466 ( );
FILL FILL_1_BUFX2_466 ( );
FILL FILL_0_BUFX2_486 ( );
FILL FILL_1_BUFX2_486 ( );
FILL FILL_0_OAI21X1_964 ( );
FILL FILL_1_OAI21X1_964 ( );
FILL FILL_2_OAI21X1_964 ( );
FILL FILL_0_BUFX2_485 ( );
FILL FILL_0_BUFX2_612 ( );
FILL FILL_0_DFFPOSX1_622 ( );
FILL FILL_1_DFFPOSX1_622 ( );
FILL FILL_2_DFFPOSX1_622 ( );
FILL FILL_3_DFFPOSX1_622 ( );
FILL FILL_4_DFFPOSX1_622 ( );
FILL FILL_5_DFFPOSX1_622 ( );
FILL FILL_6_DFFPOSX1_622 ( );
FILL FILL_0_DFFPOSX1_230 ( );
FILL FILL_1_DFFPOSX1_230 ( );
FILL FILL_2_DFFPOSX1_230 ( );
FILL FILL_3_DFFPOSX1_230 ( );
FILL FILL_4_DFFPOSX1_230 ( );
FILL FILL_5_DFFPOSX1_230 ( );
FILL FILL_6_DFFPOSX1_230 ( );
FILL FILL_0_BUFX2_617 ( );
FILL FILL_1_BUFX2_617 ( );
FILL FILL_0_NAND2X1_717 ( );
FILL FILL_1_NAND2X1_717 ( );
FILL FILL_0_DFFPOSX1_294 ( );
FILL FILL_1_DFFPOSX1_294 ( );
FILL FILL_2_DFFPOSX1_294 ( );
FILL FILL_3_DFFPOSX1_294 ( );
FILL FILL_4_DFFPOSX1_294 ( );
FILL FILL_5_DFFPOSX1_294 ( );
FILL FILL_0_OAI21X1_10 ( );
FILL FILL_1_OAI21X1_10 ( );
FILL FILL_0_BUFX2_471 ( );
FILL FILL_1_BUFX2_471 ( );
FILL FILL_0_BUFX4_233 ( );
FILL FILL_1_BUFX4_233 ( );
FILL FILL_0_NAND2X1_184 ( );
FILL FILL_1_NAND2X1_184 ( );
FILL FILL_0_DFFPOSX1_377 ( );
FILL FILL_1_DFFPOSX1_377 ( );
FILL FILL_2_DFFPOSX1_377 ( );
FILL FILL_3_DFFPOSX1_377 ( );
FILL FILL_4_DFFPOSX1_377 ( );
FILL FILL_5_DFFPOSX1_377 ( );
FILL FILL_6_DFFPOSX1_377 ( );
FILL FILL_0_NAND2X1_95 ( );
FILL FILL_1_NAND2X1_95 ( );
FILL FILL_0_NAND2X1_93 ( );
FILL FILL_1_NAND2X1_93 ( );
FILL FILL_0_OAI21X1_349 ( );
FILL FILL_1_OAI21X1_349 ( );
FILL FILL_0_INVX1_149 ( );
FILL FILL_0_BUFX2_1017 ( );
FILL FILL_1_BUFX2_1017 ( );
FILL FILL_0_DFFPOSX1_376 ( );
FILL FILL_1_DFFPOSX1_376 ( );
FILL FILL_2_DFFPOSX1_376 ( );
FILL FILL_3_DFFPOSX1_376 ( );
FILL FILL_4_DFFPOSX1_376 ( );
FILL FILL_5_DFFPOSX1_376 ( );
FILL FILL_0_DFFPOSX1_158 ( );
FILL FILL_1_DFFPOSX1_158 ( );
FILL FILL_2_DFFPOSX1_158 ( );
FILL FILL_3_DFFPOSX1_158 ( );
FILL FILL_4_DFFPOSX1_158 ( );
FILL FILL_5_DFFPOSX1_158 ( );
FILL FILL_0_OAI21X1_2 ( );
FILL FILL_1_OAI21X1_2 ( );
FILL FILL_0_BUFX2_387 ( );
FILL FILL_1_BUFX2_387 ( );
FILL FILL_0_DFFPOSX1_384 ( );
FILL FILL_1_DFFPOSX1_384 ( );
FILL FILL_2_DFFPOSX1_384 ( );
FILL FILL_3_DFFPOSX1_384 ( );
FILL FILL_4_DFFPOSX1_384 ( );
FILL FILL_5_DFFPOSX1_384 ( );
FILL FILL_6_DFFPOSX1_384 ( );
FILL FILL_0_BUFX4_190 ( );
FILL FILL_1_BUFX4_190 ( );
FILL FILL_0_BUFX2_372 ( );
FILL FILL_1_BUFX2_372 ( );
FILL FILL_0_DFFPOSX1_31 ( );
FILL FILL_1_DFFPOSX1_31 ( );
FILL FILL_2_DFFPOSX1_31 ( );
FILL FILL_3_DFFPOSX1_31 ( );
FILL FILL_4_DFFPOSX1_31 ( );
FILL FILL_5_DFFPOSX1_31 ( );
FILL FILL_6_DFFPOSX1_31 ( );
FILL FILL_0_OAI21X1_1641 ( );
FILL FILL_1_OAI21X1_1641 ( );
FILL FILL_0_DFFPOSX1_712 ( );
FILL FILL_1_DFFPOSX1_712 ( );
FILL FILL_2_DFFPOSX1_712 ( );
FILL FILL_3_DFFPOSX1_712 ( );
FILL FILL_4_DFFPOSX1_712 ( );
FILL FILL_5_DFFPOSX1_712 ( );
FILL FILL_0_OAI21X1_156 ( );
FILL FILL_1_OAI21X1_156 ( );
FILL FILL_0_OAI21X1_157 ( );
FILL FILL_1_OAI21X1_157 ( );
FILL FILL_0_OAI21X1_954 ( );
FILL FILL_1_OAI21X1_954 ( );
FILL FILL_2_OAI21X1_954 ( );
FILL FILL_0_BUFX2_667 ( );
FILL FILL_0_BUFX2_18 ( );
FILL FILL_1_BUFX2_18 ( );
FILL FILL_0_OAI21X1_942 ( );
FILL FILL_1_OAI21X1_942 ( );
FILL FILL_0_OAI21X1_943 ( );
FILL FILL_1_OAI21X1_943 ( );
FILL FILL_0_BUFX2_144 ( );
FILL FILL_0_DFFPOSX1_658 ( );
FILL FILL_1_DFFPOSX1_658 ( );
FILL FILL_2_DFFPOSX1_658 ( );
FILL FILL_3_DFFPOSX1_658 ( );
FILL FILL_4_DFFPOSX1_658 ( );
FILL FILL_5_DFFPOSX1_658 ( );
FILL FILL_0_INVX2_4 ( );
FILL FILL_0_NAND2X1_4 ( );
FILL FILL_1_NAND2X1_4 ( );
FILL FILL_0_OAI21X1_926 ( );
FILL FILL_1_OAI21X1_926 ( );
FILL FILL_0_DFFPOSX1_689 ( );
FILL FILL_1_DFFPOSX1_689 ( );
FILL FILL_2_DFFPOSX1_689 ( );
FILL FILL_3_DFFPOSX1_689 ( );
FILL FILL_4_DFFPOSX1_689 ( );
FILL FILL_5_DFFPOSX1_689 ( );
FILL FILL_6_DFFPOSX1_689 ( );
FILL FILL_0_BUFX2_79 ( );
FILL FILL_0_DFFPOSX1_206 ( );
FILL FILL_1_DFFPOSX1_206 ( );
FILL FILL_2_DFFPOSX1_206 ( );
FILL FILL_3_DFFPOSX1_206 ( );
FILL FILL_4_DFFPOSX1_206 ( );
FILL FILL_5_DFFPOSX1_206 ( );
FILL FILL_6_DFFPOSX1_206 ( );
FILL FILL_0_BUFX2_878 ( );
FILL FILL_0_BUFX2_207 ( );
FILL FILL_0_OAI21X1_1605 ( );
FILL FILL_1_OAI21X1_1605 ( );
FILL FILL_0_NAND2X1_18 ( );
FILL FILL_1_NAND2X1_18 ( );
FILL FILL_0_NAND2X1_674 ( );
FILL FILL_1_NAND2X1_674 ( );
FILL FILL_0_DFFPOSX1_1028 ( );
FILL FILL_1_DFFPOSX1_1028 ( );
FILL FILL_2_DFFPOSX1_1028 ( );
FILL FILL_3_DFFPOSX1_1028 ( );
FILL FILL_4_DFFPOSX1_1028 ( );
FILL FILL_5_DFFPOSX1_1028 ( );
FILL FILL_0_DFFPOSX1_165 ( );
FILL FILL_1_DFFPOSX1_165 ( );
FILL FILL_2_DFFPOSX1_165 ( );
FILL FILL_3_DFFPOSX1_165 ( );
FILL FILL_4_DFFPOSX1_165 ( );
FILL FILL_5_DFFPOSX1_165 ( );
FILL FILL_6_DFFPOSX1_165 ( );
FILL FILL_0_BUFX2_392 ( );
FILL FILL_1_BUFX2_392 ( );
FILL FILL_0_OAI21X1_1160 ( );
FILL FILL_1_OAI21X1_1160 ( );
FILL FILL_0_BUFX2_371 ( );
FILL FILL_0_OAI21X1_1803 ( );
FILL FILL_1_OAI21X1_1803 ( );
FILL FILL_0_NAND2X1_744 ( );
FILL FILL_1_NAND2X1_744 ( );
FILL FILL_0_DFFPOSX1_843 ( );
FILL FILL_1_DFFPOSX1_843 ( );
FILL FILL_2_DFFPOSX1_843 ( );
FILL FILL_3_DFFPOSX1_843 ( );
FILL FILL_4_DFFPOSX1_843 ( );
FILL FILL_5_DFFPOSX1_843 ( );
FILL FILL_6_DFFPOSX1_843 ( );
FILL FILL_0_NAND2X1_544 ( );
FILL FILL_1_NAND2X1_544 ( );
FILL FILL_0_OAI21X1_1816 ( );
FILL FILL_1_OAI21X1_1816 ( );
FILL FILL_0_DFFPOSX1_142 ( );
FILL FILL_1_DFFPOSX1_142 ( );
FILL FILL_2_DFFPOSX1_142 ( );
FILL FILL_3_DFFPOSX1_142 ( );
FILL FILL_4_DFFPOSX1_142 ( );
FILL FILL_5_DFFPOSX1_142 ( );
FILL FILL_0_DFFPOSX1_676 ( );
FILL FILL_1_DFFPOSX1_676 ( );
FILL FILL_2_DFFPOSX1_676 ( );
FILL FILL_3_DFFPOSX1_676 ( );
FILL FILL_4_DFFPOSX1_676 ( );
FILL FILL_5_DFFPOSX1_676 ( );
FILL FILL_6_DFFPOSX1_676 ( );
FILL FILL_0_DFFPOSX1_971 ( );
FILL FILL_1_DFFPOSX1_971 ( );
FILL FILL_2_DFFPOSX1_971 ( );
FILL FILL_3_DFFPOSX1_971 ( );
FILL FILL_4_DFFPOSX1_971 ( );
FILL FILL_5_DFFPOSX1_971 ( );
FILL FILL_6_DFFPOSX1_971 ( );
FILL FILL_0_BUFX2_222 ( );
FILL FILL_0_OAI21X1_1000 ( );
FILL FILL_1_OAI21X1_1000 ( );
FILL FILL_0_DFFPOSX1_669 ( );
FILL FILL_1_DFFPOSX1_669 ( );
FILL FILL_2_DFFPOSX1_669 ( );
FILL FILL_3_DFFPOSX1_669 ( );
FILL FILL_4_DFFPOSX1_669 ( );
FILL FILL_5_DFFPOSX1_669 ( );
FILL FILL_0_BUFX2_239 ( );
FILL FILL_1_BUFX2_239 ( );
FILL FILL_0_BUFX2_102 ( );
FILL FILL_1_BUFX2_102 ( );
FILL FILL_0_BUFX2_228 ( );
FILL FILL_0_DFFPOSX1_128 ( );
FILL FILL_1_DFFPOSX1_128 ( );
FILL FILL_2_DFFPOSX1_128 ( );
FILL FILL_3_DFFPOSX1_128 ( );
FILL FILL_4_DFFPOSX1_128 ( );
FILL FILL_5_DFFPOSX1_128 ( );
FILL FILL_6_DFFPOSX1_128 ( );
FILL FILL_0_NAND2X1_743 ( );
FILL FILL_1_NAND2X1_743 ( );
FILL FILL_0_OAI21X1_1802 ( );
FILL FILL_1_OAI21X1_1802 ( );
FILL FILL_0_OAI21X1_986 ( );
FILL FILL_1_OAI21X1_986 ( );
FILL FILL_0_OAI21X1_256 ( );
FILL FILL_1_OAI21X1_256 ( );
FILL FILL_0_OAI21X1_257 ( );
FILL FILL_1_OAI21X1_257 ( );
FILL FILL_0_DFFPOSX1_320 ( );
FILL FILL_1_DFFPOSX1_320 ( );
FILL FILL_2_DFFPOSX1_320 ( );
FILL FILL_3_DFFPOSX1_320 ( );
FILL FILL_4_DFFPOSX1_320 ( );
FILL FILL_5_DFFPOSX1_320 ( );
FILL FILL_0_NAND2X1_716 ( );
FILL FILL_1_NAND2X1_716 ( );
FILL FILL_0_CLKBUF1_82 ( );
FILL FILL_1_CLKBUF1_82 ( );
FILL FILL_2_CLKBUF1_82 ( );
FILL FILL_3_CLKBUF1_82 ( );
FILL FILL_0_BUFX2_926 ( );
FILL FILL_1_BUFX2_926 ( );
FILL FILL_0_OAI21X1_36 ( );
FILL FILL_1_OAI21X1_36 ( );
FILL FILL_0_NAND2X1_36 ( );
FILL FILL_1_NAND2X1_36 ( );
FILL FILL_0_DFFPOSX1_192 ( );
FILL FILL_1_DFFPOSX1_192 ( );
FILL FILL_2_DFFPOSX1_192 ( );
FILL FILL_3_DFFPOSX1_192 ( );
FILL FILL_4_DFFPOSX1_192 ( );
FILL FILL_5_DFFPOSX1_192 ( );
FILL FILL_0_BUFX2_886 ( );
FILL FILL_1_BUFX2_886 ( );
FILL FILL_0_BUFX2_862 ( );
FILL FILL_0_OAI21X1_71 ( );
FILL FILL_1_OAI21X1_71 ( );
FILL FILL_2_OAI21X1_71 ( );
FILL FILL_0_NAND2X1_71 ( );
FILL FILL_0_DFFPOSX1_227 ( );
FILL FILL_1_DFFPOSX1_227 ( );
FILL FILL_2_DFFPOSX1_227 ( );
FILL FILL_3_DFFPOSX1_227 ( );
FILL FILL_4_DFFPOSX1_227 ( );
FILL FILL_5_DFFPOSX1_227 ( );
FILL FILL_0_BUFX2_901 ( );
FILL FILL_0_BUFX2_1029 ( );
FILL FILL_1_BUFX2_1029 ( );
FILL FILL_0_BUFX2_352 ( );
FILL FILL_0_DFFPOSX1_623 ( );
FILL FILL_1_DFFPOSX1_623 ( );
FILL FILL_2_DFFPOSX1_623 ( );
FILL FILL_3_DFFPOSX1_623 ( );
FILL FILL_4_DFFPOSX1_623 ( );
FILL FILL_5_DFFPOSX1_623 ( );
FILL FILL_0_INVX1_52 ( );
FILL FILL_0_OAI21X1_851 ( );
FILL FILL_1_OAI21X1_851 ( );
FILL FILL_0_DFFPOSX1_653 ( );
FILL FILL_1_DFFPOSX1_653 ( );
FILL FILL_2_DFFPOSX1_653 ( );
FILL FILL_3_DFFPOSX1_653 ( );
FILL FILL_4_DFFPOSX1_653 ( );
FILL FILL_5_DFFPOSX1_653 ( );
FILL FILL_6_DFFPOSX1_653 ( );
FILL FILL_0_INVX2_122 ( );
FILL FILL_0_INVX1_95 ( );
FILL FILL_0_BUFX2_347 ( );
FILL FILL_0_INVX2_116 ( );
FILL FILL_1_INVX2_116 ( );
FILL FILL_0_INVX1_168 ( );
FILL FILL_0_INVX1_138 ( );
FILL FILL_0_DFFPOSX1_646 ( );
FILL FILL_1_DFFPOSX1_646 ( );
FILL FILL_2_DFFPOSX1_646 ( );
FILL FILL_3_DFFPOSX1_646 ( );
FILL FILL_4_DFFPOSX1_646 ( );
FILL FILL_5_DFFPOSX1_646 ( );
FILL FILL_6_DFFPOSX1_646 ( );
FILL FILL_0_INVX1_135 ( );
FILL FILL_0_OAI21X1_961 ( );
FILL FILL_1_OAI21X1_961 ( );
FILL FILL_0_OAI21X1_960 ( );
FILL FILL_1_OAI21X1_960 ( );
FILL FILL_0_DFFPOSX1_706 ( );
FILL FILL_1_DFFPOSX1_706 ( );
FILL FILL_2_DFFPOSX1_706 ( );
FILL FILL_3_DFFPOSX1_706 ( );
FILL FILL_4_DFFPOSX1_706 ( );
FILL FILL_5_DFFPOSX1_706 ( );
FILL FILL_0_INVX2_178 ( );
FILL FILL_0_BUFX2_910 ( );
FILL FILL_1_BUFX2_910 ( );
FILL FILL_0_INVX2_159 ( );
FILL FILL_0_INVX2_149 ( );
FILL FILL_0_OAI21X1_98 ( );
FILL FILL_1_OAI21X1_98 ( );
FILL FILL_0_OAI21X1_99 ( );
FILL FILL_1_OAI21X1_99 ( );
FILL FILL_0_BUFX2_770 ( );
FILL FILL_1_BUFX2_770 ( );
FILL FILL_0_DFFPOSX1_241 ( );
FILL FILL_1_DFFPOSX1_241 ( );
FILL FILL_2_DFFPOSX1_241 ( );
FILL FILL_3_DFFPOSX1_241 ( );
FILL FILL_4_DFFPOSX1_241 ( );
FILL FILL_5_DFFPOSX1_241 ( );
FILL FILL_6_DFFPOSX1_241 ( );
FILL FILL_0_OAI21X1_21 ( );
FILL FILL_1_OAI21X1_21 ( );
FILL FILL_0_NAND2X1_21 ( );
FILL FILL_1_NAND2X1_21 ( );
FILL FILL_0_DFFPOSX1_177 ( );
FILL FILL_1_DFFPOSX1_177 ( );
FILL FILL_2_DFFPOSX1_177 ( );
FILL FILL_3_DFFPOSX1_177 ( );
FILL FILL_4_DFFPOSX1_177 ( );
FILL FILL_5_DFFPOSX1_177 ( );
FILL FILL_0_BUFX2_555 ( );
FILL FILL_0_BUFX2_974 ( );
FILL FILL_0_BUFX2_641 ( );
FILL FILL_0_CLKBUF1_10 ( );
FILL FILL_1_CLKBUF1_10 ( );
FILL FILL_2_CLKBUF1_10 ( );
FILL FILL_3_CLKBUF1_10 ( );
FILL FILL_0_DFFPOSX1_426 ( );
FILL FILL_1_DFFPOSX1_426 ( );
FILL FILL_2_DFFPOSX1_426 ( );
FILL FILL_3_DFFPOSX1_426 ( );
FILL FILL_4_DFFPOSX1_426 ( );
FILL FILL_5_DFFPOSX1_426 ( );
FILL FILL_0_NAND2X1_144 ( );
FILL FILL_0_DFFPOSX1_424 ( );
FILL FILL_1_DFFPOSX1_424 ( );
FILL FILL_2_DFFPOSX1_424 ( );
FILL FILL_3_DFFPOSX1_424 ( );
FILL FILL_4_DFFPOSX1_424 ( );
FILL FILL_5_DFFPOSX1_424 ( );
FILL FILL_0_DFFPOSX1_465 ( );
FILL FILL_1_DFFPOSX1_465 ( );
FILL FILL_2_DFFPOSX1_465 ( );
FILL FILL_3_DFFPOSX1_465 ( );
FILL FILL_4_DFFPOSX1_465 ( );
FILL FILL_5_DFFPOSX1_465 ( );
FILL FILL_0_DFFPOSX1_366 ( );
FILL FILL_1_DFFPOSX1_366 ( );
FILL FILL_2_DFFPOSX1_366 ( );
FILL FILL_3_DFFPOSX1_366 ( );
FILL FILL_4_DFFPOSX1_366 ( );
FILL FILL_5_DFFPOSX1_366 ( );
FILL FILL_0_NAND2X1_82 ( );
FILL FILL_1_NAND2X1_82 ( );
FILL FILL_0_OAI21X1_338 ( );
FILL FILL_1_OAI21X1_338 ( );
FILL FILL_0_BUFX2_589 ( );
FILL FILL_0_INVX2_15 ( );
FILL FILL_0_BUFX2_562 ( );
FILL FILL_1_BUFX2_562 ( );
FILL FILL_0_XNOR2X1_3 ( );
FILL FILL_1_XNOR2X1_3 ( );
FILL FILL_2_XNOR2X1_3 ( );
FILL FILL_3_XNOR2X1_3 ( );
FILL FILL_0_INVX4_3 ( );
FILL FILL_0_DFFPOSX1_428 ( );
FILL FILL_1_DFFPOSX1_428 ( );
FILL FILL_2_DFFPOSX1_428 ( );
FILL FILL_3_DFFPOSX1_428 ( );
FILL FILL_4_DFFPOSX1_428 ( );
FILL FILL_5_DFFPOSX1_428 ( );
FILL FILL_0_OAI21X1_411 ( );
FILL FILL_1_OAI21X1_411 ( );
FILL FILL_0_BUFX4_181 ( );
FILL FILL_1_BUFX4_181 ( );
FILL FILL_0_OAI21X1_422 ( );
FILL FILL_1_OAI21X1_422 ( );
FILL FILL_0_DFFPOSX1_435 ( );
FILL FILL_1_DFFPOSX1_435 ( );
FILL FILL_2_DFFPOSX1_435 ( );
FILL FILL_3_DFFPOSX1_435 ( );
FILL FILL_4_DFFPOSX1_435 ( );
FILL FILL_5_DFFPOSX1_435 ( );
FILL FILL_0_OAI21X1_40 ( );
FILL FILL_1_OAI21X1_40 ( );
FILL FILL_0_NAND2X1_83 ( );
FILL FILL_0_BUFX2_396 ( );
FILL FILL_1_BUFX2_396 ( );
FILL FILL_0_DFFPOSX1_196 ( );
FILL FILL_1_DFFPOSX1_196 ( );
FILL FILL_2_DFFPOSX1_196 ( );
FILL FILL_3_DFFPOSX1_196 ( );
FILL FILL_4_DFFPOSX1_196 ( );
FILL FILL_5_DFFPOSX1_196 ( );
FILL FILL_0_OAI21X1_336 ( );
FILL FILL_1_OAI21X1_336 ( );
FILL FILL_0_NAND2X1_80 ( );
FILL FILL_1_NAND2X1_80 ( );
FILL FILL_0_NAND2X1_89 ( );
FILL FILL_1_NAND2X1_89 ( );
FILL FILL_0_OAI21X1_342 ( );
FILL FILL_1_OAI21X1_342 ( );
FILL FILL_0_NAND2X1_86 ( );
FILL FILL_0_DFFPOSX1_370 ( );
FILL FILL_1_DFFPOSX1_370 ( );
FILL FILL_2_DFFPOSX1_370 ( );
FILL FILL_3_DFFPOSX1_370 ( );
FILL FILL_4_DFFPOSX1_370 ( );
FILL FILL_5_DFFPOSX1_370 ( );
FILL FILL_0_BUFX2_549 ( );
FILL FILL_1_BUFX2_549 ( );
FILL FILL_0_DFFPOSX1_98 ( );
FILL FILL_1_DFFPOSX1_98 ( );
FILL FILL_2_DFFPOSX1_98 ( );
FILL FILL_3_DFFPOSX1_98 ( );
FILL FILL_4_DFFPOSX1_98 ( );
FILL FILL_5_DFFPOSX1_98 ( );
FILL FILL_6_DFFPOSX1_98 ( );
FILL FILL_0_OAI21X1_77 ( );
FILL FILL_1_OAI21X1_77 ( );
FILL FILL_2_OAI21X1_77 ( );
FILL FILL_0_OAI21X1_76 ( );
FILL FILL_1_OAI21X1_76 ( );
FILL FILL_0_BUFX2_642 ( );
FILL FILL_1_BUFX2_642 ( );
FILL FILL_0_OAI21X1_1776 ( );
FILL FILL_1_OAI21X1_1776 ( );
FILL FILL_0_DFFPOSX1_102 ( );
FILL FILL_1_DFFPOSX1_102 ( );
FILL FILL_2_DFFPOSX1_102 ( );
FILL FILL_3_DFFPOSX1_102 ( );
FILL FILL_4_DFFPOSX1_102 ( );
FILL FILL_5_DFFPOSX1_102 ( );
FILL FILL_6_DFFPOSX1_102 ( );
FILL FILL_0_OAI21X1_205 ( );
FILL FILL_1_OAI21X1_205 ( );
FILL FILL_0_BUFX2_554 ( );
FILL FILL_1_BUFX2_554 ( );
FILL FILL_0_OAI21X1_995 ( );
FILL FILL_1_OAI21X1_995 ( );
FILL FILL_0_BUFX2_536 ( );
FILL FILL_1_BUFX2_536 ( );
FILL FILL_0_OAI21X1_434 ( );
FILL FILL_1_OAI21X1_434 ( );
FILL FILL_2_OAI21X1_434 ( );
FILL FILL_0_DFFPOSX1_723 ( );
FILL FILL_1_DFFPOSX1_723 ( );
FILL FILL_2_DFFPOSX1_723 ( );
FILL FILL_3_DFFPOSX1_723 ( );
FILL FILL_4_DFFPOSX1_723 ( );
FILL FILL_5_DFFPOSX1_723 ( );
FILL FILL_0_DFFPOSX1_379 ( );
FILL FILL_1_DFFPOSX1_379 ( );
FILL FILL_2_DFFPOSX1_379 ( );
FILL FILL_3_DFFPOSX1_379 ( );
FILL FILL_4_DFFPOSX1_379 ( );
FILL FILL_5_DFFPOSX1_379 ( );
FILL FILL_0_DFFPOSX1_378 ( );
FILL FILL_1_DFFPOSX1_378 ( );
FILL FILL_2_DFFPOSX1_378 ( );
FILL FILL_3_DFFPOSX1_378 ( );
FILL FILL_4_DFFPOSX1_378 ( );
FILL FILL_5_DFFPOSX1_378 ( );
FILL FILL_0_NAND2X1_94 ( );
FILL FILL_1_NAND2X1_94 ( );
FILL FILL_0_NAND2X1_92 ( );
FILL FILL_0_OAI21X1_348 ( );
FILL FILL_1_OAI21X1_348 ( );
FILL FILL_2_OAI21X1_348 ( );
FILL FILL_0_BUFX2_479 ( );
FILL FILL_1_BUFX2_479 ( );
FILL FILL_0_DFFPOSX1_507 ( );
FILL FILL_1_DFFPOSX1_507 ( );
FILL FILL_2_DFFPOSX1_507 ( );
FILL FILL_3_DFFPOSX1_507 ( );
FILL FILL_4_DFFPOSX1_507 ( );
FILL FILL_5_DFFPOSX1_507 ( );
FILL FILL_6_DFFPOSX1_507 ( );
FILL FILL_0_BUFX2_410 ( );
FILL FILL_0_BUFX2_474 ( );
FILL FILL_1_BUFX2_474 ( );
FILL FILL_0_DFFPOSX1_446 ( );
FILL FILL_1_DFFPOSX1_446 ( );
FILL FILL_2_DFFPOSX1_446 ( );
FILL FILL_3_DFFPOSX1_446 ( );
FILL FILL_4_DFFPOSX1_446 ( );
FILL FILL_5_DFFPOSX1_446 ( );
FILL FILL_0_NAND2X1_100 ( );
FILL FILL_0_DFFPOSX1_720 ( );
FILL FILL_1_DFFPOSX1_720 ( );
FILL FILL_2_DFFPOSX1_720 ( );
FILL FILL_3_DFFPOSX1_720 ( );
FILL FILL_4_DFFPOSX1_720 ( );
FILL FILL_5_DFFPOSX1_720 ( );
FILL FILL_6_DFFPOSX1_720 ( );
FILL FILL_0_BUFX2_86 ( );
FILL FILL_1_BUFX2_86 ( );
FILL FILL_0_DFFPOSX1_268 ( );
FILL FILL_1_DFFPOSX1_268 ( );
FILL FILL_2_DFFPOSX1_268 ( );
FILL FILL_3_DFFPOSX1_268 ( );
FILL FILL_4_DFFPOSX1_268 ( );
FILL FILL_5_DFFPOSX1_268 ( );
FILL FILL_0_INVX1_141 ( );
FILL FILL_0_OAI21X1_973 ( );
FILL FILL_1_OAI21X1_973 ( );
FILL FILL_0_INVX1_163 ( );
FILL FILL_0_DFFPOSX1_270 ( );
FILL FILL_1_DFFPOSX1_270 ( );
FILL FILL_2_DFFPOSX1_270 ( );
FILL FILL_3_DFFPOSX1_270 ( );
FILL FILL_4_DFFPOSX1_270 ( );
FILL FILL_5_DFFPOSX1_270 ( );
FILL FILL_0_BUFX2_779 ( );
FILL FILL_0_DFFPOSX1_697 ( );
FILL FILL_1_DFFPOSX1_697 ( );
FILL FILL_2_DFFPOSX1_697 ( );
FILL FILL_3_DFFPOSX1_697 ( );
FILL FILL_4_DFFPOSX1_697 ( );
FILL FILL_5_DFFPOSX1_697 ( );
FILL FILL_0_BUFX2_17 ( );
FILL FILL_0_OAI21X1_4 ( );
FILL FILL_1_OAI21X1_4 ( );
FILL FILL_0_DFFPOSX1_160 ( );
FILL FILL_1_DFFPOSX1_160 ( );
FILL FILL_2_DFFPOSX1_160 ( );
FILL FILL_3_DFFPOSX1_160 ( );
FILL FILL_4_DFFPOSX1_160 ( );
FILL FILL_5_DFFPOSX1_160 ( );
FILL FILL_0_BUFX2_704 ( );
FILL FILL_1_BUFX2_704 ( );
FILL FILL_0_OAI21X1_68 ( );
FILL FILL_1_OAI21X1_68 ( );
FILL FILL_0_NAND2X1_68 ( );
FILL FILL_0_OAI21X1_50 ( );
FILL FILL_1_OAI21X1_50 ( );
FILL FILL_0_NAND2X1_50 ( );
FILL FILL_0_DFFPOSX1_174 ( );
FILL FILL_1_DFFPOSX1_174 ( );
FILL FILL_2_DFFPOSX1_174 ( );
FILL FILL_3_DFFPOSX1_174 ( );
FILL FILL_4_DFFPOSX1_174 ( );
FILL FILL_5_DFFPOSX1_174 ( );
FILL FILL_6_DFFPOSX1_174 ( );
FILL FILL_0_OAI21X1_18 ( );
FILL FILL_1_OAI21X1_18 ( );
FILL FILL_0_BUFX2_145 ( );
FILL FILL_1_BUFX2_145 ( );
FILL FILL_0_BUFX2_16 ( );
FILL FILL_1_BUFX2_16 ( );
FILL FILL_0_INVX2_156 ( );
FILL FILL_0_NAND2X1_9 ( );
FILL FILL_1_NAND2X1_9 ( );
FILL FILL_0_OAI21X1_9 ( );
FILL FILL_1_OAI21X1_9 ( );
FILL FILL_0_DFFPOSX1_717 ( );
FILL FILL_1_DFFPOSX1_717 ( );
FILL FILL_2_DFFPOSX1_717 ( );
FILL FILL_3_DFFPOSX1_717 ( );
FILL FILL_4_DFFPOSX1_717 ( );
FILL FILL_5_DFFPOSX1_717 ( );
FILL FILL_0_BUFX4_185 ( );
FILL FILL_1_BUFX4_185 ( );
FILL FILL_0_DFFPOSX1_779 ( );
FILL FILL_1_DFFPOSX1_779 ( );
FILL FILL_2_DFFPOSX1_779 ( );
FILL FILL_3_DFFPOSX1_779 ( );
FILL FILL_4_DFFPOSX1_779 ( );
FILL FILL_5_DFFPOSX1_779 ( );
FILL FILL_0_OAI21X1_983 ( );
FILL FILL_1_OAI21X1_983 ( );
FILL FILL_0_NAND2X1_437 ( );
FILL FILL_0_OAI21X1_1074 ( );
FILL FILL_1_OAI21X1_1074 ( );
FILL FILL_2_OAI21X1_1074 ( );
FILL FILL_0_NAND2X1_440 ( );
FILL FILL_0_DFFPOSX1_782 ( );
FILL FILL_1_DFFPOSX1_782 ( );
FILL FILL_2_DFFPOSX1_782 ( );
FILL FILL_3_DFFPOSX1_782 ( );
FILL FILL_4_DFFPOSX1_782 ( );
FILL FILL_5_DFFPOSX1_782 ( );
FILL FILL_0_NAND2X1_757 ( );
FILL FILL_1_NAND2X1_757 ( );
FILL FILL_0_BUFX2_34 ( );
FILL FILL_1_BUFX2_34 ( );
FILL FILL_0_BUFX4_189 ( );
FILL FILL_1_BUFX4_189 ( );
FILL FILL_2_BUFX4_189 ( );
FILL FILL_0_CLKBUF1_81 ( );
FILL FILL_1_CLKBUF1_81 ( );
FILL FILL_2_CLKBUF1_81 ( );
FILL FILL_3_CLKBUF1_81 ( );
FILL FILL_4_CLKBUF1_81 ( );
FILL FILL_0_DFFPOSX1_986 ( );
FILL FILL_1_DFFPOSX1_986 ( );
FILL FILL_2_DFFPOSX1_986 ( );
FILL FILL_3_DFFPOSX1_986 ( );
FILL FILL_4_DFFPOSX1_986 ( );
FILL FILL_5_DFFPOSX1_986 ( );
FILL FILL_6_DFFPOSX1_986 ( );
FILL FILL_0_BUFX2_240 ( );
FILL FILL_1_BUFX2_240 ( );
FILL FILL_0_BUFX2_49 ( );
FILL FILL_1_BUFX2_49 ( );
FILL FILL_0_BUFX2_47 ( );
FILL FILL_1_BUFX2_47 ( );
FILL FILL_0_OAI21X1_1011 ( );
FILL FILL_1_OAI21X1_1011 ( );
FILL FILL_2_OAI21X1_1011 ( );
FILL FILL_0_INVX1_160 ( );
FILL FILL_0_OAI21X1_1012 ( );
FILL FILL_1_OAI21X1_1012 ( );
FILL FILL_0_DFFPOSX1_732 ( );
FILL FILL_1_DFFPOSX1_732 ( );
FILL FILL_2_DFFPOSX1_732 ( );
FILL FILL_3_DFFPOSX1_732 ( );
FILL FILL_4_DFFPOSX1_732 ( );
FILL FILL_5_DFFPOSX1_732 ( );
FILL FILL_0_OAI21X1_1013 ( );
FILL FILL_1_OAI21X1_1013 ( );
FILL FILL_0_BUFX2_863 ( );
FILL FILL_1_BUFX2_863 ( );
FILL FILL_0_DFFPOSX1_256 ( );
FILL FILL_1_DFFPOSX1_256 ( );
FILL FILL_2_DFFPOSX1_256 ( );
FILL FILL_3_DFFPOSX1_256 ( );
FILL FILL_4_DFFPOSX1_256 ( );
FILL FILL_5_DFFPOSX1_256 ( );
FILL FILL_6_DFFPOSX1_256 ( );
FILL FILL_0_OAI21X1_129 ( );
FILL FILL_1_OAI21X1_129 ( );
FILL FILL_2_OAI21X1_129 ( );
FILL FILL_0_DFFPOSX1_101 ( );
FILL FILL_1_DFFPOSX1_101 ( );
FILL FILL_2_DFFPOSX1_101 ( );
FILL FILL_3_DFFPOSX1_101 ( );
FILL FILL_4_DFFPOSX1_101 ( );
FILL FILL_5_DFFPOSX1_101 ( );
FILL FILL_0_OAI21X1_1775 ( );
FILL FILL_1_OAI21X1_1775 ( );
FILL FILL_0_CLKBUF1_58 ( );
FILL FILL_1_CLKBUF1_58 ( );
FILL FILL_2_CLKBUF1_58 ( );
FILL FILL_3_CLKBUF1_58 ( );
FILL FILL_4_CLKBUF1_58 ( );
FILL FILL_0_BUFX4_196 ( );
FILL FILL_1_BUFX4_196 ( );
FILL FILL_2_BUFX4_196 ( );
FILL FILL_0_INVX2_147 ( );
FILL FILL_0_BUFX2_243 ( );
FILL FILL_0_INVX2_151 ( );
FILL FILL_0_OAI21X1_13 ( );
FILL FILL_1_OAI21X1_13 ( );
FILL FILL_0_NAND2X1_13 ( );
FILL FILL_1_NAND2X1_13 ( );
FILL FILL_0_OAI21X1_326 ( );
FILL FILL_1_OAI21X1_326 ( );
FILL FILL_0_OAI21X1_327 ( );
FILL FILL_1_OAI21X1_327 ( );
FILL FILL_0_DFFPOSX1_355 ( );
FILL FILL_1_DFFPOSX1_355 ( );
FILL FILL_2_DFFPOSX1_355 ( );
FILL FILL_3_DFFPOSX1_355 ( );
FILL FILL_4_DFFPOSX1_355 ( );
FILL FILL_5_DFFPOSX1_355 ( );
FILL FILL_0_OAI21X1_996 ( );
FILL FILL_1_OAI21X1_996 ( );
FILL FILL_0_OAI21X1_997 ( );
FILL FILL_1_OAI21X1_997 ( );
FILL FILL_0_DFFPOSX1_724 ( );
FILL FILL_1_DFFPOSX1_724 ( );
FILL FILL_2_DFFPOSX1_724 ( );
FILL FILL_3_DFFPOSX1_724 ( );
FILL FILL_4_DFFPOSX1_724 ( );
FILL FILL_5_DFFPOSX1_724 ( );
FILL FILL_6_DFFPOSX1_724 ( );
FILL FILL_0_INVX1_153 ( );
FILL FILL_1_INVX1_153 ( );
FILL FILL_0_DFFPOSX1_666 ( );
FILL FILL_1_DFFPOSX1_666 ( );
FILL FILL_2_DFFPOSX1_666 ( );
FILL FILL_3_DFFPOSX1_666 ( );
FILL FILL_4_DFFPOSX1_666 ( );
FILL FILL_5_DFFPOSX1_666 ( );
FILL FILL_6_DFFPOSX1_666 ( );
FILL FILL_0_NAND2X1_388 ( );
FILL FILL_0_OAI21X1_894 ( );
FILL FILL_1_OAI21X1_894 ( );
FILL FILL_2_OAI21X1_894 ( );
FILL FILL_0_BUFX2_303 ( );
FILL FILL_0_INVX1_134 ( );
FILL FILL_0_INVX1_114 ( );
FILL FILL_1_INVX1_114 ( );
FILL FILL_0_BUFX2_337 ( );
FILL FILL_0_BUFX2_377 ( );
FILL FILL_1_BUFX2_377 ( );
FILL FILL_0_BUFX2_967 ( );
FILL FILL_1_BUFX2_967 ( );
FILL FILL_0_OAI21X1_967 ( );
FILL FILL_1_OAI21X1_967 ( );
FILL FILL_0_OAI21X1_966 ( );
FILL FILL_1_OAI21X1_966 ( );
FILL FILL_0_BUFX2_839 ( );
FILL FILL_0_DFFPOSX1_236 ( );
FILL FILL_1_DFFPOSX1_236 ( );
FILL FILL_2_DFFPOSX1_236 ( );
FILL FILL_3_DFFPOSX1_236 ( );
FILL FILL_4_DFFPOSX1_236 ( );
FILL FILL_5_DFFPOSX1_236 ( );
FILL FILL_0_OAI21X1_88 ( );
FILL FILL_1_OAI21X1_88 ( );
FILL FILL_0_OAI21X1_89 ( );
FILL FILL_1_OAI21X1_89 ( );
FILL FILL_0_NAND2X1_723 ( );
FILL FILL_1_NAND2X1_723 ( );
FILL FILL_0_OAI21X1_1782 ( );
FILL FILL_1_OAI21X1_1782 ( );
FILL FILL_0_BUFX2_803 ( );
FILL FILL_1_BUFX2_803 ( );
FILL FILL_0_CLKBUF1_54 ( );
FILL FILL_1_CLKBUF1_54 ( );
FILL FILL_2_CLKBUF1_54 ( );
FILL FILL_3_CLKBUF1_54 ( );
FILL FILL_4_CLKBUF1_54 ( );
FILL FILL_0_NAND2X1_728 ( );
FILL FILL_1_NAND2X1_728 ( );
FILL FILL_0_BUFX2_782 ( );
FILL FILL_1_BUFX2_782 ( );
FILL FILL_0_BUFX2_674 ( );
FILL FILL_1_BUFX2_674 ( );
FILL FILL_0_DFFPOSX1_3 ( );
FILL FILL_1_DFFPOSX1_3 ( );
FILL FILL_2_DFFPOSX1_3 ( );
FILL FILL_3_DFFPOSX1_3 ( );
FILL FILL_4_DFFPOSX1_3 ( );
FILL FILL_5_DFFPOSX1_3 ( );
FILL FILL_6_DFFPOSX1_3 ( );
FILL FILL_0_NAND2X1_681 ( );
FILL FILL_0_OAI21X1_1612 ( );
FILL FILL_1_OAI21X1_1612 ( );
FILL FILL_0_BUFX2_454 ( );
FILL FILL_0_OAI21X1_227 ( );
FILL FILL_1_OAI21X1_227 ( );
FILL FILL_2_OAI21X1_227 ( );
FILL FILL_0_OAI21X1_226 ( );
FILL FILL_1_OAI21X1_226 ( );
FILL FILL_0_DFFPOSX1_305 ( );
FILL FILL_1_DFFPOSX1_305 ( );
FILL FILL_2_DFFPOSX1_305 ( );
FILL FILL_3_DFFPOSX1_305 ( );
FILL FILL_4_DFFPOSX1_305 ( );
FILL FILL_5_DFFPOSX1_305 ( );
FILL FILL_0_OAI21X1_407 ( );
FILL FILL_1_OAI21X1_407 ( );
FILL FILL_0_INVX1_8 ( );
FILL FILL_0_BUFX4_199 ( );
FILL FILL_1_BUFX4_199 ( );
FILL FILL_0_OAI21X1_401 ( );
FILL FILL_1_OAI21X1_401 ( );
FILL FILL_2_OAI21X1_401 ( );
FILL FILL_0_BUFX2_530 ( );
FILL FILL_1_BUFX2_530 ( );
FILL FILL_0_OAI21X1_467 ( );
FILL FILL_1_OAI21X1_467 ( );
FILL FILL_2_OAI21X1_467 ( );
FILL FILL_0_OAI21X1_1707 ( );
FILL FILL_1_OAI21X1_1707 ( );
FILL FILL_0_OAI21X1_1706 ( );
FILL FILL_1_OAI21X1_1706 ( );
FILL FILL_0_DFFPOSX1_66 ( );
FILL FILL_1_DFFPOSX1_66 ( );
FILL FILL_2_DFFPOSX1_66 ( );
FILL FILL_3_DFFPOSX1_66 ( );
FILL FILL_4_DFFPOSX1_66 ( );
FILL FILL_5_DFFPOSX1_66 ( );
FILL FILL_0_CLKBUF1_13 ( );
FILL FILL_1_CLKBUF1_13 ( );
FILL FILL_2_CLKBUF1_13 ( );
FILL FILL_3_CLKBUF1_13 ( );
FILL FILL_4_CLKBUF1_13 ( );
FILL FILL_0_NAND2X1_87 ( );
FILL FILL_1_NAND2X1_87 ( );
FILL FILL_0_OAI21X1_527 ( );
FILL FILL_1_OAI21X1_527 ( );
FILL FILL_2_OAI21X1_527 ( );
FILL FILL_0_OAI21X1_413 ( );
FILL FILL_1_OAI21X1_413 ( );
FILL FILL_0_OAI21X1_418 ( );
FILL FILL_1_OAI21X1_418 ( );
FILL FILL_0_NOR2X1_6 ( );
FILL FILL_1_NOR2X1_6 ( );
FILL FILL_0_INVX2_41 ( );
FILL FILL_0_OAI21X1_414 ( );
FILL FILL_1_OAI21X1_414 ( );
FILL FILL_2_OAI21X1_414 ( );
FILL FILL_0_NAND2X1_159 ( );
FILL FILL_0_OR2X2_1 ( );
FILL FILL_1_OR2X2_1 ( );
FILL FILL_2_OR2X2_1 ( );
FILL FILL_0_XNOR2X1_41 ( );
FILL FILL_1_XNOR2X1_41 ( );
FILL FILL_2_XNOR2X1_41 ( );
FILL FILL_3_XNOR2X1_41 ( );
FILL FILL_0_BUFX2_492 ( );
FILL FILL_1_BUFX2_492 ( );
FILL FILL_0_XNOR2X1_5 ( );
FILL FILL_1_XNOR2X1_5 ( );
FILL FILL_2_XNOR2X1_5 ( );
FILL FILL_3_XNOR2X1_5 ( );
FILL FILL_0_NAND2X1_228 ( );
FILL FILL_0_OAI21X1_339 ( );
FILL FILL_1_OAI21X1_339 ( );
FILL FILL_0_DFFPOSX1_367 ( );
FILL FILL_1_DFFPOSX1_367 ( );
FILL FILL_2_DFFPOSX1_367 ( );
FILL FILL_3_DFFPOSX1_367 ( );
FILL FILL_4_DFFPOSX1_367 ( );
FILL FILL_5_DFFPOSX1_367 ( );
FILL FILL_6_DFFPOSX1_367 ( );
FILL FILL_0_OAI21X1_345 ( );
FILL FILL_1_OAI21X1_345 ( );
FILL FILL_0_DFFPOSX1_411 ( );
FILL FILL_1_DFFPOSX1_411 ( );
FILL FILL_2_DFFPOSX1_411 ( );
FILL FILL_3_DFFPOSX1_411 ( );
FILL FILL_4_DFFPOSX1_411 ( );
FILL FILL_5_DFFPOSX1_411 ( );
FILL FILL_0_NAND2X1_127 ( );
FILL FILL_0_BUFX2_420 ( );
FILL FILL_0_DFFPOSX1_473 ( );
FILL FILL_1_DFFPOSX1_473 ( );
FILL FILL_2_DFFPOSX1_473 ( );
FILL FILL_3_DFFPOSX1_473 ( );
FILL FILL_4_DFFPOSX1_473 ( );
FILL FILL_5_DFFPOSX1_473 ( );
FILL FILL_6_DFFPOSX1_473 ( );
FILL FILL_0_OAI21X1_1771 ( );
FILL FILL_1_OAI21X1_1771 ( );
FILL FILL_0_OAI21X1_1770 ( );
FILL FILL_1_OAI21X1_1770 ( );
FILL FILL_0_OAI21X1_316 ( );
FILL FILL_1_OAI21X1_316 ( );
FILL FILL_0_DFFPOSX1_350 ( );
FILL FILL_1_DFFPOSX1_350 ( );
FILL FILL_2_DFFPOSX1_350 ( );
FILL FILL_3_DFFPOSX1_350 ( );
FILL FILL_4_DFFPOSX1_350 ( );
FILL FILL_5_DFFPOSX1_350 ( );
FILL FILL_0_OAI21X1_317 ( );
FILL FILL_1_OAI21X1_317 ( );
FILL FILL_0_DFFPOSX1_391 ( );
FILL FILL_1_DFFPOSX1_391 ( );
FILL FILL_2_DFFPOSX1_391 ( );
FILL FILL_3_DFFPOSX1_391 ( );
FILL FILL_4_DFFPOSX1_391 ( );
FILL FILL_5_DFFPOSX1_391 ( );
FILL FILL_0_OAI21X1_725 ( );
FILL FILL_1_OAI21X1_725 ( );
FILL FILL_0_OAI21X1_726 ( );
FILL FILL_1_OAI21X1_726 ( );
FILL FILL_2_OAI21X1_726 ( );
FILL FILL_0_BUFX2_600 ( );
FILL FILL_1_BUFX2_600 ( );
FILL FILL_0_OAI21X1_204 ( );
FILL FILL_1_OAI21X1_204 ( );
FILL FILL_0_BUFX2_594 ( );
FILL FILL_0_OAI21X1_994 ( );
FILL FILL_1_OAI21X1_994 ( );
FILL FILL_0_BUFX4_194 ( );
FILL FILL_1_BUFX4_194 ( );
FILL FILL_0_XNOR2X1_9 ( );
FILL FILL_1_XNOR2X1_9 ( );
FILL FILL_2_XNOR2X1_9 ( );
FILL FILL_0_INVX4_9 ( );
FILL FILL_0_BUFX2_467 ( );
FILL FILL_0_OAI21X1_351 ( );
FILL FILL_1_OAI21X1_351 ( );
FILL FILL_0_DFFPOSX1_442 ( );
FILL FILL_1_DFFPOSX1_442 ( );
FILL FILL_2_DFFPOSX1_442 ( );
FILL FILL_3_DFFPOSX1_442 ( );
FILL FILL_4_DFFPOSX1_442 ( );
FILL FILL_5_DFFPOSX1_442 ( );
FILL FILL_6_DFFPOSX1_442 ( );
FILL FILL_0_INVX2_21 ( );
FILL FILL_0_OAI21X1_350 ( );
FILL FILL_1_OAI21X1_350 ( );
FILL FILL_0_NAND2X1_183 ( );
FILL FILL_0_BUFX2_477 ( );
FILL FILL_0_OAI21X1_564 ( );
FILL FILL_1_OAI21X1_564 ( );
FILL FILL_0_DFFPOSX1_449 ( );
FILL FILL_1_DFFPOSX1_449 ( );
FILL FILL_2_DFFPOSX1_449 ( );
FILL FILL_3_DFFPOSX1_449 ( );
FILL FILL_4_DFFPOSX1_449 ( );
FILL FILL_5_DFFPOSX1_449 ( );
FILL FILL_6_DFFPOSX1_449 ( );
FILL FILL_0_OAI21X1_563 ( );
FILL FILL_1_OAI21X1_563 ( );
FILL FILL_2_OAI21X1_563 ( );
FILL FILL_0_OAI21X1_562 ( );
FILL FILL_1_OAI21X1_562 ( );
FILL FILL_0_NAND2X1_191 ( );
FILL FILL_1_NAND2X1_191 ( );
FILL FILL_0_NAND2X1_96 ( );
FILL FILL_0_OAI21X1_352 ( );
FILL FILL_1_OAI21X1_352 ( );
FILL FILL_2_OAI21X1_352 ( );
FILL FILL_0_OAI21X1_439 ( );
FILL FILL_1_OAI21X1_439 ( );
FILL FILL_0_BUFX2_812 ( );
FILL FILL_1_BUFX2_812 ( );
FILL FILL_0_OAI21X1_356 ( );
FILL FILL_1_OAI21X1_356 ( );
FILL FILL_2_OAI21X1_356 ( );
FILL FILL_0_OAI21X1_988 ( );
FILL FILL_1_OAI21X1_988 ( );
FILL FILL_0_OAI21X1_989 ( );
FILL FILL_1_OAI21X1_989 ( );
FILL FILL_0_BUFX2_531 ( );
FILL FILL_1_BUFX2_531 ( );
FILL FILL_0_BUFX4_333 ( );
FILL FILL_1_BUFX4_333 ( );
FILL FILL_0_NAND2X1_755 ( );
FILL FILL_1_NAND2X1_755 ( );
FILL FILL_0_OAI21X1_152 ( );
FILL FILL_1_OAI21X1_152 ( );
FILL FILL_0_OAI21X1_153 ( );
FILL FILL_1_OAI21X1_153 ( );
FILL FILL_0_OAI21X1_189 ( );
FILL FILL_1_OAI21X1_189 ( );
FILL FILL_0_OAI21X1_972 ( );
FILL FILL_1_OAI21X1_972 ( );
FILL FILL_0_OAI21X1_188 ( );
FILL FILL_1_OAI21X1_188 ( );
FILL FILL_2_OAI21X1_188 ( );
FILL FILL_0_INVX2_142 ( );
FILL FILL_0_NAND2X1_425 ( );
FILL FILL_1_NAND2X1_425 ( );
FILL FILL_0_DFFPOSX1_110 ( );
FILL FILL_1_DFFPOSX1_110 ( );
FILL FILL_2_DFFPOSX1_110 ( );
FILL FILL_3_DFFPOSX1_110 ( );
FILL FILL_4_DFFPOSX1_110 ( );
FILL FILL_5_DFFPOSX1_110 ( );
FILL FILL_0_NAND2X1_706 ( );
FILL FILL_0_NAND2X1_725 ( );
FILL FILL_0_OAI21X1_1784 ( );
FILL FILL_1_OAI21X1_1784 ( );
FILL FILL_2_OAI21X1_1784 ( );
FILL FILL_0_BUFX4_326 ( );
FILL FILL_1_BUFX4_326 ( );
FILL FILL_0_DFFPOSX1_1029 ( );
FILL FILL_1_DFFPOSX1_1029 ( );
FILL FILL_2_DFFPOSX1_1029 ( );
FILL FILL_3_DFFPOSX1_1029 ( );
FILL FILL_4_DFFPOSX1_1029 ( );
FILL FILL_5_DFFPOSX1_1029 ( );
FILL FILL_0_DFFPOSX1_224 ( );
FILL FILL_1_DFFPOSX1_224 ( );
FILL FILL_2_DFFPOSX1_224 ( );
FILL FILL_3_DFFPOSX1_224 ( );
FILL FILL_4_DFFPOSX1_224 ( );
FILL FILL_5_DFFPOSX1_224 ( );
FILL FILL_6_DFFPOSX1_224 ( );
FILL FILL_0_BUFX2_78 ( );
FILL FILL_1_BUFX2_78 ( );
FILL FILL_0_OAI21X1_1058 ( );
FILL FILL_1_OAI21X1_1058 ( );
FILL FILL_0_NAND2X1_424 ( );
FILL FILL_0_DFFPOSX1_766 ( );
FILL FILL_1_DFFPOSX1_766 ( );
FILL FILL_2_DFFPOSX1_766 ( );
FILL FILL_3_DFFPOSX1_766 ( );
FILL FILL_4_DFFPOSX1_766 ( );
FILL FILL_5_DFFPOSX1_766 ( );
FILL FILL_0_DFFPOSX1_159 ( );
FILL FILL_1_DFFPOSX1_159 ( );
FILL FILL_2_DFFPOSX1_159 ( );
FILL FILL_3_DFFPOSX1_159 ( );
FILL FILL_4_DFFPOSX1_159 ( );
FILL FILL_5_DFFPOSX1_159 ( );
FILL FILL_6_DFFPOSX1_159 ( );
FILL FILL_0_BUFX4_369 ( );
FILL FILL_1_BUFX4_369 ( );
FILL FILL_2_BUFX4_369 ( );
FILL FILL_0_BUFX2_147 ( );
FILL FILL_0_BUFX2_960 ( );
FILL FILL_1_BUFX2_960 ( );
FILL FILL_0_BUFX2_927 ( );
FILL FILL_0_DFFPOSX1_849 ( );
FILL FILL_1_DFFPOSX1_849 ( );
FILL FILL_2_DFFPOSX1_849 ( );
FILL FILL_3_DFFPOSX1_849 ( );
FILL FILL_4_DFFPOSX1_849 ( );
FILL FILL_5_DFFPOSX1_849 ( );
FILL FILL_0_NAND2X1_548 ( );
FILL FILL_1_NAND2X1_548 ( );
FILL FILL_0_OAI21X1_982 ( );
FILL FILL_1_OAI21X1_982 ( );
FILL FILL_0_OAI21X1_1071 ( );
FILL FILL_1_OAI21X1_1071 ( );
FILL FILL_0_BUFX2_159 ( );
FILL FILL_1_BUFX2_159 ( );
FILL FILL_0_OAI21X1_1164 ( );
FILL FILL_1_OAI21X1_1164 ( );
FILL FILL_0_NAND2X1_535 ( );
FILL FILL_0_NAND2X1_443 ( );
FILL FILL_1_NAND2X1_443 ( );
FILL FILL_0_BUFX4_384 ( );
FILL FILL_1_BUFX4_384 ( );
FILL FILL_0_BUFX2_101 ( );
FILL FILL_1_BUFX2_101 ( );
FILL FILL_0_NAND2X1_545 ( );
FILL FILL_1_NAND2X1_545 ( );
FILL FILL_0_INVX2_79 ( );
FILL FILL_0_NAND2X1_546 ( );
FILL FILL_0_BUFX2_100 ( );
FILL FILL_0_OAI21X1_1076 ( );
FILL FILL_1_OAI21X1_1076 ( );
FILL FILL_0_NAND2X1_442 ( );
FILL FILL_1_NAND2X1_442 ( );
FILL FILL_0_DFFPOSX1_784 ( );
FILL FILL_1_DFFPOSX1_784 ( );
FILL FILL_2_DFFPOSX1_784 ( );
FILL FILL_3_DFFPOSX1_784 ( );
FILL FILL_4_DFFPOSX1_784 ( );
FILL FILL_5_DFFPOSX1_784 ( );
FILL FILL_0_OAI21X1_1534 ( );
FILL FILL_1_OAI21X1_1534 ( );
FILL FILL_0_OAI21X1_1535 ( );
FILL FILL_1_OAI21X1_1535 ( );
FILL FILL_0_BUFX2_242 ( );
FILL FILL_1_BUFX2_242 ( );
FILL FILL_0_OAI21X1_1010 ( );
FILL FILL_1_OAI21X1_1010 ( );
FILL FILL_0_NAND2X1_37 ( );
FILL FILL_0_DFFPOSX1_731 ( );
FILL FILL_1_DFFPOSX1_731 ( );
FILL FILL_2_DFFPOSX1_731 ( );
FILL FILL_3_DFFPOSX1_731 ( );
FILL FILL_4_DFFPOSX1_731 ( );
FILL FILL_5_DFFPOSX1_731 ( );
FILL FILL_6_DFFPOSX1_731 ( );
FILL FILL_0_OAI21X1_210 ( );
FILL FILL_1_OAI21X1_210 ( );
FILL FILL_0_DFFPOSX1_297 ( );
FILL FILL_1_DFFPOSX1_297 ( );
FILL FILL_2_DFFPOSX1_297 ( );
FILL FILL_3_DFFPOSX1_297 ( );
FILL FILL_4_DFFPOSX1_297 ( );
FILL FILL_5_DFFPOSX1_297 ( );
FILL FILL_6_DFFPOSX1_297 ( );
FILL FILL_0_OAI21X1_211 ( );
FILL FILL_1_OAI21X1_211 ( );
FILL FILL_0_BUFX2_813 ( );
FILL FILL_0_OAI21X1_128 ( );
FILL FILL_1_OAI21X1_128 ( );
FILL FILL_0_DFFPOSX1_800 ( );
FILL FILL_1_DFFPOSX1_800 ( );
FILL FILL_2_DFFPOSX1_800 ( );
FILL FILL_3_DFFPOSX1_800 ( );
FILL FILL_4_DFFPOSX1_800 ( );
FILL FILL_5_DFFPOSX1_800 ( );
FILL FILL_6_DFFPOSX1_800 ( );
FILL FILL_0_BUFX2_48 ( );
FILL FILL_0_BUFX2_53 ( );
FILL FILL_0_DFFPOSX1_105 ( );
FILL FILL_1_DFFPOSX1_105 ( );
FILL FILL_2_DFFPOSX1_105 ( );
FILL FILL_3_DFFPOSX1_105 ( );
FILL FILL_4_DFFPOSX1_105 ( );
FILL FILL_5_DFFPOSX1_105 ( );
FILL FILL_0_OAI21X1_1779 ( );
FILL FILL_1_OAI21X1_1779 ( );
FILL FILL_0_NAND2X1_720 ( );
FILL FILL_0_DFFPOSX1_169 ( );
FILL FILL_1_DFFPOSX1_169 ( );
FILL FILL_2_DFFPOSX1_169 ( );
FILL FILL_3_DFFPOSX1_169 ( );
FILL FILL_4_DFFPOSX1_169 ( );
FILL FILL_5_DFFPOSX1_169 ( );
FILL FILL_6_DFFPOSX1_169 ( );
FILL FILL_0_BUFX2_246 ( );
FILL FILL_0_BUFX2_950 ( );
FILL FILL_0_BUFX4_206 ( );
FILL FILL_1_BUFX4_206 ( );
FILL FILL_0_OAI21X1_918 ( );
FILL FILL_1_OAI21X1_918 ( );
FILL FILL_0_OAI21X1_919 ( );
FILL FILL_1_OAI21X1_919 ( );
FILL FILL_0_DFFPOSX1_685 ( );
FILL FILL_1_DFFPOSX1_685 ( );
FILL FILL_2_DFFPOSX1_685 ( );
FILL FILL_3_DFFPOSX1_685 ( );
FILL FILL_4_DFFPOSX1_685 ( );
FILL FILL_5_DFFPOSX1_685 ( );
FILL FILL_6_DFFPOSX1_685 ( );
FILL FILL_0_OAI21X1_1619 ( );
FILL FILL_1_OAI21X1_1619 ( );
FILL FILL_2_OAI21X1_1619 ( );
FILL FILL_0_NAND2X1_687 ( );
FILL FILL_0_DFFPOSX1_9 ( );
FILL FILL_1_DFFPOSX1_9 ( );
FILL FILL_2_DFFPOSX1_9 ( );
FILL FILL_3_DFFPOSX1_9 ( );
FILL FILL_4_DFFPOSX1_9 ( );
FILL FILL_5_DFFPOSX1_9 ( );
FILL FILL_6_DFFPOSX1_9 ( );
FILL FILL_0_BUFX2_772 ( );
FILL FILL_1_BUFX2_772 ( );
FILL FILL_0_BUFX2_740 ( );
FILL FILL_0_BUFX2_941 ( );
FILL FILL_1_BUFX2_941 ( );
FILL FILL_0_BUFX2_365 ( );
FILL FILL_0_BUFX2_343 ( );
FILL FILL_1_BUFX2_343 ( );
FILL FILL_0_BUFX2_367 ( );
FILL FILL_1_BUFX2_367 ( );
FILL FILL_0_INVX1_111 ( );
FILL FILL_0_DFFPOSX1_709 ( );
FILL FILL_1_DFFPOSX1_709 ( );
FILL FILL_2_DFFPOSX1_709 ( );
FILL FILL_3_DFFPOSX1_709 ( );
FILL FILL_4_DFFPOSX1_709 ( );
FILL FILL_5_DFFPOSX1_709 ( );
FILL FILL_6_DFFPOSX1_709 ( );
FILL FILL_0_INVX2_123 ( );
FILL FILL_0_OAI21X1_1027 ( );
FILL FILL_1_OAI21X1_1027 ( );
FILL FILL_2_OAI21X1_1027 ( );
FILL FILL_0_DFFPOSX1_739 ( );
FILL FILL_1_DFFPOSX1_739 ( );
FILL FILL_2_DFFPOSX1_739 ( );
FILL FILL_3_DFFPOSX1_739 ( );
FILL FILL_4_DFFPOSX1_739 ( );
FILL FILL_5_DFFPOSX1_739 ( );
FILL FILL_6_DFFPOSX1_739 ( );
FILL FILL_0_DFFPOSX1_108 ( );
FILL FILL_1_DFFPOSX1_108 ( );
FILL FILL_2_DFFPOSX1_108 ( );
FILL FILL_3_DFFPOSX1_108 ( );
FILL FILL_4_DFFPOSX1_108 ( );
FILL FILL_5_DFFPOSX1_108 ( );
FILL FILL_0_DFFPOSX1_113 ( );
FILL FILL_1_DFFPOSX1_113 ( );
FILL FILL_2_DFFPOSX1_113 ( );
FILL FILL_3_DFFPOSX1_113 ( );
FILL FILL_4_DFFPOSX1_113 ( );
FILL FILL_5_DFFPOSX1_113 ( );
FILL FILL_6_DFFPOSX1_113 ( );
FILL FILL_0_OAI21X1_1787 ( );
FILL FILL_1_OAI21X1_1787 ( );
FILL FILL_0_BUFX2_995 ( );
FILL FILL_0_DFFPOSX1_99 ( );
FILL FILL_1_DFFPOSX1_99 ( );
FILL FILL_2_DFFPOSX1_99 ( );
FILL FILL_3_DFFPOSX1_99 ( );
FILL FILL_4_DFFPOSX1_99 ( );
FILL FILL_5_DFFPOSX1_99 ( );
FILL FILL_0_OAI21X1_1773 ( );
FILL FILL_1_OAI21X1_1773 ( );
FILL FILL_0_OAI21X1_1772 ( );
FILL FILL_1_OAI21X1_1772 ( );
FILL FILL_0_DFFPOSX1_363 ( );
FILL FILL_1_DFFPOSX1_363 ( );
FILL FILL_2_DFFPOSX1_363 ( );
FILL FILL_3_DFFPOSX1_363 ( );
FILL FILL_4_DFFPOSX1_363 ( );
FILL FILL_5_DFFPOSX1_363 ( );
FILL FILL_0_NAND2X1_79 ( );
FILL FILL_1_NAND2X1_79 ( );
FILL FILL_0_OAI21X1_335 ( );
FILL FILL_1_OAI21X1_335 ( );
FILL FILL_0_NAND2X1_143 ( );
FILL FILL_1_NAND2X1_143 ( );
FILL FILL_0_OAI21X1_406 ( );
FILL FILL_1_OAI21X1_406 ( );
FILL FILL_0_OAI21X1_408 ( );
FILL FILL_1_OAI21X1_408 ( );
FILL FILL_0_OAI21X1_400 ( );
FILL FILL_1_OAI21X1_400 ( );
FILL FILL_0_DFFPOSX1_494 ( );
FILL FILL_1_DFFPOSX1_494 ( );
FILL FILL_2_DFFPOSX1_494 ( );
FILL FILL_3_DFFPOSX1_494 ( );
FILL FILL_4_DFFPOSX1_494 ( );
FILL FILL_5_DFFPOSX1_494 ( );
FILL FILL_6_DFFPOSX1_494 ( );
FILL FILL_0_NAND2X1_151 ( );
FILL FILL_1_NAND2X1_151 ( );
FILL FILL_0_OAI21X1_529 ( );
FILL FILL_1_OAI21X1_529 ( );
FILL FILL_0_OAI21X1_530 ( );
FILL FILL_1_OAI21X1_530 ( );
FILL FILL_0_BUFX4_388 ( );
FILL FILL_1_BUFX4_388 ( );
FILL FILL_0_DFFPOSX1_371 ( );
FILL FILL_1_DFFPOSX1_371 ( );
FILL FILL_2_DFFPOSX1_371 ( );
FILL FILL_3_DFFPOSX1_371 ( );
FILL FILL_4_DFFPOSX1_371 ( );
FILL FILL_5_DFFPOSX1_371 ( );
FILL FILL_6_DFFPOSX1_371 ( );
FILL FILL_0_OAI21X1_528 ( );
FILL FILL_1_OAI21X1_528 ( );
FILL FILL_0_XNOR2X1_2 ( );
FILL FILL_1_XNOR2X1_2 ( );
FILL FILL_2_XNOR2X1_2 ( );
FILL FILL_3_XNOR2X1_2 ( );
FILL FILL_0_OAI21X1_417 ( );
FILL FILL_1_OAI21X1_417 ( );
FILL FILL_0_NAND2X1_157 ( );
FILL FILL_1_NAND2X1_157 ( );
FILL FILL_0_DFFPOSX1_556 ( );
FILL FILL_1_DFFPOSX1_556 ( );
FILL FILL_2_DFFPOSX1_556 ( );
FILL FILL_3_DFFPOSX1_556 ( );
FILL FILL_4_DFFPOSX1_556 ( );
FILL FILL_5_DFFPOSX1_556 ( );
FILL FILL_0_INVX2_16 ( );
FILL FILL_0_OAI21X1_684 ( );
FILL FILL_1_OAI21X1_684 ( );
FILL FILL_0_OAI21X1_685 ( );
FILL FILL_1_OAI21X1_685 ( );
FILL FILL_0_XNOR2X1_4 ( );
FILL FILL_1_XNOR2X1_4 ( );
FILL FILL_2_XNOR2X1_4 ( );
FILL FILL_0_NOR2X1_9 ( );
FILL FILL_0_BUFX2_552 ( );
FILL FILL_1_BUFX2_552 ( );
FILL FILL_0_BUFX4_387 ( );
FILL FILL_1_BUFX4_387 ( );
FILL FILL_0_DFFPOSX1_466 ( );
FILL FILL_1_DFFPOSX1_466 ( );
FILL FILL_2_DFFPOSX1_466 ( );
FILL FILL_3_DFFPOSX1_466 ( );
FILL FILL_4_DFFPOSX1_466 ( );
FILL FILL_5_DFFPOSX1_466 ( );
FILL FILL_6_DFFPOSX1_466 ( );
FILL FILL_0_DFFPOSX1_373 ( );
FILL FILL_1_DFFPOSX1_373 ( );
FILL FILL_2_DFFPOSX1_373 ( );
FILL FILL_3_DFFPOSX1_373 ( );
FILL FILL_4_DFFPOSX1_373 ( );
FILL FILL_5_DFFPOSX1_373 ( );
FILL FILL_6_DFFPOSX1_373 ( );
FILL FILL_0_OAI21X1_383 ( );
FILL FILL_1_OAI21X1_383 ( );
FILL FILL_0_DFFPOSX1_472 ( );
FILL FILL_1_DFFPOSX1_472 ( );
FILL FILL_2_DFFPOSX1_472 ( );
FILL FILL_3_DFFPOSX1_472 ( );
FILL FILL_4_DFFPOSX1_472 ( );
FILL FILL_5_DFFPOSX1_472 ( );
FILL FILL_0_NAND2X1_246 ( );
FILL FILL_1_NAND2X1_246 ( );
FILL FILL_0_BUFX4_30 ( );
FILL FILL_1_BUFX4_30 ( );
FILL FILL_0_CLKBUF1_6 ( );
FILL FILL_1_CLKBUF1_6 ( );
FILL FILL_2_CLKBUF1_6 ( );
FILL FILL_3_CLKBUF1_6 ( );
FILL FILL_4_CLKBUF1_6 ( );
FILL FILL_0_CLKBUF1_92 ( );
FILL FILL_1_CLKBUF1_92 ( );
FILL FILL_2_CLKBUF1_92 ( );
FILL FILL_3_CLKBUF1_92 ( );
FILL FILL_4_CLKBUF1_92 ( );
FILL FILL_0_INVX4_16 ( );
FILL FILL_0_NAND2X1_205 ( );
FILL FILL_0_NAND2X1_107 ( );
FILL FILL_1_NAND2X1_107 ( );
FILL FILL_0_OAI21X1_363 ( );
FILL FILL_1_OAI21X1_363 ( );
FILL FILL_0_DFFPOSX1_571 ( );
FILL FILL_1_DFFPOSX1_571 ( );
FILL FILL_2_DFFPOSX1_571 ( );
FILL FILL_3_DFFPOSX1_571 ( );
FILL FILL_4_DFFPOSX1_571 ( );
FILL FILL_5_DFFPOSX1_571 ( );
FILL FILL_0_DFFPOSX1_452 ( );
FILL FILL_1_DFFPOSX1_452 ( );
FILL FILL_2_DFFPOSX1_452 ( );
FILL FILL_3_DFFPOSX1_452 ( );
FILL FILL_4_DFFPOSX1_452 ( );
FILL FILL_5_DFFPOSX1_452 ( );
FILL FILL_0_NAND2X1_204 ( );
FILL FILL_1_NAND2X1_204 ( );
FILL FILL_0_BUFX2_599 ( );
FILL FILL_0_XNOR2X1_45 ( );
FILL FILL_1_XNOR2X1_45 ( );
FILL FILL_2_XNOR2X1_45 ( );
FILL FILL_0_NAND2X1_185 ( );
FILL FILL_1_NAND2X1_185 ( );
FILL FILL_0_DFFPOSX1_440 ( );
FILL FILL_1_DFFPOSX1_440 ( );
FILL FILL_2_DFFPOSX1_440 ( );
FILL FILL_3_DFFPOSX1_440 ( );
FILL FILL_4_DFFPOSX1_440 ( );
FILL FILL_5_DFFPOSX1_440 ( );
FILL FILL_6_DFFPOSX1_440 ( );
FILL FILL_0_DFFPOSX1_505 ( );
FILL FILL_1_DFFPOSX1_505 ( );
FILL FILL_2_DFFPOSX1_505 ( );
FILL FILL_3_DFFPOSX1_505 ( );
FILL FILL_4_DFFPOSX1_505 ( );
FILL FILL_5_DFFPOSX1_505 ( );
FILL FILL_6_DFFPOSX1_505 ( );
FILL FILL_0_DFFPOSX1_508 ( );
FILL FILL_1_DFFPOSX1_508 ( );
FILL FILL_2_DFFPOSX1_508 ( );
FILL FILL_3_DFFPOSX1_508 ( );
FILL FILL_4_DFFPOSX1_508 ( );
FILL FILL_5_DFFPOSX1_508 ( );
FILL FILL_0_NAND2X1_179 ( );
FILL FILL_1_NAND2X1_179 ( );
FILL FILL_0_BUFX2_953 ( );
FILL FILL_0_OAI21X1_565 ( );
FILL FILL_1_OAI21X1_565 ( );
FILL FILL_0_NAND2X1_198 ( );
FILL FILL_1_NAND2X1_198 ( );
FILL FILL_0_OAI21X1_444 ( );
FILL FILL_1_OAI21X1_444 ( );
FILL FILL_0_DFFPOSX1_380 ( );
FILL FILL_1_DFFPOSX1_380 ( );
FILL FILL_2_DFFPOSX1_380 ( );
FILL FILL_3_DFFPOSX1_380 ( );
FILL FILL_4_DFFPOSX1_380 ( );
FILL FILL_5_DFFPOSX1_380 ( );
FILL FILL_6_DFFPOSX1_380 ( );
FILL FILL_0_DFFPOSX1_140 ( );
FILL FILL_1_DFFPOSX1_140 ( );
FILL FILL_2_DFFPOSX1_140 ( );
FILL FILL_3_DFFPOSX1_140 ( );
FILL FILL_4_DFFPOSX1_140 ( );
FILL FILL_5_DFFPOSX1_140 ( );
FILL FILL_0_DFFPOSX1_286 ( );
FILL FILL_1_DFFPOSX1_286 ( );
FILL FILL_2_DFFPOSX1_286 ( );
FILL FILL_3_DFFPOSX1_286 ( );
FILL FILL_4_DFFPOSX1_286 ( );
FILL FILL_5_DFFPOSX1_286 ( );
FILL FILL_6_DFFPOSX1_286 ( );
FILL FILL_0_NAND2X1_675 ( );
FILL FILL_1_NAND2X1_675 ( );
FILL FILL_0_OAI21X1_1606 ( );
FILL FILL_1_OAI21X1_1606 ( );
FILL FILL_0_DFFPOSX1_767 ( );
FILL FILL_1_DFFPOSX1_767 ( );
FILL FILL_2_DFFPOSX1_767 ( );
FILL FILL_3_DFFPOSX1_767 ( );
FILL FILL_4_DFFPOSX1_767 ( );
FILL FILL_5_DFFPOSX1_767 ( );
FILL FILL_6_DFFPOSX1_767 ( );
FILL FILL_0_OAI21X1_1059 ( );
FILL FILL_1_OAI21X1_1059 ( );
FILL FILL_0_INVX1_174 ( );
FILL FILL_0_DFFPOSX1_28 ( );
FILL FILL_1_DFFPOSX1_28 ( );
FILL FILL_2_DFFPOSX1_28 ( );
FILL FILL_3_DFFPOSX1_28 ( );
FILL FILL_4_DFFPOSX1_28 ( );
FILL FILL_5_DFFPOSX1_28 ( );
FILL FILL_0_OAI21X1_1638 ( );
FILL FILL_1_OAI21X1_1638 ( );
FILL FILL_2_OAI21X1_1638 ( );
FILL FILL_0_NAND2X1_685 ( );
FILL FILL_1_NAND2X1_685 ( );
FILL FILL_0_OAI21X1_1617 ( );
FILL FILL_1_OAI21X1_1617 ( );
FILL FILL_0_DFFPOSX1_7 ( );
FILL FILL_1_DFFPOSX1_7 ( );
FILL FILL_2_DFFPOSX1_7 ( );
FILL FILL_3_DFFPOSX1_7 ( );
FILL FILL_4_DFFPOSX1_7 ( );
FILL FILL_5_DFFPOSX1_7 ( );
FILL FILL_6_DFFPOSX1_7 ( );
FILL FILL_0_NAND2X1_511 ( );
FILL FILL_0_DFFPOSX1_287 ( );
FILL FILL_1_DFFPOSX1_287 ( );
FILL FILL_2_DFFPOSX1_287 ( );
FILL FILL_3_DFFPOSX1_287 ( );
FILL FILL_4_DFFPOSX1_287 ( );
FILL FILL_5_DFFPOSX1_287 ( );
FILL FILL_0_DFFPOSX1_257 ( );
FILL FILL_1_DFFPOSX1_257 ( );
FILL FILL_2_DFFPOSX1_257 ( );
FILL FILL_3_DFFPOSX1_257 ( );
FILL FILL_4_DFFPOSX1_257 ( );
FILL FILL_5_DFFPOSX1_257 ( );
FILL FILL_0_NAND2X1_3 ( );
FILL FILL_1_NAND2X1_3 ( );
FILL FILL_0_OAI21X1_3 ( );
FILL FILL_1_OAI21X1_3 ( );
FILL FILL_0_BUFX2_140 ( );
FILL FILL_1_BUFX2_140 ( );
FILL FILL_0_BUFX4_152 ( );
FILL FILL_1_BUFX4_152 ( );
FILL FILL_0_OAI21X1_131 ( );
FILL FILL_1_OAI21X1_131 ( );
FILL FILL_0_DFFPOSX1_785 ( );
FILL FILL_1_DFFPOSX1_785 ( );
FILL FILL_2_DFFPOSX1_785 ( );
FILL FILL_3_DFFPOSX1_785 ( );
FILL FILL_4_DFFPOSX1_785 ( );
FILL FILL_5_DFFPOSX1_785 ( );
FILL FILL_6_DFFPOSX1_785 ( );
FILL FILL_0_INVX1_162 ( );
FILL FILL_0_DFFPOSX1_848 ( );
FILL FILL_1_DFFPOSX1_848 ( );
FILL FILL_2_DFFPOSX1_848 ( );
FILL FILL_3_DFFPOSX1_848 ( );
FILL FILL_4_DFFPOSX1_848 ( );
FILL FILL_5_DFFPOSX1_848 ( );
FILL FILL_6_DFFPOSX1_848 ( );
FILL FILL_0_INVX8_3 ( );
FILL FILL_1_INVX8_3 ( );
FILL FILL_0_OAI21X1_1167 ( );
FILL FILL_1_OAI21X1_1167 ( );
FILL FILL_0_OAI21X1_1159 ( );
FILL FILL_1_OAI21X1_1159 ( );
FILL FILL_2_OAI21X1_1159 ( );
FILL FILL_0_OAI21X1_1075 ( );
FILL FILL_1_OAI21X1_1075 ( );
FILL FILL_0_NAND2X1_441 ( );
FILL FILL_1_NAND2X1_441 ( );
FILL FILL_0_DFFPOSX1_783 ( );
FILL FILL_1_DFFPOSX1_783 ( );
FILL FILL_2_DFFPOSX1_783 ( );
FILL FILL_3_DFFPOSX1_783 ( );
FILL FILL_4_DFFPOSX1_783 ( );
FILL FILL_5_DFFPOSX1_783 ( );
FILL FILL_6_DFFPOSX1_783 ( );
FILL FILL_0_DFFPOSX1_976 ( );
FILL FILL_1_DFFPOSX1_976 ( );
FILL FILL_2_DFFPOSX1_976 ( );
FILL FILL_3_DFFPOSX1_976 ( );
FILL FILL_4_DFFPOSX1_976 ( );
FILL FILL_5_DFFPOSX1_976 ( );
FILL FILL_0_OAI21X1_1505 ( );
FILL FILL_1_OAI21X1_1505 ( );
FILL FILL_0_OAI21X1_1504 ( );
FILL FILL_1_OAI21X1_1504 ( );
FILL FILL_0_BUFX4_158 ( );
FILL FILL_1_BUFX4_158 ( );
FILL FILL_0_OAI21X1_1487 ( );
FILL FILL_1_OAI21X1_1487 ( );
FILL FILL_0_DFFPOSX1_141 ( );
FILL FILL_1_DFFPOSX1_141 ( );
FILL FILL_2_DFFPOSX1_141 ( );
FILL FILL_3_DFFPOSX1_141 ( );
FILL FILL_4_DFFPOSX1_141 ( );
FILL FILL_5_DFFPOSX1_141 ( );
FILL FILL_6_DFFPOSX1_141 ( );
FILL FILL_0_BUFX4_343 ( );
FILL FILL_1_BUFX4_343 ( );
FILL FILL_2_BUFX4_343 ( );
FILL FILL_0_NAND2X1_756 ( );
FILL FILL_1_NAND2X1_756 ( );
FILL FILL_0_BUFX4_28 ( );
FILL FILL_1_BUFX4_28 ( );
FILL FILL_0_BUFX2_115 ( );
FILL FILL_1_BUFX2_115 ( );
FILL FILL_0_OAI21X1_1092 ( );
FILL FILL_1_OAI21X1_1092 ( );
FILL FILL_2_OAI21X1_1092 ( );
FILL FILL_0_NAND2X1_458 ( );
FILL FILL_0_DFFPOSX1_801 ( );
FILL FILL_1_DFFPOSX1_801 ( );
FILL FILL_2_DFFPOSX1_801 ( );
FILL FILL_3_DFFPOSX1_801 ( );
FILL FILL_4_DFFPOSX1_801 ( );
FILL FILL_5_DFFPOSX1_801 ( );
FILL FILL_0_OAI21X1_1093 ( );
FILL FILL_1_OAI21X1_1093 ( );
FILL FILL_0_NAND2X1_459 ( );
FILL FILL_0_BUFX4_139 ( );
FILL FILL_1_BUFX4_139 ( );
FILL FILL_0_OAI21X1_82 ( );
FILL FILL_1_OAI21X1_82 ( );
FILL FILL_0_OAI21X1_83 ( );
FILL FILL_1_OAI21X1_83 ( );
FILL FILL_0_DFFPOSX1_233 ( );
FILL FILL_1_DFFPOSX1_233 ( );
FILL FILL_2_DFFPOSX1_233 ( );
FILL FILL_3_DFFPOSX1_233 ( );
FILL FILL_4_DFFPOSX1_233 ( );
FILL FILL_5_DFFPOSX1_233 ( );
FILL FILL_0_BUFX2_118 ( );
FILL FILL_0_DFFPOSX1_73 ( );
FILL FILL_1_DFFPOSX1_73 ( );
FILL FILL_2_DFFPOSX1_73 ( );
FILL FILL_3_DFFPOSX1_73 ( );
FILL FILL_4_DFFPOSX1_73 ( );
FILL FILL_5_DFFPOSX1_73 ( );
FILL FILL_0_OAI21X1_1720 ( );
FILL FILL_1_OAI21X1_1720 ( );
FILL FILL_0_OAI21X1_1721 ( );
FILL FILL_1_OAI21X1_1721 ( );
FILL FILL_0_DFFPOSX1_41 ( );
FILL FILL_1_DFFPOSX1_41 ( );
FILL FILL_2_DFFPOSX1_41 ( );
FILL FILL_3_DFFPOSX1_41 ( );
FILL FILL_4_DFFPOSX1_41 ( );
FILL FILL_5_DFFPOSX1_41 ( );
FILL FILL_0_BUFX2_51 ( );
FILL FILL_0_OAI21X1_1657 ( );
FILL FILL_1_OAI21X1_1657 ( );
FILL FILL_0_OAI21X1_1656 ( );
FILL FILL_1_OAI21X1_1656 ( );
FILL FILL_0_DFFPOSX1_1009 ( );
FILL FILL_1_DFFPOSX1_1009 ( );
FILL FILL_2_DFFPOSX1_1009 ( );
FILL FILL_3_DFFPOSX1_1009 ( );
FILL FILL_4_DFFPOSX1_1009 ( );
FILL FILL_5_DFFPOSX1_1009 ( );
FILL FILL_0_OAI21X1_1586 ( );
FILL FILL_1_OAI21X1_1586 ( );
FILL FILL_0_OAI21X1_958 ( );
FILL FILL_1_OAI21X1_958 ( );
FILL FILL_0_OAI21X1_959 ( );
FILL FILL_1_OAI21X1_959 ( );
FILL FILL_2_OAI21X1_959 ( );
FILL FILL_0_BUFX2_361 ( );
FILL FILL_1_BUFX2_361 ( );
FILL FILL_0_DFFPOSX1_738 ( );
FILL FILL_1_DFFPOSX1_738 ( );
FILL FILL_2_DFFPOSX1_738 ( );
FILL FILL_3_DFFPOSX1_738 ( );
FILL FILL_4_DFFPOSX1_738 ( );
FILL FILL_5_DFFPOSX1_738 ( );
FILL FILL_0_OAI21X1_1024 ( );
FILL FILL_1_OAI21X1_1024 ( );
FILL FILL_0_OAI21X1_1025 ( );
FILL FILL_1_OAI21X1_1025 ( );
FILL FILL_0_DFFPOSX1_705 ( );
FILL FILL_1_DFFPOSX1_705 ( );
FILL FILL_2_DFFPOSX1_705 ( );
FILL FILL_3_DFFPOSX1_705 ( );
FILL FILL_4_DFFPOSX1_705 ( );
FILL FILL_5_DFFPOSX1_705 ( );
FILL FILL_6_DFFPOSX1_705 ( );
FILL FILL_0_BUFX2_773 ( );
FILL FILL_1_BUFX2_773 ( );
FILL FILL_0_BUFX2_706 ( );
FILL FILL_0_OAI21X1_913 ( );
FILL FILL_1_OAI21X1_913 ( );
FILL FILL_0_OAI21X1_912 ( );
FILL FILL_1_OAI21X1_912 ( );
FILL FILL_2_OAI21X1_912 ( );
FILL FILL_0_DFFPOSX1_682 ( );
FILL FILL_1_DFFPOSX1_682 ( );
FILL FILL_2_DFFPOSX1_682 ( );
FILL FILL_3_DFFPOSX1_682 ( );
FILL FILL_4_DFFPOSX1_682 ( );
FILL FILL_5_DFFPOSX1_682 ( );
FILL FILL_0_OAI21X1_1026 ( );
FILL FILL_1_OAI21X1_1026 ( );
FILL FILL_0_BUFX2_449 ( );
FILL FILL_0_BUFX2_544 ( );
FILL FILL_1_BUFX2_544 ( );
FILL FILL_0_BUFX2_931 ( );
FILL FILL_1_BUFX2_931 ( );
FILL FILL_0_DFFPOSX1_260 ( );
FILL FILL_1_DFFPOSX1_260 ( );
FILL FILL_2_DFFPOSX1_260 ( );
FILL FILL_3_DFFPOSX1_260 ( );
FILL FILL_4_DFFPOSX1_260 ( );
FILL FILL_5_DFFPOSX1_260 ( );
FILL FILL_6_DFFPOSX1_260 ( );
FILL FILL_0_BUFX4_153 ( );
FILL FILL_1_BUFX4_153 ( );
FILL FILL_0_BUFX4_315 ( );
FILL FILL_1_BUFX4_315 ( );
FILL FILL_0_CLKBUF1_56 ( );
FILL FILL_1_CLKBUF1_56 ( );
FILL FILL_2_CLKBUF1_56 ( );
FILL FILL_3_CLKBUF1_56 ( );
FILL FILL_0_NAND2X1_747 ( );
FILL FILL_1_NAND2X1_747 ( );
FILL FILL_0_OAI21X1_1806 ( );
FILL FILL_1_OAI21X1_1806 ( );
FILL FILL_0_DFFPOSX1_362 ( );
FILL FILL_1_DFFPOSX1_362 ( );
FILL FILL_2_DFFPOSX1_362 ( );
FILL FILL_3_DFFPOSX1_362 ( );
FILL FILL_4_DFFPOSX1_362 ( );
FILL FILL_5_DFFPOSX1_362 ( );
FILL FILL_6_DFFPOSX1_362 ( );
FILL FILL_0_NAND2X1_78 ( );
FILL FILL_1_NAND2X1_78 ( );
FILL FILL_0_OAI21X1_334 ( );
FILL FILL_1_OAI21X1_334 ( );
FILL FILL_0_DFFPOSX1_361 ( );
FILL FILL_1_DFFPOSX1_361 ( );
FILL FILL_2_DFFPOSX1_361 ( );
FILL FILL_3_DFFPOSX1_361 ( );
FILL FILL_4_DFFPOSX1_361 ( );
FILL FILL_5_DFFPOSX1_361 ( );
FILL FILL_0_NAND2X1_77 ( );
FILL FILL_0_OAI21X1_333 ( );
FILL FILL_1_OAI21X1_333 ( );
FILL FILL_2_OAI21X1_333 ( );
FILL FILL_0_BUFX4_355 ( );
FILL FILL_1_BUFX4_355 ( );
FILL FILL_0_NAND2X1_88 ( );
FILL FILL_0_NAND2X1_147 ( );
FILL FILL_1_NAND2X1_147 ( );
FILL FILL_0_BUFX2_582 ( );
FILL FILL_1_BUFX2_582 ( );
FILL FILL_0_NOR2X1_60 ( );
FILL FILL_1_NOR2X1_60 ( );
FILL FILL_0_NAND2X1_270 ( );
FILL FILL_1_NAND2X1_270 ( );
FILL FILL_0_INVX2_13 ( );
FILL FILL_0_NAND2X1_149 ( );
FILL FILL_1_NAND2X1_149 ( );
FILL FILL_0_BUFX2_583 ( );
FILL FILL_1_BUFX2_583 ( );
FILL FILL_0_OAI21X1_523 ( );
FILL FILL_1_OAI21X1_523 ( );
FILL FILL_0_DFFPOSX1_492 ( );
FILL FILL_1_DFFPOSX1_492 ( );
FILL FILL_2_DFFPOSX1_492 ( );
FILL FILL_3_DFFPOSX1_492 ( );
FILL FILL_4_DFFPOSX1_492 ( );
FILL FILL_5_DFFPOSX1_492 ( );
FILL FILL_6_DFFPOSX1_492 ( );
FILL FILL_0_OAI21X1_524 ( );
FILL FILL_1_OAI21X1_524 ( );
FILL FILL_0_OAI21X1_343 ( );
FILL FILL_1_OAI21X1_343 ( );
FILL FILL_0_BUFX2_550 ( );
FILL FILL_0_OAI21X1_699 ( );
FILL FILL_1_OAI21X1_699 ( );
FILL FILL_0_INVX2_14 ( );
FILL FILL_0_NAND2X1_155 ( );
FILL FILL_0_BUFX2_528 ( );
FILL FILL_1_BUFX2_528 ( );
FILL FILL_0_AOI21X1_30 ( );
FILL FILL_1_AOI21X1_30 ( );
FILL FILL_0_INVX1_35 ( );
FILL FILL_0_OAI21X1_687 ( );
FILL FILL_1_OAI21X1_687 ( );
FILL FILL_2_OAI21X1_687 ( );
FILL FILL_0_NOR2X1_5 ( );
FILL FILL_1_NOR2X1_5 ( );
FILL FILL_0_OAI21X1_682 ( );
FILL FILL_1_OAI21X1_682 ( );
FILL FILL_0_OAI21X1_683 ( );
FILL FILL_1_OAI21X1_683 ( );
FILL FILL_0_NAND2X1_312 ( );
FILL FILL_1_NAND2X1_312 ( );
FILL FILL_0_DFFPOSX1_557 ( );
FILL FILL_1_DFFPOSX1_557 ( );
FILL FILL_2_DFFPOSX1_557 ( );
FILL FILL_3_DFFPOSX1_557 ( );
FILL FILL_4_DFFPOSX1_557 ( );
FILL FILL_5_DFFPOSX1_557 ( );
FILL FILL_6_DFFPOSX1_557 ( );
FILL FILL_0_BUFX2_496 ( );
FILL FILL_1_BUFX2_496 ( );
FILL FILL_0_OAI21X1_468 ( );
FILL FILL_1_OAI21X1_468 ( );
FILL FILL_0_OAI21X1_469 ( );
FILL FILL_1_OAI21X1_469 ( );
FILL FILL_0_BUFX2_398 ( );
FILL FILL_1_BUFX2_398 ( );
FILL FILL_0_BUFX2_508 ( );
FILL FILL_0_NAND2X1_226 ( );
FILL FILL_1_NAND2X1_226 ( );
FILL FILL_0_DFFPOSX1_467 ( );
FILL FILL_1_DFFPOSX1_467 ( );
FILL FILL_2_DFFPOSX1_467 ( );
FILL FILL_3_DFFPOSX1_467 ( );
FILL FILL_4_DFFPOSX1_467 ( );
FILL FILL_5_DFFPOSX1_467 ( );
FILL FILL_0_NAND2X1_229 ( );
FILL FILL_1_NAND2X1_229 ( );
FILL FILL_0_BUFX4_131 ( );
FILL FILL_1_BUFX4_131 ( );
FILL FILL_2_BUFX4_131 ( );
FILL FILL_0_OAI21X1_481 ( );
FILL FILL_1_OAI21X1_481 ( );
FILL FILL_0_BUFX2_593 ( );
FILL FILL_1_BUFX2_593 ( );
FILL FILL_0_BUFX2_510 ( );
FILL FILL_1_BUFX2_510 ( );
FILL FILL_0_BUFX2_509 ( );
FILL FILL_1_BUFX2_509 ( );
FILL FILL_0_NAND2X1_245 ( );
FILL FILL_1_NAND2X1_245 ( );
FILL FILL_0_CLKBUF1_48 ( );
FILL FILL_1_CLKBUF1_48 ( );
FILL FILL_2_CLKBUF1_48 ( );
FILL FILL_3_CLKBUF1_48 ( );
FILL FILL_4_CLKBUF1_48 ( );
FILL FILL_0_NAND2X1_106 ( );
FILL FILL_1_NAND2X1_106 ( );
FILL FILL_0_OAI21X1_362 ( );
FILL FILL_1_OAI21X1_362 ( );
FILL FILL_0_INVX1_2 ( );
FILL FILL_0_DFFPOSX1_453 ( );
FILL FILL_1_DFFPOSX1_453 ( );
FILL FILL_2_DFFPOSX1_453 ( );
FILL FILL_3_DFFPOSX1_453 ( );
FILL FILL_4_DFFPOSX1_453 ( );
FILL FILL_5_DFFPOSX1_453 ( );
FILL FILL_6_DFFPOSX1_453 ( );
FILL FILL_0_OAI21X1_450 ( );
FILL FILL_1_OAI21X1_450 ( );
FILL FILL_0_NAND2X1_207 ( );
FILL FILL_1_NAND2X1_207 ( );
FILL FILL_0_NAND2X1_133 ( );
FILL FILL_1_NAND2X1_133 ( );
FILL FILL_0_INVX1_15 ( );
FILL FILL_0_OAI21X1_449 ( );
FILL FILL_1_OAI21X1_449 ( );
FILL FILL_0_OAI21X1_453 ( );
FILL FILL_1_OAI21X1_453 ( );
FILL FILL_0_NAND2X1_208 ( );
FILL FILL_0_OAI21X1_560 ( );
FILL FILL_1_OAI21X1_560 ( );
FILL FILL_0_DFFPOSX1_506 ( );
FILL FILL_1_DFFPOSX1_506 ( );
FILL FILL_2_DFFPOSX1_506 ( );
FILL FILL_3_DFFPOSX1_506 ( );
FILL FILL_4_DFFPOSX1_506 ( );
FILL FILL_5_DFFPOSX1_506 ( );
FILL FILL_0_NAND2X1_180 ( );
FILL FILL_1_NAND2X1_180 ( );
FILL FILL_0_BUFX2_465 ( );
FILL FILL_1_BUFX2_465 ( );
FILL FILL_0_BUFX4_236 ( );
FILL FILL_1_BUFX4_236 ( );
FILL FILL_0_BUFX4_337 ( );
FILL FILL_1_BUFX4_337 ( );
FILL FILL_2_BUFX4_337 ( );
FILL FILL_0_OAI21X1_433 ( );
FILL FILL_1_OAI21X1_433 ( );
FILL FILL_0_XNOR2X1_8 ( );
FILL FILL_1_XNOR2X1_8 ( );
FILL FILL_2_XNOR2X1_8 ( );
FILL FILL_3_XNOR2X1_8 ( );
FILL FILL_0_OAI21X1_431 ( );
FILL FILL_1_OAI21X1_431 ( );
FILL FILL_0_INVX2_20 ( );
FILL FILL_0_BUFX2_413 ( );
FILL FILL_1_BUFX2_413 ( );
FILL FILL_0_XNOR2X1_31 ( );
FILL FILL_1_XNOR2X1_31 ( );
FILL FILL_2_XNOR2X1_31 ( );
FILL FILL_3_XNOR2X1_31 ( );
FILL FILL_0_NAND2X1_193 ( );
FILL FILL_1_NAND2X1_193 ( );
FILL FILL_0_BUFX4_383 ( );
FILL FILL_1_BUFX4_383 ( );
FILL FILL_0_BUFX2_553 ( );
FILL FILL_0_BUFX2_417 ( );
FILL FILL_0_BUFX4_214 ( );
FILL FILL_1_BUFX4_214 ( );
FILL FILL_0_DFFPOSX1_448 ( );
FILL FILL_1_DFFPOSX1_448 ( );
FILL FILL_2_DFFPOSX1_448 ( );
FILL FILL_3_DFFPOSX1_448 ( );
FILL FILL_4_DFFPOSX1_448 ( );
FILL FILL_5_DFFPOSX1_448 ( );
FILL FILL_0_BUFX2_541 ( );
FILL FILL_1_BUFX2_541 ( );
FILL FILL_0_DFFPOSX1_344 ( );
FILL FILL_1_DFFPOSX1_344 ( );
FILL FILL_2_DFFPOSX1_344 ( );
FILL FILL_3_DFFPOSX1_344 ( );
FILL FILL_4_DFFPOSX1_344 ( );
FILL FILL_5_DFFPOSX1_344 ( );
FILL FILL_0_OAI21X1_1814 ( );
FILL FILL_1_OAI21X1_1814 ( );
FILL FILL_0_BUFX2_415 ( );
FILL FILL_0_BUFX2_1006 ( );
FILL FILL_1_BUFX2_1006 ( );
FILL FILL_0_BUFX2_602 ( );
FILL FILL_0_BUFX2_962 ( );
FILL FILL_1_BUFX2_962 ( );
FILL FILL_0_BUFX2_15 ( );
FILL FILL_1_BUFX2_15 ( );
FILL FILL_0_BUFX2_610 ( );
FILL FILL_0_CLKBUF1_52 ( );
FILL FILL_1_CLKBUF1_52 ( );
FILL FILL_2_CLKBUF1_52 ( );
FILL FILL_3_CLKBUF1_52 ( );
FILL FILL_4_CLKBUF1_52 ( );
FILL FILL_0_DFFPOSX1_830 ( );
FILL FILL_1_DFFPOSX1_830 ( );
FILL FILL_2_DFFPOSX1_830 ( );
FILL FILL_3_DFFPOSX1_830 ( );
FILL FILL_4_DFFPOSX1_830 ( );
FILL FILL_5_DFFPOSX1_830 ( );
FILL FILL_6_DFFPOSX1_830 ( );
FILL FILL_0_NAND2X1_426 ( );
FILL FILL_1_NAND2X1_426 ( );
FILL FILL_0_NAND2X1_504 ( );
FILL FILL_1_NAND2X1_504 ( );
FILL FILL_0_DFFPOSX1_831 ( );
FILL FILL_1_DFFPOSX1_831 ( );
FILL FILL_2_DFFPOSX1_831 ( );
FILL FILL_3_DFFPOSX1_831 ( );
FILL FILL_4_DFFPOSX1_831 ( );
FILL FILL_5_DFFPOSX1_831 ( );
FILL FILL_0_OAI21X1_1142 ( );
FILL FILL_1_OAI21X1_1142 ( );
FILL FILL_2_OAI21X1_1142 ( );
FILL FILL_0_BUFX4_228 ( );
FILL FILL_1_BUFX4_228 ( );
FILL FILL_2_BUFX4_228 ( );
FILL FILL_0_BUFX4_192 ( );
FILL FILL_1_BUFX4_192 ( );
FILL FILL_0_NAND2X1_508 ( );
FILL FILL_0_CLKBUF1_51 ( );
FILL FILL_1_CLKBUF1_51 ( );
FILL FILL_2_CLKBUF1_51 ( );
FILL FILL_3_CLKBUF1_51 ( );
FILL FILL_4_CLKBUF1_51 ( );
FILL FILL_0_OAI21X1_191 ( );
FILL FILL_1_OAI21X1_191 ( );
FILL FILL_0_OAI21X1_190 ( );
FILL FILL_1_OAI21X1_190 ( );
FILL FILL_0_NAND2X1_503 ( );
FILL FILL_0_OAI21X1_130 ( );
FILL FILL_1_OAI21X1_130 ( );
FILL FILL_0_CLKBUF1_62 ( );
FILL FILL_1_CLKBUF1_62 ( );
FILL FILL_2_CLKBUF1_62 ( );
FILL FILL_3_CLKBUF1_62 ( );
FILL FILL_0_BUFX2_226 ( );
FILL FILL_1_BUFX2_226 ( );
FILL FILL_0_BUFX2_75 ( );
FILL FILL_1_BUFX2_75 ( );
FILL FILL_0_BUFX2_32 ( );
FILL FILL_1_BUFX2_32 ( );
FILL FILL_0_OAI21X1_1314 ( );
FILL FILL_1_OAI21X1_1314 ( );
FILL FILL_0_OAI21X1_1315 ( );
FILL FILL_1_OAI21X1_1315 ( );
FILL FILL_0_XNOR2X1_84 ( );
FILL FILL_1_XNOR2X1_84 ( );
FILL FILL_2_XNOR2X1_84 ( );
FILL FILL_3_XNOR2X1_84 ( );
FILL FILL_0_XNOR2X1_71 ( );
FILL FILL_1_XNOR2X1_71 ( );
FILL FILL_2_XNOR2X1_71 ( );
FILL FILL_3_XNOR2X1_71 ( );
FILL FILL_0_OAI21X1_1077 ( );
FILL FILL_1_OAI21X1_1077 ( );
FILL FILL_0_NAND3X1_43 ( );
FILL FILL_1_NAND3X1_43 ( );
FILL FILL_0_NOR2X1_158 ( );
FILL FILL_0_XNOR2X1_70 ( );
FILL FILL_1_XNOR2X1_70 ( );
FILL FILL_2_XNOR2X1_70 ( );
FILL FILL_0_OAI21X1_1317 ( );
FILL FILL_1_OAI21X1_1317 ( );
FILL FILL_0_OAI21X1_1318 ( );
FILL FILL_1_OAI21X1_1318 ( );
FILL FILL_2_OAI21X1_1318 ( );
FILL FILL_0_OAI21X1_1319 ( );
FILL FILL_1_OAI21X1_1319 ( );
FILL FILL_0_OAI21X1_1166 ( );
FILL FILL_1_OAI21X1_1166 ( );
FILL FILL_0_OAI21X1_1316 ( );
FILL FILL_1_OAI21X1_1316 ( );
FILL FILL_0_OAI21X1_1488 ( );
FILL FILL_1_OAI21X1_1488 ( );
FILL FILL_0_DFFPOSX1_912 ( );
FILL FILL_1_DFFPOSX1_912 ( );
FILL FILL_2_DFFPOSX1_912 ( );
FILL FILL_3_DFFPOSX1_912 ( );
FILL FILL_4_DFFPOSX1_912 ( );
FILL FILL_5_DFFPOSX1_912 ( );
FILL FILL_0_BUFX2_164 ( );
FILL FILL_1_BUFX2_164 ( );
FILL FILL_0_BUFX4_364 ( );
FILL FILL_1_BUFX4_364 ( );
FILL FILL_0_OAI21X1_1815 ( );
FILL FILL_1_OAI21X1_1815 ( );
FILL FILL_0_DFFPOSX1_795 ( );
FILL FILL_1_DFFPOSX1_795 ( );
FILL FILL_2_DFFPOSX1_795 ( );
FILL FILL_3_DFFPOSX1_795 ( );
FILL FILL_4_DFFPOSX1_795 ( );
FILL FILL_5_DFFPOSX1_795 ( );
FILL FILL_0_OAI21X1_37 ( );
FILL FILL_1_OAI21X1_37 ( );
FILL FILL_0_BUFX2_113 ( );
FILL FILL_0_BUFX4_68 ( );
FILL FILL_1_BUFX4_68 ( );
FILL FILL_0_BUFX2_183 ( );
FILL FILL_0_CLKBUF1_71 ( );
FILL FILL_1_CLKBUF1_71 ( );
FILL FILL_2_CLKBUF1_71 ( );
FILL FILL_3_CLKBUF1_71 ( );
FILL FILL_4_CLKBUF1_71 ( );
FILL FILL_0_DFFPOSX1_863 ( );
FILL FILL_1_DFFPOSX1_863 ( );
FILL FILL_2_DFFPOSX1_863 ( );
FILL FILL_3_DFFPOSX1_863 ( );
FILL FILL_4_DFFPOSX1_863 ( );
FILL FILL_5_DFFPOSX1_863 ( );
FILL FILL_6_DFFPOSX1_863 ( );
FILL FILL_0_NAND2X1_577 ( );
FILL FILL_1_NAND2X1_577 ( );
FILL FILL_0_BUFX2_116 ( );
FILL FILL_0_NAND2X1_576 ( );
FILL FILL_0_OAI21X1_1549 ( );
FILL FILL_1_OAI21X1_1549 ( );
FILL FILL_0_DFFPOSX1_990 ( );
FILL FILL_1_DFFPOSX1_990 ( );
FILL FILL_2_DFFPOSX1_990 ( );
FILL FILL_3_DFFPOSX1_990 ( );
FILL FILL_4_DFFPOSX1_990 ( );
FILL FILL_5_DFFPOSX1_990 ( );
FILL FILL_0_OAI21X1_1548 ( );
FILL FILL_1_OAI21X1_1548 ( );
FILL FILL_0_BUFX2_259 ( );
FILL FILL_0_OAI21X1_1090 ( );
FILL FILL_1_OAI21X1_1090 ( );
FILL FILL_0_NAND2X1_456 ( );
FILL FILL_0_DFFPOSX1_798 ( );
FILL FILL_1_DFFPOSX1_798 ( );
FILL FILL_2_DFFPOSX1_798 ( );
FILL FILL_3_DFFPOSX1_798 ( );
FILL FILL_4_DFFPOSX1_798 ( );
FILL FILL_5_DFFPOSX1_798 ( );
FILL FILL_6_DFFPOSX1_798 ( );
FILL FILL_0_OAI21X1_1550 ( );
FILL FILL_1_OAI21X1_1550 ( );
FILL FILL_0_BUFX4_338 ( );
FILL FILL_1_BUFX4_338 ( );
FILL FILL_0_BUFX2_181 ( );
FILL FILL_0_BUFX2_244 ( );
FILL FILL_1_BUFX2_244 ( );
FILL FILL_0_OAI21X1_154 ( );
FILL FILL_1_OAI21X1_154 ( );
FILL FILL_0_OAI21X1_155 ( );
FILL FILL_1_OAI21X1_155 ( );
FILL FILL_2_OAI21X1_155 ( );
FILL FILL_0_NAND2X1_655 ( );
FILL FILL_0_BUFX4_154 ( );
FILL FILL_1_BUFX4_154 ( );
FILL FILL_0_DFFPOSX1_269 ( );
FILL FILL_1_DFFPOSX1_269 ( );
FILL FILL_2_DFFPOSX1_269 ( );
FILL FILL_3_DFFPOSX1_269 ( );
FILL FILL_4_DFFPOSX1_269 ( );
FILL FILL_5_DFFPOSX1_269 ( );
FILL FILL_6_DFFPOSX1_269 ( );
FILL FILL_0_OAI21X1_946 ( );
FILL FILL_1_OAI21X1_946 ( );
FILL FILL_0_BUFX2_353 ( );
FILL FILL_1_BUFX2_353 ( );
FILL FILL_0_OAI21X1_947 ( );
FILL FILL_1_OAI21X1_947 ( );
FILL FILL_0_DFFPOSX1_699 ( );
FILL FILL_1_DFFPOSX1_699 ( );
FILL FILL_2_DFFPOSX1_699 ( );
FILL FILL_3_DFFPOSX1_699 ( );
FILL FILL_4_DFFPOSX1_699 ( );
FILL FILL_5_DFFPOSX1_699 ( );
FILL FILL_0_BUFX2_351 ( );
FILL FILL_1_BUFX2_351 ( );
FILL FILL_0_INVX1_159 ( );
FILL FILL_0_BUFX2_741 ( );
FILL FILL_1_BUFX2_741 ( );
FILL FILL_0_DFFPOSX1_74 ( );
FILL FILL_1_DFFPOSX1_74 ( );
FILL FILL_2_DFFPOSX1_74 ( );
FILL FILL_3_DFFPOSX1_74 ( );
FILL FILL_4_DFFPOSX1_74 ( );
FILL FILL_5_DFFPOSX1_74 ( );
FILL FILL_6_DFFPOSX1_74 ( );
FILL FILL_0_OAI21X1_1723 ( );
FILL FILL_1_OAI21X1_1723 ( );
FILL FILL_2_OAI21X1_1723 ( );
FILL FILL_0_OAI21X1_1722 ( );
FILL FILL_1_OAI21X1_1722 ( );
FILL FILL_0_DFFPOSX1_730 ( );
FILL FILL_1_DFFPOSX1_730 ( );
FILL FILL_2_DFFPOSX1_730 ( );
FILL FILL_3_DFFPOSX1_730 ( );
FILL FILL_4_DFFPOSX1_730 ( );
FILL FILL_5_DFFPOSX1_730 ( );
FILL FILL_0_OAI21X1_1009 ( );
FILL FILL_1_OAI21X1_1009 ( );
FILL FILL_0_OAI21X1_136 ( );
FILL FILL_1_OAI21X1_136 ( );
FILL FILL_2_OAI21X1_136 ( );
FILL FILL_0_OAI21X1_137 ( );
FILL FILL_1_OAI21X1_137 ( );
FILL FILL_0_OAI21X1_264 ( );
FILL FILL_1_OAI21X1_264 ( );
FILL FILL_0_OAI21X1_265 ( );
FILL FILL_1_OAI21X1_265 ( );
FILL FILL_0_DFFPOSX1_324 ( );
FILL FILL_1_DFFPOSX1_324 ( );
FILL FILL_2_DFFPOSX1_324 ( );
FILL FILL_3_DFFPOSX1_324 ( );
FILL FILL_4_DFFPOSX1_324 ( );
FILL FILL_5_DFFPOSX1_324 ( );
FILL FILL_0_DFFPOSX1_132 ( );
FILL FILL_1_DFFPOSX1_132 ( );
FILL FILL_2_DFFPOSX1_132 ( );
FILL FILL_3_DFFPOSX1_132 ( );
FILL FILL_4_DFFPOSX1_132 ( );
FILL FILL_5_DFFPOSX1_132 ( );
FILL FILL_0_BUFX2_522 ( );
FILL FILL_1_BUFX2_522 ( );
FILL FILL_0_BUFX2_738 ( );
FILL FILL_1_BUFX2_738 ( );
FILL FILL_0_BUFX4_320 ( );
FILL FILL_1_BUFX4_320 ( );
FILL FILL_0_DFFPOSX1_488 ( );
FILL FILL_1_DFFPOSX1_488 ( );
FILL FILL_2_DFFPOSX1_488 ( );
FILL FILL_3_DFFPOSX1_488 ( );
FILL FILL_4_DFFPOSX1_488 ( );
FILL FILL_5_DFFPOSX1_488 ( );
FILL FILL_6_DFFPOSX1_488 ( );
FILL FILL_0_OAI21X1_511 ( );
FILL FILL_1_OAI21X1_511 ( );
FILL FILL_0_OAI21X1_512 ( );
FILL FILL_1_OAI21X1_512 ( );
FILL FILL_0_INVX2_12 ( );
FILL FILL_0_OAI21X1_344 ( );
FILL FILL_1_OAI21X1_344 ( );
FILL FILL_2_OAI21X1_344 ( );
FILL FILL_0_DFFPOSX1_372 ( );
FILL FILL_1_DFFPOSX1_372 ( );
FILL FILL_2_DFFPOSX1_372 ( );
FILL FILL_3_DFFPOSX1_372 ( );
FILL FILL_4_DFFPOSX1_372 ( );
FILL FILL_5_DFFPOSX1_372 ( );
FILL FILL_0_BUFX2_397 ( );
FILL FILL_0_INVX4_2 ( );
FILL FILL_0_BUFX4_163 ( );
FILL FILL_1_BUFX4_163 ( );
FILL FILL_2_BUFX4_163 ( );
FILL FILL_0_BUFX2_577 ( );
FILL FILL_1_BUFX2_577 ( );
FILL FILL_0_OAI21X1_516 ( );
FILL FILL_1_OAI21X1_516 ( );
FILL FILL_2_OAI21X1_516 ( );
FILL FILL_0_CLKBUF1_75 ( );
FILL FILL_1_CLKBUF1_75 ( );
FILL FILL_2_CLKBUF1_75 ( );
FILL FILL_3_CLKBUF1_75 ( );
FILL FILL_0_NAND2X1_271 ( );
FILL FILL_1_NAND2X1_271 ( );
FILL FILL_0_DFFPOSX1_562 ( );
FILL FILL_1_DFFPOSX1_562 ( );
FILL FILL_2_DFFPOSX1_562 ( );
FILL FILL_3_DFFPOSX1_562 ( );
FILL FILL_4_DFFPOSX1_562 ( );
FILL FILL_5_DFFPOSX1_562 ( );
FILL FILL_6_DFFPOSX1_562 ( );
FILL FILL_0_OAI21X1_700 ( );
FILL FILL_1_OAI21X1_700 ( );
FILL FILL_0_INVX4_6 ( );
FILL FILL_1_INVX4_6 ( );
FILL FILL_0_OAI21X1_686 ( );
FILL FILL_1_OAI21X1_686 ( );
FILL FILL_0_OAI21X1_688 ( );
FILL FILL_1_OAI21X1_688 ( );
FILL FILL_0_INVX4_5 ( );
FILL FILL_1_INVX4_5 ( );
FILL FILL_0_DFFPOSX1_558 ( );
FILL FILL_1_DFFPOSX1_558 ( );
FILL FILL_2_DFFPOSX1_558 ( );
FILL FILL_3_DFFPOSX1_558 ( );
FILL FILL_4_DFFPOSX1_558 ( );
FILL FILL_5_DFFPOSX1_558 ( );
FILL FILL_0_NAND2X1_311 ( );
FILL FILL_1_NAND2X1_311 ( );
FILL FILL_0_BUFX2_529 ( );
FILL FILL_0_BUFX2_525 ( );
FILL FILL_1_BUFX2_525 ( );
FILL FILL_0_INVX4_4 ( );
FILL FILL_1_INVX4_4 ( );
FILL FILL_0_XNOR2X1_20 ( );
FILL FILL_1_XNOR2X1_20 ( );
FILL FILL_2_XNOR2X1_20 ( );
FILL FILL_3_XNOR2X1_20 ( );
FILL FILL_0_AND2X2_9 ( );
FILL FILL_1_AND2X2_9 ( );
FILL FILL_0_BUFX4_182 ( );
FILL FILL_1_BUFX4_182 ( );
FILL FILL_0_DFFPOSX1_464 ( );
FILL FILL_1_DFFPOSX1_464 ( );
FILL FILL_2_DFFPOSX1_464 ( );
FILL FILL_3_DFFPOSX1_464 ( );
FILL FILL_4_DFFPOSX1_464 ( );
FILL FILL_5_DFFPOSX1_464 ( );
FILL FILL_6_DFFPOSX1_464 ( );
FILL FILL_0_DFFPOSX1_549 ( );
FILL FILL_1_DFFPOSX1_549 ( );
FILL FILL_2_DFFPOSX1_549 ( );
FILL FILL_3_DFFPOSX1_549 ( );
FILL FILL_4_DFFPOSX1_549 ( );
FILL FILL_5_DFFPOSX1_549 ( );
FILL FILL_6_DFFPOSX1_549 ( );
FILL FILL_0_DFFPOSX1_517 ( );
FILL FILL_1_DFFPOSX1_517 ( );
FILL FILL_2_DFFPOSX1_517 ( );
FILL FILL_3_DFFPOSX1_517 ( );
FILL FILL_4_DFFPOSX1_517 ( );
FILL FILL_5_DFFPOSX1_517 ( );
FILL FILL_0_DFFPOSX1_518 ( );
FILL FILL_1_DFFPOSX1_518 ( );
FILL FILL_2_DFFPOSX1_518 ( );
FILL FILL_3_DFFPOSX1_518 ( );
FILL FILL_4_DFFPOSX1_518 ( );
FILL FILL_5_DFFPOSX1_518 ( );
FILL FILL_6_DFFPOSX1_518 ( );
FILL FILL_0_DFFPOSX1_390 ( );
FILL FILL_1_DFFPOSX1_390 ( );
FILL FILL_2_DFFPOSX1_390 ( );
FILL FILL_3_DFFPOSX1_390 ( );
FILL FILL_4_DFFPOSX1_390 ( );
FILL FILL_5_DFFPOSX1_390 ( );
FILL FILL_6_DFFPOSX1_390 ( );
FILL FILL_0_DFFPOSX1_454 ( );
FILL FILL_1_DFFPOSX1_454 ( );
FILL FILL_2_DFFPOSX1_454 ( );
FILL FILL_3_DFFPOSX1_454 ( );
FILL FILL_4_DFFPOSX1_454 ( );
FILL FILL_5_DFFPOSX1_454 ( );
FILL FILL_0_XNOR2X1_13 ( );
FILL FILL_1_XNOR2X1_13 ( );
FILL FILL_2_XNOR2X1_13 ( );
FILL FILL_3_XNOR2X1_13 ( );
FILL FILL_0_OAI21X1_452 ( );
FILL FILL_1_OAI21X1_452 ( );
FILL FILL_0_XNOR2X1_14 ( );
FILL FILL_1_XNOR2X1_14 ( );
FILL FILL_2_XNOR2X1_14 ( );
FILL FILL_3_XNOR2X1_14 ( );
FILL FILL_0_DFFPOSX1_455 ( );
FILL FILL_1_DFFPOSX1_455 ( );
FILL FILL_2_DFFPOSX1_455 ( );
FILL FILL_3_DFFPOSX1_455 ( );
FILL FILL_4_DFFPOSX1_455 ( );
FILL FILL_5_DFFPOSX1_455 ( );
FILL FILL_6_DFFPOSX1_455 ( );
FILL FILL_0_OAI21X1_561 ( );
FILL FILL_1_OAI21X1_561 ( );
FILL FILL_0_DFFPOSX1_441 ( );
FILL FILL_1_DFFPOSX1_441 ( );
FILL FILL_2_DFFPOSX1_441 ( );
FILL FILL_3_DFFPOSX1_441 ( );
FILL FILL_4_DFFPOSX1_441 ( );
FILL FILL_5_DFFPOSX1_441 ( );
FILL FILL_0_OAI21X1_432 ( );
FILL FILL_1_OAI21X1_432 ( );
FILL FILL_0_XNOR2X1_29 ( );
FILL FILL_1_XNOR2X1_29 ( );
FILL FILL_2_XNOR2X1_29 ( );
FILL FILL_3_XNOR2X1_29 ( );
FILL FILL_0_NOR2X1_66 ( );
FILL FILL_1_NOR2X1_66 ( );
FILL FILL_0_MUX2X1_1 ( );
FILL FILL_1_MUX2X1_1 ( );
FILL FILL_2_MUX2X1_1 ( );
FILL FILL_0_INVX4_8 ( );
FILL FILL_0_XNOR2X1_30 ( );
FILL FILL_1_XNOR2X1_30 ( );
FILL FILL_2_XNOR2X1_30 ( );
FILL FILL_0_NAND2X1_280 ( );
FILL FILL_0_DFFPOSX1_447 ( );
FILL FILL_1_DFFPOSX1_447 ( );
FILL FILL_2_DFFPOSX1_447 ( );
FILL FILL_3_DFFPOSX1_447 ( );
FILL FILL_4_DFFPOSX1_447 ( );
FILL FILL_5_DFFPOSX1_447 ( );
FILL FILL_6_DFFPOSX1_447 ( );
FILL FILL_0_OAI21X1_601 ( );
FILL FILL_1_OAI21X1_601 ( );
FILL FILL_0_OAI21X1_443 ( );
FILL FILL_1_OAI21X1_443 ( );
FILL FILL_0_NAND2X1_197 ( );
FILL FILL_0_NAND2X1_188 ( );
FILL FILL_0_DFFPOSX1_444 ( );
FILL FILL_1_DFFPOSX1_444 ( );
FILL FILL_2_DFFPOSX1_444 ( );
FILL FILL_3_DFFPOSX1_444 ( );
FILL FILL_4_DFFPOSX1_444 ( );
FILL FILL_5_DFFPOSX1_444 ( );
FILL FILL_0_OAI21X1_305 ( );
FILL FILL_1_OAI21X1_305 ( );
FILL FILL_2_OAI21X1_305 ( );
FILL FILL_0_OAI21X1_176 ( );
FILL FILL_1_OAI21X1_176 ( );
FILL FILL_0_OAI21X1_177 ( );
FILL FILL_1_OAI21X1_177 ( );
FILL FILL_0_NAND2X1_103 ( );
FILL FILL_0_DFFPOSX1_280 ( );
FILL FILL_1_DFFPOSX1_280 ( );
FILL FILL_2_DFFPOSX1_280 ( );
FILL FILL_3_DFFPOSX1_280 ( );
FILL FILL_4_DFFPOSX1_280 ( );
FILL FILL_5_DFFPOSX1_280 ( );
FILL FILL_6_DFFPOSX1_280 ( );
FILL FILL_0_CLKBUF1_2 ( );
FILL FILL_1_CLKBUF1_2 ( );
FILL FILL_2_CLKBUF1_2 ( );
FILL FILL_3_CLKBUF1_2 ( );
FILL FILL_4_CLKBUF1_2 ( );
FILL FILL_0_DFFPOSX1_288 ( );
FILL FILL_1_DFFPOSX1_288 ( );
FILL FILL_2_DFFPOSX1_288 ( );
FILL FILL_3_DFFPOSX1_288 ( );
FILL FILL_4_DFFPOSX1_288 ( );
FILL FILL_5_DFFPOSX1_288 ( );
FILL FILL_0_OAI21X1_192 ( );
FILL FILL_1_OAI21X1_192 ( );
FILL FILL_0_OAI21X1_193 ( );
FILL FILL_1_OAI21X1_193 ( );
FILL FILL_0_BUFX2_971 ( );
FILL FILL_0_OAI21X1_1134 ( );
FILL FILL_1_OAI21X1_1134 ( );
FILL FILL_0_DFFPOSX1_768 ( );
FILL FILL_1_DFFPOSX1_768 ( );
FILL FILL_2_DFFPOSX1_768 ( );
FILL FILL_3_DFFPOSX1_768 ( );
FILL FILL_4_DFFPOSX1_768 ( );
FILL FILL_5_DFFPOSX1_768 ( );
FILL FILL_0_OAI21X1_1141 ( );
FILL FILL_1_OAI21X1_1141 ( );
FILL FILL_0_DFFPOSX1_827 ( );
FILL FILL_1_DFFPOSX1_827 ( );
FILL FILL_2_DFFPOSX1_827 ( );
FILL FILL_3_DFFPOSX1_827 ( );
FILL FILL_4_DFFPOSX1_827 ( );
FILL FILL_5_DFFPOSX1_827 ( );
FILL FILL_0_OAI21X1_1138 ( );
FILL FILL_1_OAI21X1_1138 ( );
FILL FILL_2_OAI21X1_1138 ( );
FILL FILL_0_NAND2X1_510 ( );
FILL FILL_0_BUFX4_186 ( );
FILL FILL_1_BUFX4_186 ( );
FILL FILL_0_DFFPOSX1_829 ( );
FILL FILL_1_DFFPOSX1_829 ( );
FILL FILL_2_DFFPOSX1_829 ( );
FILL FILL_3_DFFPOSX1_829 ( );
FILL FILL_4_DFFPOSX1_829 ( );
FILL FILL_5_DFFPOSX1_829 ( );
FILL FILL_0_OAI21X1_1500 ( );
FILL FILL_1_OAI21X1_1500 ( );
FILL FILL_0_OAI21X1_1501 ( );
FILL FILL_1_OAI21X1_1501 ( );
FILL FILL_0_DFFPOSX1_826 ( );
FILL FILL_1_DFFPOSX1_826 ( );
FILL FILL_2_DFFPOSX1_826 ( );
FILL FILL_3_DFFPOSX1_826 ( );
FILL FILL_4_DFFPOSX1_826 ( );
FILL FILL_5_DFFPOSX1_826 ( );
FILL FILL_6_DFFPOSX1_826 ( );
FILL FILL_0_OAI21X1_319 ( );
FILL FILL_1_OAI21X1_319 ( );
FILL FILL_0_OAI21X1_318 ( );
FILL FILL_1_OAI21X1_318 ( );
FILL FILL_2_OAI21X1_318 ( );
FILL FILL_0_BUFX2_209 ( );
FILL FILL_0_OAI21X1_1308 ( );
FILL FILL_1_OAI21X1_1308 ( );
FILL FILL_0_DFFPOSX1_908 ( );
FILL FILL_1_DFFPOSX1_908 ( );
FILL FILL_2_DFFPOSX1_908 ( );
FILL FILL_3_DFFPOSX1_908 ( );
FILL FILL_4_DFFPOSX1_908 ( );
FILL FILL_5_DFFPOSX1_908 ( );
FILL FILL_6_DFFPOSX1_908 ( );
FILL FILL_0_NAND2X1_543 ( );
FILL FILL_0_DFFPOSX1_911 ( );
FILL FILL_1_DFFPOSX1_911 ( );
FILL FILL_2_DFFPOSX1_911 ( );
FILL FILL_3_DFFPOSX1_911 ( );
FILL FILL_4_DFFPOSX1_911 ( );
FILL FILL_5_DFFPOSX1_911 ( );
FILL FILL_0_XNOR2X1_68 ( );
FILL FILL_1_XNOR2X1_68 ( );
FILL FILL_2_XNOR2X1_68 ( );
FILL FILL_3_XNOR2X1_68 ( );
FILL FILL_0_NOR2X1_157 ( );
FILL FILL_1_NOR2X1_157 ( );
FILL FILL_0_XNOR2X1_67 ( );
FILL FILL_1_XNOR2X1_67 ( );
FILL FILL_2_XNOR2X1_67 ( );
FILL FILL_3_XNOR2X1_67 ( );
FILL FILL_0_BUFX4_226 ( );
FILL FILL_1_BUFX4_226 ( );
FILL FILL_0_XNOR2X1_101 ( );
FILL FILL_1_XNOR2X1_101 ( );
FILL FILL_2_XNOR2X1_101 ( );
FILL FILL_3_XNOR2X1_101 ( );
FILL FILL_0_OAI21X1_1165 ( );
FILL FILL_1_OAI21X1_1165 ( );
FILL FILL_0_NAND2X1_547 ( );
FILL FILL_1_NAND2X1_547 ( );
FILL FILL_0_OAI21X1_1502 ( );
FILL FILL_1_OAI21X1_1502 ( );
FILL FILL_0_OAI21X1_1503 ( );
FILL FILL_1_OAI21X1_1503 ( );
FILL FILL_2_OAI21X1_1503 ( );
FILL FILL_0_DFFPOSX1_907 ( );
FILL FILL_1_DFFPOSX1_907 ( );
FILL FILL_2_DFFPOSX1_907 ( );
FILL FILL_3_DFFPOSX1_907 ( );
FILL FILL_4_DFFPOSX1_907 ( );
FILL FILL_5_DFFPOSX1_907 ( );
FILL FILL_0_OAI21X1_1087 ( );
FILL FILL_1_OAI21X1_1087 ( );
FILL FILL_0_NAND2X1_453 ( );
FILL FILL_1_NAND2X1_453 ( );
FILL FILL_0_DFFPOSX1_193 ( );
FILL FILL_1_DFFPOSX1_193 ( );
FILL FILL_2_DFFPOSX1_193 ( );
FILL FILL_3_DFFPOSX1_193 ( );
FILL FILL_4_DFFPOSX1_193 ( );
FILL FILL_5_DFFPOSX1_193 ( );
FILL FILL_6_DFFPOSX1_193 ( );
FILL FILL_0_OAI21X1_1355 ( );
FILL FILL_1_OAI21X1_1355 ( );
FILL FILL_0_CLKBUF1_76 ( );
FILL FILL_1_CLKBUF1_76 ( );
FILL FILL_2_CLKBUF1_76 ( );
FILL FILL_3_CLKBUF1_76 ( );
FILL FILL_4_CLKBUF1_76 ( );
FILL FILL_0_OAI21X1_1191 ( );
FILL FILL_1_OAI21X1_1191 ( );
FILL FILL_0_OAI21X1_1189 ( );
FILL FILL_1_OAI21X1_1189 ( );
FILL FILL_0_BUFX4_201 ( );
FILL FILL_1_BUFX4_201 ( );
FILL FILL_0_NOR2X1_170 ( );
FILL FILL_1_NOR2X1_170 ( );
FILL FILL_0_DFFPOSX1_614 ( );
FILL FILL_1_DFFPOSX1_614 ( );
FILL FILL_2_DFFPOSX1_614 ( );
FILL FILL_3_DFFPOSX1_614 ( );
FILL FILL_4_DFFPOSX1_614 ( );
FILL FILL_5_DFFPOSX1_614 ( );
FILL FILL_6_DFFPOSX1_614 ( );
FILL FILL_0_INVX2_88 ( );
FILL FILL_0_BUFX4_73 ( );
FILL FILL_1_BUFX4_73 ( );
FILL FILL_0_DFFPOSX1_862 ( );
FILL FILL_1_DFFPOSX1_862 ( );
FILL FILL_2_DFFPOSX1_862 ( );
FILL FILL_3_DFFPOSX1_862 ( );
FILL FILL_4_DFFPOSX1_862 ( );
FILL FILL_5_DFFPOSX1_862 ( );
FILL FILL_0_OAI21X1_1361 ( );
FILL FILL_1_OAI21X1_1361 ( );
FILL FILL_0_DFFPOSX1_928 ( );
FILL FILL_1_DFFPOSX1_928 ( );
FILL FILL_2_DFFPOSX1_928 ( );
FILL FILL_3_DFFPOSX1_928 ( );
FILL FILL_4_DFFPOSX1_928 ( );
FILL FILL_5_DFFPOSX1_928 ( );
FILL FILL_6_DFFPOSX1_928 ( );
FILL FILL_0_BUFX4_374 ( );
FILL FILL_1_BUFX4_374 ( );
FILL FILL_0_BUFX2_179 ( );
FILL FILL_1_BUFX2_179 ( );
FILL FILL_0_CLKBUF1_37 ( );
FILL FILL_1_CLKBUF1_37 ( );
FILL FILL_2_CLKBUF1_37 ( );
FILL FILL_3_CLKBUF1_37 ( );
FILL FILL_4_CLKBUF1_37 ( );
FILL FILL_0_OAI21X1_921 ( );
FILL FILL_1_OAI21X1_921 ( );
FILL FILL_0_DFFPOSX1_686 ( );
FILL FILL_1_DFFPOSX1_686 ( );
FILL FILL_2_DFFPOSX1_686 ( );
FILL FILL_3_DFFPOSX1_686 ( );
FILL FILL_4_DFFPOSX1_686 ( );
FILL FILL_5_DFFPOSX1_686 ( );
FILL FILL_0_OAI21X1_917 ( );
FILL FILL_1_OAI21X1_917 ( );
FILL FILL_0_DFFPOSX1_684 ( );
FILL FILL_1_DFFPOSX1_684 ( );
FILL FILL_2_DFFPOSX1_684 ( );
FILL FILL_3_DFFPOSX1_684 ( );
FILL FILL_4_DFFPOSX1_684 ( );
FILL FILL_5_DFFPOSX1_684 ( );
FILL FILL_0_INVX1_172 ( );
FILL FILL_0_BUFX2_676 ( );
FILL FILL_1_BUFX2_676 ( );
FILL FILL_0_INVX1_113 ( );
FILL FILL_0_BUFX2_319 ( );
FILL FILL_0_BUFX2_709 ( );
FILL FILL_0_OAI21X1_1645 ( );
FILL FILL_1_OAI21X1_1645 ( );
FILL FILL_0_DFFPOSX1_35 ( );
FILL FILL_1_DFFPOSX1_35 ( );
FILL FILL_2_DFFPOSX1_35 ( );
FILL FILL_3_DFFPOSX1_35 ( );
FILL FILL_4_DFFPOSX1_35 ( );
FILL FILL_5_DFFPOSX1_35 ( );
FILL FILL_6_DFFPOSX1_35 ( );
FILL FILL_0_BUFX2_864 ( );
FILL FILL_1_BUFX2_864 ( );
FILL FILL_0_BUFX2_677 ( );
FILL FILL_0_OAI21X1_1658 ( );
FILL FILL_1_OAI21X1_1658 ( );
FILL FILL_0_OAI21X1_1659 ( );
FILL FILL_1_OAI21X1_1659 ( );
FILL FILL_0_DFFPOSX1_42 ( );
FILL FILL_1_DFFPOSX1_42 ( );
FILL FILL_2_DFFPOSX1_42 ( );
FILL FILL_3_DFFPOSX1_42 ( );
FILL FILL_4_DFFPOSX1_42 ( );
FILL FILL_5_DFFPOSX1_42 ( );
FILL FILL_6_DFFPOSX1_42 ( );
FILL FILL_0_OAI21X1_1008 ( );
FILL FILL_1_OAI21X1_1008 ( );
FILL FILL_0_BUFX2_630 ( );
FILL FILL_1_BUFX2_630 ( );
FILL FILL_0_BUFX4_173 ( );
FILL FILL_1_BUFX4_173 ( );
FILL FILL_0_NAND2X1_11 ( );
FILL FILL_0_OAI21X1_11 ( );
FILL FILL_1_OAI21X1_11 ( );
FILL FILL_0_DFFPOSX1_167 ( );
FILL FILL_1_DFFPOSX1_167 ( );
FILL FILL_2_DFFPOSX1_167 ( );
FILL FILL_3_DFFPOSX1_167 ( );
FILL FILL_4_DFFPOSX1_167 ( );
FILL FILL_5_DFFPOSX1_167 ( );
FILL FILL_6_DFFPOSX1_167 ( );
FILL FILL_0_BUFX2_502 ( );
FILL FILL_1_BUFX2_502 ( );
FILL FILL_0_BUFX2_566 ( );
FILL FILL_0_OAI21X1_1709 ( );
FILL FILL_1_OAI21X1_1709 ( );
FILL FILL_0_OAI21X1_1708 ( );
FILL FILL_1_OAI21X1_1708 ( );
FILL FILL_0_DFFPOSX1_67 ( );
FILL FILL_1_DFFPOSX1_67 ( );
FILL FILL_2_DFFPOSX1_67 ( );
FILL FILL_3_DFFPOSX1_67 ( );
FILL FILL_4_DFFPOSX1_67 ( );
FILL FILL_5_DFFPOSX1_67 ( );
FILL FILL_0_CLKBUF1_66 ( );
FILL FILL_1_CLKBUF1_66 ( );
FILL FILL_2_CLKBUF1_66 ( );
FILL FILL_3_CLKBUF1_66 ( );
FILL FILL_4_CLKBUF1_66 ( );
FILL FILL_0_OAI21X1_403 ( );
FILL FILL_1_OAI21X1_403 ( );
FILL FILL_2_OAI21X1_403 ( );
FILL FILL_0_OAI21X1_402 ( );
FILL FILL_1_OAI21X1_402 ( );
FILL FILL_0_OAI21X1_672 ( );
FILL FILL_1_OAI21X1_672 ( );
FILL FILL_0_OAI21X1_673 ( );
FILL FILL_1_OAI21X1_673 ( );
FILL FILL_0_OAI21X1_405 ( );
FILL FILL_1_OAI21X1_405 ( );
FILL FILL_0_INVX2_40 ( );
FILL FILL_0_NOR2X1_102 ( );
FILL FILL_0_OAI21X1_676 ( );
FILL FILL_1_OAI21X1_676 ( );
FILL FILL_0_AND2X2_11 ( );
FILL FILL_1_AND2X2_11 ( );
FILL FILL_0_OAI21X1_517 ( );
FILL FILL_1_OAI21X1_517 ( );
FILL FILL_0_XNOR2X1_24 ( );
FILL FILL_1_XNOR2X1_24 ( );
FILL FILL_2_XNOR2X1_24 ( );
FILL FILL_0_OAI21X1_522 ( );
FILL FILL_1_OAI21X1_522 ( );
FILL FILL_0_DFFPOSX1_490 ( );
FILL FILL_1_DFFPOSX1_490 ( );
FILL FILL_2_DFFPOSX1_490 ( );
FILL FILL_3_DFFPOSX1_490 ( );
FILL FILL_4_DFFPOSX1_490 ( );
FILL FILL_5_DFFPOSX1_490 ( );
FILL FILL_6_DFFPOSX1_490 ( );
FILL FILL_0_BUFX2_626 ( );
FILL FILL_1_BUFX2_626 ( );
FILL FILL_0_CLKBUF1_46 ( );
FILL FILL_1_CLKBUF1_46 ( );
FILL FILL_2_CLKBUF1_46 ( );
FILL FILL_3_CLKBUF1_46 ( );
FILL FILL_4_CLKBUF1_46 ( );
FILL FILL_0_OAI21X1_532 ( );
FILL FILL_1_OAI21X1_532 ( );
FILL FILL_0_OAI21X1_531 ( );
FILL FILL_1_OAI21X1_531 ( );
FILL FILL_0_INVX4_30 ( );
FILL FILL_0_OAI21X1_690 ( );
FILL FILL_1_OAI21X1_690 ( );
FILL FILL_0_NOR2X1_10 ( );
FILL FILL_0_NAND2X1_166 ( );
FILL FILL_1_NAND2X1_166 ( );
FILL FILL_0_OAI21X1_689 ( );
FILL FILL_1_OAI21X1_689 ( );
FILL FILL_0_NAND2X1_310 ( );
FILL FILL_0_OAI21X1_410 ( );
FILL FILL_1_OAI21X1_410 ( );
FILL FILL_0_NAND2X1_162 ( );
FILL FILL_0_NOR2X1_7 ( );
FILL FILL_1_NOR2X1_7 ( );
FILL FILL_0_NAND3X1_1 ( );
FILL FILL_1_NAND3X1_1 ( );
FILL FILL_2_NAND3X1_1 ( );
FILL FILL_0_NOR2X1_40 ( );
FILL FILL_1_NOR2X1_40 ( );
FILL FILL_0_DFFPOSX1_500 ( );
FILL FILL_1_DFFPOSX1_500 ( );
FILL FILL_2_DFFPOSX1_500 ( );
FILL FILL_3_DFFPOSX1_500 ( );
FILL FILL_4_DFFPOSX1_500 ( );
FILL FILL_5_DFFPOSX1_500 ( );
FILL FILL_0_OAI21X1_466 ( );
FILL FILL_1_OAI21X1_466 ( );
FILL FILL_0_NAND2X1_248 ( );
FILL FILL_0_OAI21X1_471 ( );
FILL FILL_1_OAI21X1_471 ( );
FILL FILL_0_NAND2X1_318 ( );
FILL FILL_1_NAND2X1_318 ( );
FILL FILL_0_NAND2X1_181 ( );
FILL FILL_1_NAND2X1_181 ( );
FILL FILL_0_OAI21X1_661 ( );
FILL FILL_1_OAI21X1_661 ( );
FILL FILL_0_OAI21X1_660 ( );
FILL FILL_1_OAI21X1_660 ( );
FILL FILL_0_OAI21X1_585 ( );
FILL FILL_1_OAI21X1_585 ( );
FILL FILL_0_OAI21X1_586 ( );
FILL FILL_1_OAI21X1_586 ( );
FILL FILL_0_OAI21X1_589 ( );
FILL FILL_1_OAI21X1_589 ( );
FILL FILL_0_NAND2X1_247 ( );
FILL FILL_0_BUFX2_507 ( );
FILL FILL_1_BUFX2_507 ( );
FILL FILL_0_BUFX2_419 ( );
FILL FILL_1_BUFX2_419 ( );
FILL FILL_0_OAI21X1_590 ( );
FILL FILL_1_OAI21X1_590 ( );
FILL FILL_0_NAND2X1_105 ( );
FILL FILL_1_NAND2X1_105 ( );
FILL FILL_0_OAI21X1_587 ( );
FILL FILL_1_OAI21X1_587 ( );
FILL FILL_0_OAI21X1_588 ( );
FILL FILL_1_OAI21X1_588 ( );
FILL FILL_0_XNOR2X1_34 ( );
FILL FILL_1_XNOR2X1_34 ( );
FILL FILL_2_XNOR2X1_34 ( );
FILL FILL_3_XNOR2X1_34 ( );
FILL FILL_0_OAI21X1_451 ( );
FILL FILL_1_OAI21X1_451 ( );
FILL FILL_0_OAI21X1_389 ( );
FILL FILL_1_OAI21X1_389 ( );
FILL FILL_0_NOR2X1_24 ( );
FILL FILL_1_NOR2X1_24 ( );
FILL FILL_0_NAND2X1_203 ( );
FILL FILL_1_NAND2X1_203 ( );
FILL FILL_0_OAI21X1_448 ( );
FILL FILL_1_OAI21X1_448 ( );
FILL FILL_0_DFFPOSX1_417 ( );
FILL FILL_1_DFFPOSX1_417 ( );
FILL FILL_2_DFFPOSX1_417 ( );
FILL FILL_3_DFFPOSX1_417 ( );
FILL FILL_4_DFFPOSX1_417 ( );
FILL FILL_5_DFFPOSX1_417 ( );
FILL FILL_0_NAND2X1_170 ( );
FILL FILL_0_XNOR2X1_6 ( );
FILL FILL_1_XNOR2X1_6 ( );
FILL FILL_2_XNOR2X1_6 ( );
FILL FILL_3_XNOR2X1_6 ( );
FILL FILL_0_NAND2X1_169 ( );
FILL FILL_1_NAND2X1_169 ( );
FILL FILL_0_NAND2X1_173 ( );
FILL FILL_0_DFFPOSX1_438 ( );
FILL FILL_1_DFFPOSX1_438 ( );
FILL FILL_2_DFFPOSX1_438 ( );
FILL FILL_3_DFFPOSX1_438 ( );
FILL FILL_4_DFFPOSX1_438 ( );
FILL FILL_5_DFFPOSX1_438 ( );
FILL FILL_6_DFFPOSX1_438 ( );
FILL FILL_0_NOR2X1_14 ( );
FILL FILL_1_NOR2X1_14 ( );
FILL FILL_0_AND2X2_3 ( );
FILL FILL_1_AND2X2_3 ( );
FILL FILL_0_OAI21X1_430 ( );
FILL FILL_1_OAI21X1_430 ( );
FILL FILL_0_NAND3X1_27 ( );
FILL FILL_1_NAND3X1_27 ( );
FILL FILL_2_NAND3X1_27 ( );
FILL FILL_0_NOR2X1_107 ( );
FILL FILL_0_NOR2X1_65 ( );
FILL FILL_0_NAND2X1_99 ( );
FILL FILL_1_NAND2X1_99 ( );
FILL FILL_0_OAI21X1_441 ( );
FILL FILL_1_OAI21X1_441 ( );
FILL FILL_0_INVX4_13 ( );
FILL FILL_1_INVX4_13 ( );
FILL FILL_0_OAI21X1_602 ( );
FILL FILL_1_OAI21X1_602 ( );
FILL FILL_0_DFFPOSX1_522 ( );
FILL FILL_1_DFFPOSX1_522 ( );
FILL FILL_2_DFFPOSX1_522 ( );
FILL FILL_3_DFFPOSX1_522 ( );
FILL FILL_4_DFFPOSX1_522 ( );
FILL FILL_5_DFFPOSX1_522 ( );
FILL FILL_0_OAI21X1_436 ( );
FILL FILL_1_OAI21X1_436 ( );
FILL FILL_0_OAI21X1_435 ( );
FILL FILL_1_OAI21X1_435 ( );
FILL FILL_2_OAI21X1_435 ( );
FILL FILL_0_OAI21X1_304 ( );
FILL FILL_1_OAI21X1_304 ( );
FILL FILL_0_OAI21X1_572 ( );
FILL FILL_1_OAI21X1_572 ( );
FILL FILL_0_OAI21X1_359 ( );
FILL FILL_1_OAI21X1_359 ( );
FILL FILL_2_OAI21X1_359 ( );
FILL FILL_0_BUFX4_314 ( );
FILL FILL_1_BUFX4_314 ( );
FILL FILL_0_DFFPOSX1_334 ( );
FILL FILL_1_DFFPOSX1_334 ( );
FILL FILL_2_DFFPOSX1_334 ( );
FILL FILL_3_DFFPOSX1_334 ( );
FILL FILL_4_DFFPOSX1_334 ( );
FILL FILL_5_DFFPOSX1_334 ( );
FILL FILL_6_DFFPOSX1_334 ( );
FILL FILL_0_NAND2X1_423 ( );
FILL FILL_0_DFFPOSX1_387 ( );
FILL FILL_1_DFFPOSX1_387 ( );
FILL FILL_2_DFFPOSX1_387 ( );
FILL FILL_3_DFFPOSX1_387 ( );
FILL FILL_4_DFFPOSX1_387 ( );
FILL FILL_5_DFFPOSX1_387 ( );
FILL FILL_0_CLKBUF1_15 ( );
FILL FILL_1_CLKBUF1_15 ( );
FILL FILL_2_CLKBUF1_15 ( );
FILL FILL_3_CLKBUF1_15 ( );
FILL FILL_4_CLKBUF1_15 ( );
FILL FILL_0_BUFX2_1004 ( );
FILL FILL_1_BUFX2_1004 ( );
FILL FILL_0_NAND2X1_422 ( );
FILL FILL_1_NAND2X1_422 ( );
FILL FILL_0_OAI21X1_1060 ( );
FILL FILL_1_OAI21X1_1060 ( );
FILL FILL_0_BUFX4_354 ( );
FILL FILL_1_BUFX4_354 ( );
FILL FILL_0_BUFX2_835 ( );
FILL FILL_1_BUFX2_835 ( );
FILL FILL_0_OAI21X1_1140 ( );
FILL FILL_1_OAI21X1_1140 ( );
FILL FILL_2_OAI21X1_1140 ( );
FILL FILL_0_OAI21X1_1139 ( );
FILL FILL_1_OAI21X1_1139 ( );
FILL FILL_0_NAND2X1_506 ( );
FILL FILL_0_OAI21X1_1137 ( );
FILL FILL_1_OAI21X1_1137 ( );
FILL FILL_0_NOR2X1_138 ( );
FILL FILL_1_NOR2X1_138 ( );
FILL FILL_0_XNOR2X1_61 ( );
FILL FILL_1_XNOR2X1_61 ( );
FILL FILL_2_XNOR2X1_61 ( );
FILL FILL_3_XNOR2X1_61 ( );
FILL FILL_0_INVX1_187 ( );
FILL FILL_0_BUFX4_124 ( );
FILL FILL_1_BUFX4_124 ( );
FILL FILL_2_BUFX4_124 ( );
FILL FILL_0_OAI21X1_1133 ( );
FILL FILL_1_OAI21X1_1133 ( );
FILL FILL_0_DFFPOSX1_975 ( );
FILL FILL_1_DFFPOSX1_975 ( );
FILL FILL_2_DFFPOSX1_975 ( );
FILL FILL_3_DFFPOSX1_975 ( );
FILL FILL_4_DFFPOSX1_975 ( );
FILL FILL_5_DFFPOSX1_975 ( );
FILL FILL_6_DFFPOSX1_975 ( );
FILL FILL_0_NAND2X1_439 ( );
FILL FILL_1_NAND2X1_439 ( );
FILL FILL_0_OAI21X1_203 ( );
FILL FILL_1_OAI21X1_203 ( );
FILL FILL_0_OAI21X1_202 ( );
FILL FILL_1_OAI21X1_202 ( );
FILL FILL_0_DFFPOSX1_351 ( );
FILL FILL_1_DFFPOSX1_351 ( );
FILL FILL_2_DFFPOSX1_351 ( );
FILL FILL_3_DFFPOSX1_351 ( );
FILL FILL_4_DFFPOSX1_351 ( );
FILL FILL_5_DFFPOSX1_351 ( );
FILL FILL_6_DFFPOSX1_351 ( );
FILL FILL_0_OAI21X1_1309 ( );
FILL FILL_1_OAI21X1_1309 ( );
FILL FILL_0_CLKBUF1_53 ( );
FILL FILL_1_CLKBUF1_53 ( );
FILL FILL_2_CLKBUF1_53 ( );
FILL FILL_3_CLKBUF1_53 ( );
FILL FILL_4_CLKBUF1_53 ( );
FILL FILL_0_BUFX2_161 ( );
FILL FILL_1_BUFX2_161 ( );
FILL FILL_0_OAI21X1_1163 ( );
FILL FILL_1_OAI21X1_1163 ( );
FILL FILL_2_OAI21X1_1163 ( );
FILL FILL_0_INVX1_193 ( );
FILL FILL_0_OAI21X1_1162 ( );
FILL FILL_1_OAI21X1_1162 ( );
FILL FILL_0_NAND2X1_542 ( );
FILL FILL_1_NAND2X1_542 ( );
FILL FILL_0_OAI21X1_1498 ( );
FILL FILL_1_OAI21X1_1498 ( );
FILL FILL_0_DFFPOSX1_780 ( );
FILL FILL_1_DFFPOSX1_780 ( );
FILL FILL_2_DFFPOSX1_780 ( );
FILL FILL_3_DFFPOSX1_780 ( );
FILL FILL_4_DFFPOSX1_780 ( );
FILL FILL_5_DFFPOSX1_780 ( );
FILL FILL_6_DFFPOSX1_780 ( );
FILL FILL_0_BUFX2_160 ( );
FILL FILL_0_INVX4_42 ( );
FILL FILL_0_BUFX4_350 ( );
FILL FILL_1_BUFX4_350 ( );
FILL FILL_2_BUFX4_350 ( );
FILL FILL_0_OAI21X1_1304 ( );
FILL FILL_1_OAI21X1_1304 ( );
FILL FILL_0_OAI21X1_1305 ( );
FILL FILL_1_OAI21X1_1305 ( );
FILL FILL_2_OAI21X1_1305 ( );
FILL FILL_0_BUFX2_31 ( );
FILL FILL_1_BUFX2_31 ( );
FILL FILL_0_NAND2X1_454 ( );
FILL FILL_0_DFFPOSX1_794 ( );
FILL FILL_1_DFFPOSX1_794 ( );
FILL FILL_2_DFFPOSX1_794 ( );
FILL FILL_3_DFFPOSX1_794 ( );
FILL FILL_4_DFFPOSX1_794 ( );
FILL FILL_5_DFFPOSX1_794 ( );
FILL FILL_0_NAND2X1_452 ( );
FILL FILL_1_NAND2X1_452 ( );
FILL FILL_0_OAI21X1_1086 ( );
FILL FILL_1_OAI21X1_1086 ( );
FILL FILL_0_DFFPOSX1_859 ( );
FILL FILL_1_DFFPOSX1_859 ( );
FILL FILL_2_DFFPOSX1_859 ( );
FILL FILL_3_DFFPOSX1_859 ( );
FILL FILL_4_DFFPOSX1_859 ( );
FILL FILL_5_DFFPOSX1_859 ( );
FILL FILL_0_OAI21X1_1183 ( );
FILL FILL_1_OAI21X1_1183 ( );
FILL FILL_0_NAND2X1_569 ( );
FILL FILL_1_NAND2X1_569 ( );
FILL FILL_0_DFFPOSX1_926 ( );
FILL FILL_1_DFFPOSX1_926 ( );
FILL FILL_2_DFFPOSX1_926 ( );
FILL FILL_3_DFFPOSX1_926 ( );
FILL FILL_4_DFFPOSX1_926 ( );
FILL FILL_5_DFFPOSX1_926 ( );
FILL FILL_6_DFFPOSX1_926 ( );
FILL FILL_0_NOR2X1_171 ( );
FILL FILL_0_NAND2X1_579 ( );
FILL FILL_0_DFFPOSX1_865 ( );
FILL FILL_1_DFFPOSX1_865 ( );
FILL FILL_2_DFFPOSX1_865 ( );
FILL FILL_3_DFFPOSX1_865 ( );
FILL FILL_4_DFFPOSX1_865 ( );
FILL FILL_5_DFFPOSX1_865 ( );
FILL FILL_6_DFFPOSX1_865 ( );
FILL FILL_0_OAI21X1_1363 ( );
FILL FILL_1_OAI21X1_1363 ( );
FILL FILL_0_OAI21X1_1362 ( );
FILL FILL_1_OAI21X1_1362 ( );
FILL FILL_2_OAI21X1_1362 ( );
FILL FILL_0_AOI21X1_64 ( );
FILL FILL_1_AOI21X1_64 ( );
FILL FILL_2_AOI21X1_64 ( );
FILL FILL_0_INVX1_226 ( );
FILL FILL_0_AOI21X1_42 ( );
FILL FILL_1_AOI21X1_42 ( );
FILL FILL_0_NOR2X1_230 ( );
FILL FILL_1_NOR2X1_230 ( );
FILL FILL_0_OAI21X1_1364 ( );
FILL FILL_1_OAI21X1_1364 ( );
FILL FILL_0_OAI21X1_1552 ( );
FILL FILL_1_OAI21X1_1552 ( );
FILL FILL_0_DFFPOSX1_991 ( );
FILL FILL_1_DFFPOSX1_991 ( );
FILL FILL_2_DFFPOSX1_991 ( );
FILL FILL_3_DFFPOSX1_991 ( );
FILL FILL_4_DFFPOSX1_991 ( );
FILL FILL_5_DFFPOSX1_991 ( );
FILL FILL_6_DFFPOSX1_991 ( );
FILL FILL_0_BUFX2_245 ( );
FILL FILL_1_BUFX2_245 ( );
FILL FILL_0_BUFX2_117 ( );
FILL FILL_1_BUFX2_117 ( );
FILL FILL_0_CLKBUF1_38 ( );
FILL FILL_1_CLKBUF1_38 ( );
FILL FILL_2_CLKBUF1_38 ( );
FILL FILL_3_CLKBUF1_38 ( );
FILL FILL_4_CLKBUF1_38 ( );
FILL FILL_0_BUFX2_837 ( );
FILL FILL_1_BUFX2_837 ( );
FILL FILL_0_OAI21X1_920 ( );
FILL FILL_1_OAI21X1_920 ( );
FILL FILL_0_BUFX2_50 ( );
FILL FILL_1_BUFX2_50 ( );
FILL FILL_0_OAI21X1_916 ( );
FILL FILL_1_OAI21X1_916 ( );
FILL FILL_0_OAI21X1_1004 ( );
FILL FILL_1_OAI21X1_1004 ( );
FILL FILL_0_BUFX2_758 ( );
FILL FILL_0_OAI21X1_1005 ( );
FILL FILL_1_OAI21X1_1005 ( );
FILL FILL_0_OAI21X1_1034 ( );
FILL FILL_1_OAI21X1_1034 ( );
FILL FILL_0_OAI21X1_1035 ( );
FILL FILL_1_OAI21X1_1035 ( );
FILL FILL_0_BUFX2_743 ( );
FILL FILL_1_BUFX2_743 ( );
FILL FILL_0_NAND2X1_351 ( );
FILL FILL_1_NAND2X1_351 ( );
FILL FILL_0_BUFX2_1028 ( );
FILL FILL_0_INVX1_81 ( );
FILL FILL_0_NAND2X1_713 ( );
FILL FILL_0_INVX2_6 ( );
FILL FILL_0_BUFX2_900 ( );
FILL FILL_1_BUFX2_900 ( );
FILL FILL_0_NAND2X1_688 ( );
FILL FILL_0_OAI21X1_1620 ( );
FILL FILL_1_OAI21X1_1620 ( );
FILL FILL_0_DFFPOSX1_10 ( );
FILL FILL_1_DFFPOSX1_10 ( );
FILL FILL_2_DFFPOSX1_10 ( );
FILL FILL_3_DFFPOSX1_10 ( );
FILL FILL_4_DFFPOSX1_10 ( );
FILL FILL_5_DFFPOSX1_10 ( );
FILL FILL_0_NAND2X1_656 ( );
FILL FILL_1_NAND2X1_656 ( );
FILL FILL_0_OAI21X1_1587 ( );
FILL FILL_1_OAI21X1_1587 ( );
FILL FILL_0_DFFPOSX1_1010 ( );
FILL FILL_1_DFFPOSX1_1010 ( );
FILL FILL_2_DFFPOSX1_1010 ( );
FILL FILL_3_DFFPOSX1_1010 ( );
FILL FILL_4_DFFPOSX1_1010 ( );
FILL FILL_5_DFFPOSX1_1010 ( );
FILL FILL_6_DFFPOSX1_1010 ( );
FILL FILL_0_BUFX4_217 ( );
FILL FILL_1_BUFX4_217 ( );
FILL FILL_0_OAI21X1_674 ( );
FILL FILL_1_OAI21X1_674 ( );
FILL FILL_0_DFFPOSX1_553 ( );
FILL FILL_1_DFFPOSX1_553 ( );
FILL FILL_2_DFFPOSX1_553 ( );
FILL FILL_3_DFFPOSX1_553 ( );
FILL FILL_4_DFFPOSX1_553 ( );
FILL FILL_5_DFFPOSX1_553 ( );
FILL FILL_6_DFFPOSX1_553 ( );
FILL FILL_0_OAI21X1_675 ( );
FILL FILL_1_OAI21X1_675 ( );
FILL FILL_2_OAI21X1_675 ( );
FILL FILL_0_NAND2X1_146 ( );
FILL FILL_0_OAI21X1_404 ( );
FILL FILL_1_OAI21X1_404 ( );
FILL FILL_0_DFFPOSX1_425 ( );
FILL FILL_1_DFFPOSX1_425 ( );
FILL FILL_2_DFFPOSX1_425 ( );
FILL FILL_3_DFFPOSX1_425 ( );
FILL FILL_4_DFFPOSX1_425 ( );
FILL FILL_5_DFFPOSX1_425 ( );
FILL FILL_6_DFFPOSX1_425 ( );
FILL FILL_0_INVX2_11 ( );
FILL FILL_0_OAI21X1_677 ( );
FILL FILL_1_OAI21X1_677 ( );
FILL FILL_0_DFFPOSX1_554 ( );
FILL FILL_1_DFFPOSX1_554 ( );
FILL FILL_2_DFFPOSX1_554 ( );
FILL FILL_3_DFFPOSX1_554 ( );
FILL FILL_4_DFFPOSX1_554 ( );
FILL FILL_5_DFFPOSX1_554 ( );
FILL FILL_0_NAND2X1_145 ( );
FILL FILL_0_OAI21X1_678 ( );
FILL FILL_1_OAI21X1_678 ( );
FILL FILL_0_NOR2X1_103 ( );
FILL FILL_1_NOR2X1_103 ( );
FILL FILL_0_INVX2_52 ( );
FILL FILL_0_OAI21X1_679 ( );
FILL FILL_1_OAI21X1_679 ( );
FILL FILL_0_INVX1_34 ( );
FILL FILL_0_OAI21X1_521 ( );
FILL FILL_1_OAI21X1_521 ( );
FILL FILL_0_OAI21X1_518 ( );
FILL FILL_1_OAI21X1_518 ( );
FILL FILL_0_OAI21X1_519 ( );
FILL FILL_1_OAI21X1_519 ( );
FILL FILL_0_NOR2X1_4 ( );
FILL FILL_0_AND2X2_1 ( );
FILL FILL_1_AND2X2_1 ( );
FILL FILL_0_AND2X2_18 ( );
FILL FILL_1_AND2X2_18 ( );
FILL FILL_0_DFFPOSX1_561 ( );
FILL FILL_1_DFFPOSX1_561 ( );
FILL FILL_2_DFFPOSX1_561 ( );
FILL FILL_3_DFFPOSX1_561 ( );
FILL FILL_4_DFFPOSX1_561 ( );
FILL FILL_5_DFFPOSX1_561 ( );
FILL FILL_0_AND2X2_19 ( );
FILL FILL_1_AND2X2_19 ( );
FILL FILL_0_NOR2X1_104 ( );
FILL FILL_1_NOR2X1_104 ( );
FILL FILL_0_OAI21X1_698 ( );
FILL FILL_1_OAI21X1_698 ( );
FILL FILL_2_OAI21X1_698 ( );
FILL FILL_0_AND2X2_20 ( );
FILL FILL_1_AND2X2_20 ( );
FILL FILL_0_NAND2X1_272 ( );
FILL FILL_1_NAND2X1_272 ( );
FILL FILL_0_INVX1_9 ( );
FILL FILL_0_AND2X2_12 ( );
FILL FILL_1_AND2X2_12 ( );
FILL FILL_0_NAND3X1_14 ( );
FILL FILL_1_NAND3X1_14 ( );
FILL FILL_0_NAND2X1_165 ( );
FILL FILL_1_NAND2X1_165 ( );
FILL FILL_0_NAND2X1_167 ( );
FILL FILL_1_NAND2X1_167 ( );
FILL FILL_0_AND2X2_2 ( );
FILL FILL_1_AND2X2_2 ( );
FILL FILL_0_NAND3X1_15 ( );
FILL FILL_1_NAND3X1_15 ( );
FILL FILL_2_NAND3X1_15 ( );
FILL FILL_0_NOR2X1_62 ( );
FILL FILL_0_DFFPOSX1_496 ( );
FILL FILL_1_DFFPOSX1_496 ( );
FILL FILL_2_DFFPOSX1_496 ( );
FILL FILL_3_DFFPOSX1_496 ( );
FILL FILL_4_DFFPOSX1_496 ( );
FILL FILL_5_DFFPOSX1_496 ( );
FILL FILL_0_DFFPOSX1_369 ( );
FILL FILL_1_DFFPOSX1_369 ( );
FILL FILL_2_DFFPOSX1_369 ( );
FILL FILL_3_DFFPOSX1_369 ( );
FILL FILL_4_DFFPOSX1_369 ( );
FILL FILL_5_DFFPOSX1_369 ( );
FILL FILL_6_DFFPOSX1_369 ( );
FILL FILL_0_BUFX2_564 ( );
FILL FILL_1_BUFX2_564 ( );
FILL FILL_0_DFFPOSX1_475 ( );
FILL FILL_1_DFFPOSX1_475 ( );
FILL FILL_2_DFFPOSX1_475 ( );
FILL FILL_3_DFFPOSX1_475 ( );
FILL FILL_4_DFFPOSX1_475 ( );
FILL FILL_5_DFFPOSX1_475 ( );
FILL FILL_6_DFFPOSX1_475 ( );
FILL FILL_0_OAI21X1_480 ( );
FILL FILL_1_OAI21X1_480 ( );
FILL FILL_0_OAI21X1_470 ( );
FILL FILL_1_OAI21X1_470 ( );
FILL FILL_2_OAI21X1_470 ( );
FILL FILL_0_BUFX4_335 ( );
FILL FILL_1_BUFX4_335 ( );
FILL FILL_0_OAI21X1_705 ( );
FILL FILL_1_OAI21X1_705 ( );
FILL FILL_0_BUFX2_571 ( );
FILL FILL_0_DFFPOSX1_474 ( );
FILL FILL_1_DFFPOSX1_474 ( );
FILL FILL_2_DFFPOSX1_474 ( );
FILL FILL_3_DFFPOSX1_474 ( );
FILL FILL_4_DFFPOSX1_474 ( );
FILL FILL_5_DFFPOSX1_474 ( );
FILL FILL_0_DFFPOSX1_389 ( );
FILL FILL_1_DFFPOSX1_389 ( );
FILL FILL_2_DFFPOSX1_389 ( );
FILL FILL_3_DFFPOSX1_389 ( );
FILL FILL_4_DFFPOSX1_389 ( );
FILL FILL_5_DFFPOSX1_389 ( );
FILL FILL_0_OAI21X1_361 ( );
FILL FILL_1_OAI21X1_361 ( );
FILL FILL_0_INVX4_15 ( );
FILL FILL_1_INVX4_15 ( );
FILL FILL_0_NAND2X1_206 ( );
FILL FILL_1_NAND2X1_206 ( );
FILL FILL_0_OAI21X1_833 ( );
FILL FILL_1_OAI21X1_833 ( );
FILL FILL_0_NOR2X1_26 ( );
FILL FILL_1_NOR2X1_26 ( );
FILL FILL_0_INVX1_16 ( );
FILL FILL_0_DFFPOSX1_581 ( );
FILL FILL_1_DFFPOSX1_581 ( );
FILL FILL_2_DFFPOSX1_581 ( );
FILL FILL_3_DFFPOSX1_581 ( );
FILL FILL_4_DFFPOSX1_581 ( );
FILL FILL_5_DFFPOSX1_581 ( );
FILL FILL_6_DFFPOSX1_581 ( );
FILL FILL_0_NOR2X1_23 ( );
FILL FILL_0_BUFX2_424 ( );
FILL FILL_1_BUFX2_424 ( );
FILL FILL_0_DFFPOSX1_437 ( );
FILL FILL_1_DFFPOSX1_437 ( );
FILL FILL_2_DFFPOSX1_437 ( );
FILL FILL_3_DFFPOSX1_437 ( );
FILL FILL_4_DFFPOSX1_437 ( );
FILL FILL_5_DFFPOSX1_437 ( );
FILL FILL_0_OAI21X1_425 ( );
FILL FILL_1_OAI21X1_425 ( );
FILL FILL_2_OAI21X1_425 ( );
FILL FILL_0_DFFPOSX1_436 ( );
FILL FILL_1_DFFPOSX1_436 ( );
FILL FILL_2_DFFPOSX1_436 ( );
FILL FILL_3_DFFPOSX1_436 ( );
FILL FILL_4_DFFPOSX1_436 ( );
FILL FILL_5_DFFPOSX1_436 ( );
FILL FILL_6_DFFPOSX1_436 ( );
FILL FILL_0_XNOR2X1_7 ( );
FILL FILL_1_XNOR2X1_7 ( );
FILL FILL_2_XNOR2X1_7 ( );
FILL FILL_3_XNOR2X1_7 ( );
FILL FILL_0_NAND2X1_277 ( );
FILL FILL_1_NAND2X1_277 ( );
FILL FILL_0_NOR2X1_13 ( );
FILL FILL_0_NAND2X1_177 ( );
FILL FILL_1_NAND2X1_177 ( );
FILL FILL_0_NOR2X1_15 ( );
FILL FILL_1_NOR2X1_15 ( );
FILL FILL_0_DFFPOSX1_383 ( );
FILL FILL_1_DFFPOSX1_383 ( );
FILL FILL_2_DFFPOSX1_383 ( );
FILL FILL_3_DFFPOSX1_383 ( );
FILL FILL_4_DFFPOSX1_383 ( );
FILL FILL_5_DFFPOSX1_383 ( );
FILL FILL_0_OAI21X1_440 ( );
FILL FILL_1_OAI21X1_440 ( );
FILL FILL_0_OAI21X1_442 ( );
FILL FILL_1_OAI21X1_442 ( );
FILL FILL_0_NAND2X1_196 ( );
FILL FILL_1_NAND2X1_196 ( );
FILL FILL_0_XNOR2X1_11 ( );
FILL FILL_1_XNOR2X1_11 ( );
FILL FILL_2_XNOR2X1_11 ( );
FILL FILL_3_XNOR2X1_11 ( );
FILL FILL_0_NOR2X1_71 ( );
FILL FILL_0_NAND2X1_190 ( );
FILL FILL_0_OAI21X1_574 ( );
FILL FILL_1_OAI21X1_574 ( );
FILL FILL_0_DFFPOSX1_511 ( );
FILL FILL_1_DFFPOSX1_511 ( );
FILL FILL_2_DFFPOSX1_511 ( );
FILL FILL_3_DFFPOSX1_511 ( );
FILL FILL_4_DFFPOSX1_511 ( );
FILL FILL_5_DFFPOSX1_511 ( );
FILL FILL_0_BUFX2_607 ( );
FILL FILL_0_NAND2X1_101 ( );
FILL FILL_1_NAND2X1_101 ( );
FILL FILL_0_OAI21X1_284 ( );
FILL FILL_1_OAI21X1_284 ( );
FILL FILL_0_OAI21X1_285 ( );
FILL FILL_1_OAI21X1_285 ( );
FILL FILL_2_OAI21X1_285 ( );
FILL FILL_0_DFFPOSX1_765 ( );
FILL FILL_1_DFFPOSX1_765 ( );
FILL FILL_2_DFFPOSX1_765 ( );
FILL FILL_3_DFFPOSX1_765 ( );
FILL FILL_4_DFFPOSX1_765 ( );
FILL FILL_5_DFFPOSX1_765 ( );
FILL FILL_6_DFFPOSX1_765 ( );
FILL FILL_0_OAI21X1_1057 ( );
FILL FILL_1_OAI21X1_1057 ( );
FILL FILL_0_DFFPOSX1_764 ( );
FILL FILL_1_DFFPOSX1_764 ( );
FILL FILL_2_DFFPOSX1_764 ( );
FILL FILL_3_DFFPOSX1_764 ( );
FILL FILL_4_DFFPOSX1_764 ( );
FILL FILL_5_DFFPOSX1_764 ( );
FILL FILL_0_OAI21X1_1056 ( );
FILL FILL_1_OAI21X1_1056 ( );
FILL FILL_0_XNOR2X1_60 ( );
FILL FILL_1_XNOR2X1_60 ( );
FILL FILL_2_XNOR2X1_60 ( );
FILL FILL_3_XNOR2X1_60 ( );
FILL FILL_0_NAND2X1_507 ( );
FILL FILL_1_NAND2X1_507 ( );
FILL FILL_0_OAI21X1_1135 ( );
FILL FILL_1_OAI21X1_1135 ( );
FILL FILL_2_OAI21X1_1135 ( );
FILL FILL_0_INVX4_35 ( );
FILL FILL_0_OAI21X1_1136 ( );
FILL FILL_1_OAI21X1_1136 ( );
FILL FILL_0_DFFPOSX1_828 ( );
FILL FILL_1_DFFPOSX1_828 ( );
FILL FILL_2_DFFPOSX1_828 ( );
FILL FILL_3_DFFPOSX1_828 ( );
FILL FILL_4_DFFPOSX1_828 ( );
FILL FILL_5_DFFPOSX1_828 ( );
FILL FILL_6_DFFPOSX1_828 ( );
FILL FILL_0_NOR2X1_139 ( );
FILL FILL_1_NOR2X1_139 ( );
FILL FILL_0_DFFPOSX1_293 ( );
FILL FILL_1_DFFPOSX1_293 ( );
FILL FILL_2_DFFPOSX1_293 ( );
FILL FILL_3_DFFPOSX1_293 ( );
FILL FILL_4_DFFPOSX1_293 ( );
FILL FILL_5_DFFPOSX1_293 ( );
FILL FILL_6_DFFPOSX1_293 ( );
FILL FILL_0_INVX2_113 ( );
FILL FILL_0_BUFX2_208 ( );
FILL FILL_1_BUFX2_208 ( );
FILL FILL_0_DFFPOSX1_781 ( );
FILL FILL_1_DFFPOSX1_781 ( );
FILL FILL_2_DFFPOSX1_781 ( );
FILL FILL_3_DFFPOSX1_781 ( );
FILL FILL_4_DFFPOSX1_781 ( );
FILL FILL_5_DFFPOSX1_781 ( );
FILL FILL_0_CLKBUF1_28 ( );
FILL FILL_1_CLKBUF1_28 ( );
FILL FILL_2_CLKBUF1_28 ( );
FILL FILL_3_CLKBUF1_28 ( );
FILL FILL_4_CLKBUF1_28 ( );
FILL FILL_0_BUFX2_142 ( );
FILL FILL_0_DFFPOSX1_846 ( );
FILL FILL_1_DFFPOSX1_846 ( );
FILL FILL_2_DFFPOSX1_846 ( );
FILL FILL_3_DFFPOSX1_846 ( );
FILL FILL_4_DFFPOSX1_846 ( );
FILL FILL_5_DFFPOSX1_846 ( );
FILL FILL_0_OAI21X1_1072 ( );
FILL FILL_1_OAI21X1_1072 ( );
FILL FILL_0_INVX2_77 ( );
FILL FILL_1_INVX2_77 ( );
FILL FILL_0_NAND2X1_438 ( );
FILL FILL_0_INVX2_76 ( );
FILL FILL_0_NAND2X1_638 ( );
FILL FILL_1_NAND2X1_638 ( );
FILL FILL_0_OAI21X1_1499 ( );
FILL FILL_1_OAI21X1_1499 ( );
FILL FILL_0_DFFPOSX1_974 ( );
FILL FILL_1_DFFPOSX1_974 ( );
FILL FILL_2_DFFPOSX1_974 ( );
FILL FILL_3_DFFPOSX1_974 ( );
FILL FILL_4_DFFPOSX1_974 ( );
FILL FILL_5_DFFPOSX1_974 ( );
FILL FILL_0_DFFPOSX1_913 ( );
FILL FILL_1_DFFPOSX1_913 ( );
FILL FILL_2_DFFPOSX1_913 ( );
FILL FILL_3_DFFPOSX1_913 ( );
FILL FILL_4_DFFPOSX1_913 ( );
FILL FILL_5_DFFPOSX1_913 ( );
FILL FILL_6_DFFPOSX1_913 ( );
FILL FILL_0_OAI21X1_1545 ( );
FILL FILL_1_OAI21X1_1545 ( );
FILL FILL_2_OAI21X1_1545 ( );
FILL FILL_0_DFFPOSX1_796 ( );
FILL FILL_1_DFFPOSX1_796 ( );
FILL FILL_2_DFFPOSX1_796 ( );
FILL FILL_3_DFFPOSX1_796 ( );
FILL FILL_4_DFFPOSX1_796 ( );
FILL FILL_5_DFFPOSX1_796 ( );
FILL FILL_6_DFFPOSX1_796 ( );
FILL FILL_0_BUFX2_223 ( );
FILL FILL_1_BUFX2_223 ( );
FILL FILL_0_XNOR2X1_103 ( );
FILL FILL_1_XNOR2X1_103 ( );
FILL FILL_2_XNOR2X1_103 ( );
FILL FILL_3_XNOR2X1_103 ( );
FILL FILL_0_DFFPOSX1_860 ( );
FILL FILL_1_DFFPOSX1_860 ( );
FILL FILL_2_DFFPOSX1_860 ( );
FILL FILL_3_DFFPOSX1_860 ( );
FILL FILL_4_DFFPOSX1_860 ( );
FILL FILL_5_DFFPOSX1_860 ( );
FILL FILL_0_NAND2X1_570 ( );
FILL FILL_1_NAND2X1_570 ( );
FILL FILL_0_DFFPOSX1_861 ( );
FILL FILL_1_DFFPOSX1_861 ( );
FILL FILL_2_DFFPOSX1_861 ( );
FILL FILL_3_DFFPOSX1_861 ( );
FILL FILL_4_DFFPOSX1_861 ( );
FILL FILL_5_DFFPOSX1_861 ( );
FILL FILL_6_DFFPOSX1_861 ( );
FILL FILL_0_NAND2X1_573 ( );
FILL FILL_1_NAND2X1_573 ( );
FILL FILL_0_BUFX2_114 ( );
FILL FILL_1_BUFX2_114 ( );
FILL FILL_0_NAND2X1_575 ( );
FILL FILL_1_NAND2X1_575 ( );
FILL FILL_0_OAI21X1_1192 ( );
FILL FILL_1_OAI21X1_1192 ( );
FILL FILL_2_OAI21X1_1192 ( );
FILL FILL_0_OAI21X1_1190 ( );
FILL FILL_1_OAI21X1_1190 ( );
FILL FILL_0_AOI21X1_43 ( );
FILL FILL_1_AOI21X1_43 ( );
FILL FILL_2_AOI21X1_43 ( );
FILL FILL_0_OAI21X1_1195 ( );
FILL FILL_1_OAI21X1_1195 ( );
FILL FILL_0_NAND2X1_644 ( );
FILL FILL_1_NAND2X1_644 ( );
FILL FILL_0_INVX4_45 ( );
FILL FILL_1_INVX4_45 ( );
FILL FILL_0_OAI21X1_1554 ( );
FILL FILL_1_OAI21X1_1554 ( );
FILL FILL_0_OAI21X1_1555 ( );
FILL FILL_1_OAI21X1_1555 ( );
FILL FILL_0_DFFPOSX1_992 ( );
FILL FILL_1_DFFPOSX1_992 ( );
FILL FILL_2_DFFPOSX1_992 ( );
FILL FILL_3_DFFPOSX1_992 ( );
FILL FILL_4_DFFPOSX1_992 ( );
FILL FILL_5_DFFPOSX1_992 ( );
FILL FILL_0_OAI21X1_1551 ( );
FILL FILL_1_OAI21X1_1551 ( );
FILL FILL_0_OAI21X1_1193 ( );
FILL FILL_1_OAI21X1_1193 ( );
FILL FILL_0_DFFPOSX1_864 ( );
FILL FILL_1_DFFPOSX1_864 ( );
FILL FILL_2_DFFPOSX1_864 ( );
FILL FILL_3_DFFPOSX1_864 ( );
FILL FILL_4_DFFPOSX1_864 ( );
FILL FILL_5_DFFPOSX1_864 ( );
FILL FILL_0_NAND2X1_578 ( );
FILL FILL_1_NAND2X1_578 ( );
FILL FILL_0_OAI21X1_7 ( );
FILL FILL_1_OAI21X1_7 ( );
FILL FILL_0_NAND2X1_7 ( );
FILL FILL_0_DFFPOSX1_163 ( );
FILL FILL_1_DFFPOSX1_163 ( );
FILL FILL_2_DFFPOSX1_163 ( );
FILL FILL_3_DFFPOSX1_163 ( );
FILL FILL_4_DFFPOSX1_163 ( );
FILL FILL_5_DFFPOSX1_163 ( );
FILL FILL_6_DFFPOSX1_163 ( );
FILL FILL_0_BUFX2_176 ( );
FILL FILL_0_OAI21X1_1610 ( );
FILL FILL_1_OAI21X1_1610 ( );
FILL FILL_2_OAI21X1_1610 ( );
FILL FILL_0_INVX1_115 ( );
FILL FILL_0_NAND2X1_679 ( );
FILL FILL_0_DFFPOSX1_1 ( );
FILL FILL_1_DFFPOSX1_1 ( );
FILL FILL_2_DFFPOSX1_1 ( );
FILL FILL_3_DFFPOSX1_1 ( );
FILL FILL_4_DFFPOSX1_1 ( );
FILL FILL_5_DFFPOSX1_1 ( );
FILL FILL_0_DFFPOSX1_728 ( );
FILL FILL_1_DFFPOSX1_728 ( );
FILL FILL_2_DFFPOSX1_728 ( );
FILL FILL_3_DFFPOSX1_728 ( );
FILL FILL_4_DFFPOSX1_728 ( );
FILL FILL_5_DFFPOSX1_728 ( );
FILL FILL_6_DFFPOSX1_728 ( );
FILL FILL_0_INVX2_114 ( );
FILL FILL_0_BUFX2_333 ( );
FILL FILL_1_BUFX2_333 ( );
FILL FILL_0_NAND2X1_374 ( );
FILL FILL_1_NAND2X1_374 ( );
FILL FILL_0_OAI21X1_880 ( );
FILL FILL_1_OAI21X1_880 ( );
FILL FILL_0_BUFX2_1031 ( );
FILL FILL_0_BUFX2_836 ( );
FILL FILL_0_BUFX2_882 ( );
FILL FILL_1_BUFX2_882 ( );
FILL FILL_0_DFFPOSX1_226 ( );
FILL FILL_1_DFFPOSX1_226 ( );
FILL FILL_2_DFFPOSX1_226 ( );
FILL FILL_3_DFFPOSX1_226 ( );
FILL FILL_4_DFFPOSX1_226 ( );
FILL FILL_5_DFFPOSX1_226 ( );
FILL FILL_6_DFFPOSX1_226 ( );
FILL FILL_0_OAI21X1_70 ( );
FILL FILL_1_OAI21X1_70 ( );
FILL FILL_0_NAND2X1_70 ( );
FILL FILL_1_NAND2X1_70 ( );
FILL FILL_0_BUFX2_818 ( );
FILL FILL_0_DFFPOSX1_146 ( );
FILL FILL_1_DFFPOSX1_146 ( );
FILL FILL_2_DFFPOSX1_146 ( );
FILL FILL_3_DFFPOSX1_146 ( );
FILL FILL_4_DFFPOSX1_146 ( );
FILL FILL_5_DFFPOSX1_146 ( );
FILL FILL_6_DFFPOSX1_146 ( );
FILL FILL_0_BUFX2_427 ( );
FILL FILL_1_BUFX2_427 ( );
FILL FILL_0_NAND2X1_76 ( );
FILL FILL_1_NAND2X1_76 ( );
FILL FILL_0_DFFPOSX1_360 ( );
FILL FILL_1_DFFPOSX1_360 ( );
FILL FILL_2_DFFPOSX1_360 ( );
FILL FILL_3_DFFPOSX1_360 ( );
FILL FILL_4_DFFPOSX1_360 ( );
FILL FILL_5_DFFPOSX1_360 ( );
FILL FILL_6_DFFPOSX1_360 ( );
FILL FILL_0_OAI21X1_332 ( );
FILL FILL_1_OAI21X1_332 ( );
FILL FILL_0_DFFPOSX1_487 ( );
FILL FILL_1_DFFPOSX1_487 ( );
FILL FILL_2_DFFPOSX1_487 ( );
FILL FILL_3_DFFPOSX1_487 ( );
FILL FILL_4_DFFPOSX1_487 ( );
FILL FILL_5_DFFPOSX1_487 ( );
FILL FILL_0_OAI21X1_507 ( );
FILL FILL_1_OAI21X1_507 ( );
FILL FILL_0_OAI21X1_508 ( );
FILL FILL_1_OAI21X1_508 ( );
FILL FILL_0_INVX1_25 ( );
FILL FILL_0_XNOR2X1_40 ( );
FILL FILL_1_XNOR2X1_40 ( );
FILL FILL_2_XNOR2X1_40 ( );
FILL FILL_3_XNOR2X1_40 ( );
FILL FILL_0_NAND2X1_268 ( );
FILL FILL_1_NAND2X1_268 ( );
FILL FILL_0_NAND2X1_269 ( );
FILL FILL_1_NAND2X1_269 ( );
FILL FILL_0_NOR2X1_58 ( );
FILL FILL_1_NOR2X1_58 ( );
FILL FILL_0_INVX4_29 ( );
FILL FILL_1_INVX4_29 ( );
FILL FILL_0_BUFX2_800 ( );
FILL FILL_0_BUFX2_524 ( );
FILL FILL_0_DFFPOSX1_491 ( );
FILL FILL_1_DFFPOSX1_491 ( );
FILL FILL_2_DFFPOSX1_491 ( );
FILL FILL_3_DFFPOSX1_491 ( );
FILL FILL_4_DFFPOSX1_491 ( );
FILL FILL_5_DFFPOSX1_491 ( );
FILL FILL_0_OAI21X1_520 ( );
FILL FILL_1_OAI21X1_520 ( );
FILL FILL_0_NAND2X1_309 ( );
FILL FILL_0_BUFX2_434 ( );
FILL FILL_1_BUFX2_434 ( );
FILL FILL_0_NAND2X1_150 ( );
FILL FILL_1_NAND2X1_150 ( );
FILL FILL_0_NAND2X1_308 ( );
FILL FILL_1_NAND2X1_308 ( );
FILL FILL_0_OAI21X1_696 ( );
FILL FILL_1_OAI21X1_696 ( );
FILL FILL_2_OAI21X1_696 ( );
FILL FILL_0_OAI21X1_697 ( );
FILL FILL_1_OAI21X1_697 ( );
FILL FILL_0_XNOR2X1_42 ( );
FILL FILL_1_XNOR2X1_42 ( );
FILL FILL_2_XNOR2X1_42 ( );
FILL FILL_0_NAND2X1_314 ( );
FILL FILL_1_NAND2X1_314 ( );
FILL FILL_0_INVX2_17 ( );
FILL FILL_0_OAI21X1_693 ( );
FILL FILL_1_OAI21X1_693 ( );
FILL FILL_0_NAND2X1_313 ( );
FILL FILL_0_XNOR2X1_27 ( );
FILL FILL_1_XNOR2X1_27 ( );
FILL FILL_2_XNOR2X1_27 ( );
FILL FILL_3_XNOR2X1_27 ( );
FILL FILL_0_OAI21X1_545 ( );
FILL FILL_1_OAI21X1_545 ( );
FILL FILL_0_OAI21X1_704 ( );
FILL FILL_1_OAI21X1_704 ( );
FILL FILL_0_OAI21X1_539 ( );
FILL FILL_1_OAI21X1_539 ( );
FILL FILL_0_INVX1_26 ( );
FILL FILL_0_NOR2X1_8 ( );
FILL FILL_0_INVX1_1 ( );
FILL FILL_0_NAND2X1_276 ( );
FILL FILL_0_OAI21X1_546 ( );
FILL FILL_1_OAI21X1_546 ( );
FILL FILL_2_OAI21X1_546 ( );
FILL FILL_0_OAI21X1_544 ( );
FILL FILL_1_OAI21X1_544 ( );
FILL FILL_0_OAI21X1_341 ( );
FILL FILL_1_OAI21X1_341 ( );
FILL FILL_2_OAI21X1_341 ( );
FILL FILL_0_NAND2X1_85 ( );
FILL FILL_0_DFFPOSX1_404 ( );
FILL FILL_1_DFFPOSX1_404 ( );
FILL FILL_2_DFFPOSX1_404 ( );
FILL FILL_3_DFFPOSX1_404 ( );
FILL FILL_4_DFFPOSX1_404 ( );
FILL FILL_5_DFFPOSX1_404 ( );
FILL FILL_0_NAND2X1_120 ( );
FILL FILL_0_BUFX2_573 ( );
FILL FILL_0_OAI21X1_484 ( );
FILL FILL_1_OAI21X1_484 ( );
FILL FILL_0_OAI21X1_485 ( );
FILL FILL_1_OAI21X1_485 ( );
FILL FILL_0_XNOR2X1_22 ( );
FILL FILL_1_XNOR2X1_22 ( );
FILL FILL_2_XNOR2X1_22 ( );
FILL FILL_3_XNOR2X1_22 ( );
FILL FILL_0_DFFPOSX1_564 ( );
FILL FILL_1_DFFPOSX1_564 ( );
FILL FILL_2_DFFPOSX1_564 ( );
FILL FILL_3_DFFPOSX1_564 ( );
FILL FILL_4_DFFPOSX1_564 ( );
FILL FILL_5_DFFPOSX1_564 ( );
FILL FILL_6_DFFPOSX1_564 ( );
FILL FILL_0_OAI21X1_706 ( );
FILL FILL_1_OAI21X1_706 ( );
FILL FILL_0_OAI21X1_483 ( );
FILL FILL_1_OAI21X1_483 ( );
FILL FILL_0_BUFX2_551 ( );
FILL FILL_1_BUFX2_551 ( );
FILL FILL_0_BUFX2_453 ( );
FILL FILL_1_BUFX2_453 ( );
FILL FILL_0_BUFX4_373 ( );
FILL FILL_1_BUFX4_373 ( );
FILL FILL_0_NAND2X1_135 ( );
FILL FILL_1_NAND2X1_135 ( );
FILL FILL_0_BUFX2_634 ( );
FILL FILL_1_BUFX2_634 ( );
FILL FILL_0_OAI21X1_751 ( );
FILL FILL_1_OAI21X1_751 ( );
FILL FILL_0_OAI21X1_752 ( );
FILL FILL_1_OAI21X1_752 ( );
FILL FILL_2_OAI21X1_752 ( );
FILL FILL_0_OAI21X1_834 ( );
FILL FILL_1_OAI21X1_834 ( );
FILL FILL_2_OAI21X1_834 ( );
FILL FILL_0_DFFPOSX1_608 ( );
FILL FILL_1_DFFPOSX1_608 ( );
FILL FILL_2_DFFPOSX1_608 ( );
FILL FILL_3_DFFPOSX1_608 ( );
FILL FILL_4_DFFPOSX1_608 ( );
FILL FILL_5_DFFPOSX1_608 ( );
FILL FILL_0_OAI21X1_754 ( );
FILL FILL_1_OAI21X1_754 ( );
FILL FILL_0_OAI21X1_753 ( );
FILL FILL_1_OAI21X1_753 ( );
FILL FILL_0_INVX1_29 ( );
FILL FILL_0_BUFX2_534 ( );
FILL FILL_0_DFFPOSX1_393 ( );
FILL FILL_1_DFFPOSX1_393 ( );
FILL FILL_2_DFFPOSX1_393 ( );
FILL FILL_3_DFFPOSX1_393 ( );
FILL FILL_4_DFFPOSX1_393 ( );
FILL FILL_5_DFFPOSX1_393 ( );
FILL FILL_6_DFFPOSX1_393 ( );
FILL FILL_0_BUFX2_482 ( );
FILL FILL_0_AND2X2_5 ( );
FILL FILL_1_AND2X2_5 ( );
FILL FILL_0_INVX1_10 ( );
FILL FILL_0_OAI21X1_424 ( );
FILL FILL_1_OAI21X1_424 ( );
FILL FILL_0_OAI21X1_427 ( );
FILL FILL_1_OAI21X1_427 ( );
FILL FILL_0_NAND2X1_278 ( );
FILL FILL_1_NAND2X1_278 ( );
FILL FILL_0_AND2X2_4 ( );
FILL FILL_1_AND2X2_4 ( );
FILL FILL_0_NAND2X1_186 ( );
FILL FILL_0_NOR2X1_16 ( );
FILL FILL_1_NOR2X1_16 ( );
FILL FILL_0_CLKBUF1_33 ( );
FILL FILL_1_CLKBUF1_33 ( );
FILL FILL_2_CLKBUF1_33 ( );
FILL FILL_3_CLKBUF1_33 ( );
FILL FILL_4_CLKBUF1_33 ( );
FILL FILL_0_INVX4_12 ( );
FILL FILL_0_OAI21X1_355 ( );
FILL FILL_1_OAI21X1_355 ( );
FILL FILL_0_NAND2X1_194 ( );
FILL FILL_1_NAND2X1_194 ( );
FILL FILL_0_NOR2X1_19 ( );
FILL FILL_0_NOR2X1_70 ( );
FILL FILL_1_NOR2X1_70 ( );
FILL FILL_0_INVX2_24 ( );
FILL FILL_0_OAI21X1_573 ( );
FILL FILL_1_OAI21X1_573 ( );
FILL FILL_0_NAND2X1_102 ( );
FILL FILL_1_NAND2X1_102 ( );
FILL FILL_0_NAND2X1_195 ( );
FILL FILL_1_NAND2X1_195 ( );
FILL FILL_0_DFFPOSX1_386 ( );
FILL FILL_1_DFFPOSX1_386 ( );
FILL FILL_2_DFFPOSX1_386 ( );
FILL FILL_3_DFFPOSX1_386 ( );
FILL FILL_4_DFFPOSX1_386 ( );
FILL FILL_5_DFFPOSX1_386 ( );
FILL FILL_6_DFFPOSX1_386 ( );
FILL FILL_0_INVX1_14 ( );
FILL FILL_0_XNOR2X1_10 ( );
FILL FILL_1_XNOR2X1_10 ( );
FILL FILL_2_XNOR2X1_10 ( );
FILL FILL_3_XNOR2X1_10 ( );
FILL FILL_0_OAI21X1_551 ( );
FILL FILL_1_OAI21X1_551 ( );
FILL FILL_0_OAI21X1_357 ( );
FILL FILL_1_OAI21X1_357 ( );
FILL FILL_0_BUFX2_204 ( );
FILL FILL_0_DFFPOSX1_385 ( );
FILL FILL_1_DFFPOSX1_385 ( );
FILL FILL_2_DFFPOSX1_385 ( );
FILL FILL_3_DFFPOSX1_385 ( );
FILL FILL_4_DFFPOSX1_385 ( );
FILL FILL_5_DFFPOSX1_385 ( );
FILL FILL_0_OAI21X1_1017 ( );
FILL FILL_1_OAI21X1_1017 ( );
FILL FILL_0_OAI21X1_1016 ( );
FILL FILL_1_OAI21X1_1016 ( );
FILL FILL_2_OAI21X1_1016 ( );
FILL FILL_0_OAI21X1_281 ( );
FILL FILL_1_OAI21X1_281 ( );
FILL FILL_0_DFFPOSX1_332 ( );
FILL FILL_1_DFFPOSX1_332 ( );
FILL FILL_2_DFFPOSX1_332 ( );
FILL FILL_3_DFFPOSX1_332 ( );
FILL FILL_4_DFFPOSX1_332 ( );
FILL FILL_5_DFFPOSX1_332 ( );
FILL FILL_6_DFFPOSX1_332 ( );
FILL FILL_0_OAI21X1_280 ( );
FILL FILL_1_OAI21X1_280 ( );
FILL FILL_0_OAI21X1_220 ( );
FILL FILL_1_OAI21X1_220 ( );
FILL FILL_2_OAI21X1_220 ( );
FILL FILL_0_OAI21X1_1275 ( );
FILL FILL_1_OAI21X1_1275 ( );
FILL FILL_0_INVX1_175 ( );
FILL FILL_0_INVX1_173 ( );
FILL FILL_0_BUFX4_4 ( );
FILL FILL_1_BUFX4_4 ( );
FILL FILL_0_NAND2X1_505 ( );
FILL FILL_0_NOR2X1_135 ( );
FILL FILL_1_NOR2X1_135 ( );
FILL FILL_0_INVX2_70 ( );
FILL FILL_1_INVX2_70 ( );
FILL FILL_0_OAI21X1_1447 ( );
FILL FILL_1_OAI21X1_1447 ( );
FILL FILL_0_DFFPOSX1_957 ( );
FILL FILL_1_DFFPOSX1_957 ( );
FILL FILL_2_DFFPOSX1_957 ( );
FILL FILL_3_DFFPOSX1_957 ( );
FILL FILL_4_DFFPOSX1_957 ( );
FILL FILL_5_DFFPOSX1_957 ( );
FILL FILL_0_OAI21X1_1446 ( );
FILL FILL_1_OAI21X1_1446 ( );
FILL FILL_2_OAI21X1_1446 ( );
FILL FILL_0_BUFX4_169 ( );
FILL FILL_1_BUFX4_169 ( );
FILL FILL_0_BUFX4_78 ( );
FILL FILL_1_BUFX4_78 ( );
FILL FILL_0_OAI21X1_1452 ( );
FILL FILL_1_OAI21X1_1452 ( );
FILL FILL_0_OAI21X1_1073 ( );
FILL FILL_1_OAI21X1_1073 ( );
FILL FILL_0_OAI21X1_1015 ( );
FILL FILL_1_OAI21X1_1015 ( );
FILL FILL_0_DFFPOSX1_910 ( );
FILL FILL_1_DFFPOSX1_910 ( );
FILL FILL_2_DFFPOSX1_910 ( );
FILL FILL_3_DFFPOSX1_910 ( );
FILL FILL_4_DFFPOSX1_910 ( );
FILL FILL_5_DFFPOSX1_910 ( );
FILL FILL_6_DFFPOSX1_910 ( );
FILL FILL_0_BUFX2_143 ( );
FILL FILL_1_BUFX2_143 ( );
FILL FILL_0_BUFX2_224 ( );
FILL FILL_1_BUFX2_224 ( );
FILL FILL_0_BUFX2_96 ( );
FILL FILL_1_BUFX2_96 ( );
FILL FILL_0_OAI21X1_1307 ( );
FILL FILL_1_OAI21X1_1307 ( );
FILL FILL_0_OAI21X1_1306 ( );
FILL FILL_1_OAI21X1_1306 ( );
FILL FILL_0_NAND2X1_539 ( );
FILL FILL_1_NAND2X1_539 ( );
FILL FILL_0_NAND2X1_540 ( );
FILL FILL_1_NAND2X1_540 ( );
FILL FILL_0_INVX4_41 ( );
FILL FILL_1_INVX4_41 ( );
FILL FILL_0_INVX2_78 ( );
FILL FILL_0_NAND2X1_609 ( );
FILL FILL_1_NAND2X1_609 ( );
FILL FILL_0_NAND2X1_536 ( );
FILL FILL_0_XNOR2X1_82 ( );
FILL FILL_1_XNOR2X1_82 ( );
FILL FILL_2_XNOR2X1_82 ( );
FILL FILL_0_NAND2X1_541 ( );
FILL FILL_1_NAND2X1_541 ( );
FILL FILL_0_OAI21X1_1320 ( );
FILL FILL_1_OAI21X1_1320 ( );
FILL FILL_0_OAI21X1_1322 ( );
FILL FILL_1_OAI21X1_1322 ( );
FILL FILL_0_OAI21X1_1321 ( );
FILL FILL_1_OAI21X1_1321 ( );
FILL FILL_0_DFFPOSX1_989 ( );
FILL FILL_1_DFFPOSX1_989 ( );
FILL FILL_2_DFFPOSX1_989 ( );
FILL FILL_3_DFFPOSX1_989 ( );
FILL FILL_4_DFFPOSX1_989 ( );
FILL FILL_5_DFFPOSX1_989 ( );
FILL FILL_0_OAI21X1_1546 ( );
FILL FILL_1_OAI21X1_1546 ( );
FILL FILL_0_BUFX2_241 ( );
FILL FILL_0_OAI21X1_1088 ( );
FILL FILL_1_OAI21X1_1088 ( );
FILL FILL_2_OAI21X1_1088 ( );
FILL FILL_0_OAI21X1_1370 ( );
FILL FILL_1_OAI21X1_1370 ( );
FILL FILL_0_OAI21X1_1544 ( );
FILL FILL_1_OAI21X1_1544 ( );
FILL FILL_0_NAND2X1_572 ( );
FILL FILL_0_OAI21X1_1184 ( );
FILL FILL_1_OAI21X1_1184 ( );
FILL FILL_2_OAI21X1_1184 ( );
FILL FILL_0_OAI21X1_1185 ( );
FILL FILL_1_OAI21X1_1185 ( );
FILL FILL_0_OAI21X1_1186 ( );
FILL FILL_1_OAI21X1_1186 ( );
FILL FILL_0_OAI21X1_1187 ( );
FILL FILL_1_OAI21X1_1187 ( );
FILL FILL_2_OAI21X1_1187 ( );
FILL FILL_0_INVX4_48 ( );
FILL FILL_0_OAI21X1_1188 ( );
FILL FILL_1_OAI21X1_1188 ( );
FILL FILL_0_NAND3X1_48 ( );
FILL FILL_1_NAND3X1_48 ( );
FILL FILL_0_OAI21X1_1357 ( );
FILL FILL_1_OAI21X1_1357 ( );
FILL FILL_0_OAI21X1_1547 ( );
FILL FILL_1_OAI21X1_1547 ( );
FILL FILL_0_XNOR2X1_86 ( );
FILL FILL_1_XNOR2X1_86 ( );
FILL FILL_2_XNOR2X1_86 ( );
FILL FILL_3_XNOR2X1_86 ( );
FILL FILL_0_INVX1_180 ( );
FILL FILL_0_INVX2_104 ( );
FILL FILL_0_OAI21X1_1556 ( );
FILL FILL_1_OAI21X1_1556 ( );
FILL FILL_0_DFFPOSX1_799 ( );
FILL FILL_1_DFFPOSX1_799 ( );
FILL FILL_2_DFFPOSX1_799 ( );
FILL FILL_3_DFFPOSX1_799 ( );
FILL FILL_4_DFFPOSX1_799 ( );
FILL FILL_5_DFFPOSX1_799 ( );
FILL FILL_0_OAI21X1_1553 ( );
FILL FILL_1_OAI21X1_1553 ( );
FILL FILL_0_CLKBUF1_20 ( );
FILL FILL_1_CLKBUF1_20 ( );
FILL FILL_2_CLKBUF1_20 ( );
FILL FILL_3_CLKBUF1_20 ( );
FILL FILL_4_CLKBUF1_20 ( );
FILL FILL_0_BUFX2_52 ( );
FILL FILL_1_BUFX2_52 ( );
FILL FILL_0_BUFX2_180 ( );
FILL FILL_1_BUFX2_180 ( );
FILL FILL_0_OAI21X1_1349 ( );
FILL FILL_1_OAI21X1_1349 ( );
FILL FILL_2_OAI21X1_1349 ( );
FILL FILL_0_DFFPOSX1_923 ( );
FILL FILL_1_DFFPOSX1_923 ( );
FILL FILL_2_DFFPOSX1_923 ( );
FILL FILL_3_DFFPOSX1_923 ( );
FILL FILL_4_DFFPOSX1_923 ( );
FILL FILL_5_DFFPOSX1_923 ( );
FILL FILL_6_DFFPOSX1_923 ( );
FILL FILL_0_OAI21X1_1348 ( );
FILL FILL_1_OAI21X1_1348 ( );
FILL FILL_0_BUFX2_59 ( );
FILL FILL_0_DFFPOSX1_279 ( );
FILL FILL_1_DFFPOSX1_279 ( );
FILL FILL_2_DFFPOSX1_279 ( );
FILL FILL_3_DFFPOSX1_279 ( );
FILL FILL_4_DFFPOSX1_279 ( );
FILL FILL_5_DFFPOSX1_279 ( );
FILL FILL_0_OAI21X1_175 ( );
FILL FILL_1_OAI21X1_175 ( );
FILL FILL_2_OAI21X1_175 ( );
FILL FILL_0_OAI21X1_174 ( );
FILL FILL_1_OAI21X1_174 ( );
FILL FILL_0_BUFX2_735 ( );
FILL FILL_0_NAND2X1_711 ( );
FILL FILL_1_NAND2X1_711 ( );
FILL FILL_0_OAI21X1_49 ( );
FILL FILL_1_OAI21X1_49 ( );
FILL FILL_0_NAND2X1_49 ( );
FILL FILL_1_NAND2X1_49 ( );
FILL FILL_0_DFFPOSX1_205 ( );
FILL FILL_1_DFFPOSX1_205 ( );
FILL FILL_2_DFFPOSX1_205 ( );
FILL FILL_3_DFFPOSX1_205 ( );
FILL FILL_4_DFFPOSX1_205 ( );
FILL FILL_5_DFFPOSX1_205 ( );
FILL FILL_0_BUFX2_703 ( );
FILL FILL_0_INVX1_128 ( );
FILL FILL_0_DFFPOSX1_652 ( );
FILL FILL_1_DFFPOSX1_652 ( );
FILL FILL_2_DFFPOSX1_652 ( );
FILL FILL_3_DFFPOSX1_652 ( );
FILL FILL_4_DFFPOSX1_652 ( );
FILL FILL_5_DFFPOSX1_652 ( );
FILL FILL_0_INVX2_192 ( );
FILL FILL_0_DFFPOSX1_162 ( );
FILL FILL_1_DFFPOSX1_162 ( );
FILL FILL_2_DFFPOSX1_162 ( );
FILL FILL_3_DFFPOSX1_162 ( );
FILL FILL_4_DFFPOSX1_162 ( );
FILL FILL_5_DFFPOSX1_162 ( );
FILL FILL_0_NAND2X1_6 ( );
FILL FILL_0_OAI21X1_6 ( );
FILL FILL_1_OAI21X1_6 ( );
FILL FILL_2_OAI21X1_6 ( );
FILL FILL_0_BUFX2_1010 ( );
FILL FILL_0_NAND2X1_761 ( );
FILL FILL_1_NAND2X1_761 ( );
FILL FILL_0_OAI21X1_1820 ( );
FILL FILL_1_OAI21X1_1820 ( );
FILL FILL_0_DFFPOSX1_210 ( );
FILL FILL_1_DFFPOSX1_210 ( );
FILL FILL_2_DFFPOSX1_210 ( );
FILL FILL_3_DFFPOSX1_210 ( );
FILL FILL_4_DFFPOSX1_210 ( );
FILL FILL_5_DFFPOSX1_210 ( );
FILL FILL_0_OAI21X1_54 ( );
FILL FILL_1_OAI21X1_54 ( );
FILL FILL_2_OAI21X1_54 ( );
FILL FILL_0_NAND2X1_54 ( );
FILL FILL_0_BUFX4_327 ( );
FILL FILL_1_BUFX4_327 ( );
FILL FILL_0_CLKBUF1_41 ( );
FILL FILL_1_CLKBUF1_41 ( );
FILL FILL_2_CLKBUF1_41 ( );
FILL FILL_3_CLKBUF1_41 ( );
FILL FILL_4_CLKBUF1_41 ( );
FILL FILL_0_BUFX4_222 ( );
FILL FILL_1_BUFX4_222 ( );
FILL FILL_2_BUFX4_222 ( );
FILL FILL_0_BUFX2_619 ( );
FILL FILL_1_BUFX2_619 ( );
FILL FILL_0_DFFPOSX1_489 ( );
FILL FILL_1_DFFPOSX1_489 ( );
FILL FILL_2_DFFPOSX1_489 ( );
FILL FILL_3_DFFPOSX1_489 ( );
FILL FILL_4_DFFPOSX1_489 ( );
FILL FILL_5_DFFPOSX1_489 ( );
FILL FILL_0_OAI21X1_514 ( );
FILL FILL_1_OAI21X1_514 ( );
FILL FILL_0_OAI21X1_515 ( );
FILL FILL_1_OAI21X1_515 ( );
FILL FILL_0_INVX1_24 ( );
FILL FILL_0_OAI21X1_506 ( );
FILL FILL_1_OAI21X1_506 ( );
FILL FILL_0_OAI21X1_510 ( );
FILL FILL_1_OAI21X1_510 ( );
FILL FILL_0_NOR2X1_59 ( );
FILL FILL_1_NOR2X1_59 ( );
FILL FILL_0_OAI21X1_513 ( );
FILL FILL_1_OAI21X1_513 ( );
FILL FILL_0_NAND2X1_718 ( );
FILL FILL_1_NAND2X1_718 ( );
FILL FILL_0_OAI21X1_1777 ( );
FILL FILL_1_OAI21X1_1777 ( );
FILL FILL_0_DFFPOSX1_103 ( );
FILL FILL_1_DFFPOSX1_103 ( );
FILL FILL_2_DFFPOSX1_103 ( );
FILL FILL_3_DFFPOSX1_103 ( );
FILL FILL_4_DFFPOSX1_103 ( );
FILL FILL_5_DFFPOSX1_103 ( );
FILL FILL_0_DFFPOSX1_368 ( );
FILL FILL_1_DFFPOSX1_368 ( );
FILL FILL_2_DFFPOSX1_368 ( );
FILL FILL_3_DFFPOSX1_368 ( );
FILL FILL_4_DFFPOSX1_368 ( );
FILL FILL_5_DFFPOSX1_368 ( );
FILL FILL_0_NAND2X1_84 ( );
FILL FILL_1_NAND2X1_84 ( );
FILL FILL_0_OAI21X1_340 ( );
FILL FILL_1_OAI21X1_340 ( );
FILL FILL_0_OAI21X1_537 ( );
FILL FILL_1_OAI21X1_537 ( );
FILL FILL_0_OAI21X1_701 ( );
FILL FILL_1_OAI21X1_701 ( );
FILL FILL_0_DFFPOSX1_497 ( );
FILL FILL_1_DFFPOSX1_497 ( );
FILL FILL_2_DFFPOSX1_497 ( );
FILL FILL_3_DFFPOSX1_497 ( );
FILL FILL_4_DFFPOSX1_497 ( );
FILL FILL_5_DFFPOSX1_497 ( );
FILL FILL_6_DFFPOSX1_497 ( );
FILL FILL_0_OAI21X1_538 ( );
FILL FILL_1_OAI21X1_538 ( );
FILL FILL_0_NAND2X1_274 ( );
FILL FILL_1_NAND2X1_274 ( );
FILL FILL_0_OAI21X1_543 ( );
FILL FILL_1_OAI21X1_543 ( );
FILL FILL_0_OAI21X1_542 ( );
FILL FILL_1_OAI21X1_542 ( );
FILL FILL_0_OAI22X1_1 ( );
FILL FILL_1_OAI22X1_1 ( );
FILL FILL_2_OAI22X1_1 ( );
FILL FILL_0_NAND2X1_273 ( );
FILL FILL_1_NAND2X1_273 ( );
FILL FILL_0_NOR2X1_61 ( );
FILL FILL_0_NAND2X1_275 ( );
FILL FILL_1_NAND2X1_275 ( );
FILL FILL_0_BUFX4_167 ( );
FILL FILL_1_BUFX4_167 ( );
FILL FILL_0_XNOR2X1_26 ( );
FILL FILL_1_XNOR2X1_26 ( );
FILL FILL_2_XNOR2X1_26 ( );
FILL FILL_3_XNOR2X1_26 ( );
FILL FILL_0_OAI21X1_536 ( );
FILL FILL_1_OAI21X1_536 ( );
FILL FILL_2_OAI21X1_536 ( );
FILL FILL_0_NOR2X1_11 ( );
FILL FILL_0_NOR2X1_105 ( );
FILL FILL_1_NOR2X1_105 ( );
FILL FILL_0_AND2X2_8 ( );
FILL FILL_1_AND2X2_8 ( );
FILL FILL_0_OAI21X1_376 ( );
FILL FILL_1_OAI21X1_376 ( );
FILL FILL_0_BUFX4_345 ( );
FILL FILL_1_BUFX4_345 ( );
FILL FILL_0_NAND2X1_225 ( );
FILL FILL_0_NAND2X1_244 ( );
FILL FILL_0_BUFX2_561 ( );
FILL FILL_1_BUFX2_561 ( );
FILL FILL_0_INVX2_36 ( );
FILL FILL_1_INVX2_36 ( );
FILL FILL_0_AOI21X1_3 ( );
FILL FILL_1_AOI21X1_3 ( );
FILL FILL_2_AOI21X1_3 ( );
FILL FILL_0_INVX1_20 ( );
FILL FILL_0_NOR2X1_49 ( );
FILL FILL_1_NOR2X1_49 ( );
FILL FILL_0_BUFX2_635 ( );
FILL FILL_1_BUFX2_635 ( );
FILL FILL_0_NAND2X1_316 ( );
FILL FILL_1_NAND2X1_316 ( );
FILL FILL_0_DFFPOSX1_410 ( );
FILL FILL_1_DFFPOSX1_410 ( );
FILL FILL_2_DFFPOSX1_410 ( );
FILL FILL_3_DFFPOSX1_410 ( );
FILL FILL_4_DFFPOSX1_410 ( );
FILL FILL_5_DFFPOSX1_410 ( );
FILL FILL_6_DFFPOSX1_410 ( );
FILL FILL_0_DFFPOSX1_419 ( );
FILL FILL_1_DFFPOSX1_419 ( );
FILL FILL_2_DFFPOSX1_419 ( );
FILL FILL_3_DFFPOSX1_419 ( );
FILL FILL_4_DFFPOSX1_419 ( );
FILL FILL_5_DFFPOSX1_419 ( );
FILL FILL_6_DFFPOSX1_419 ( );
FILL FILL_0_DFFPOSX1_524 ( );
FILL FILL_1_DFFPOSX1_524 ( );
FILL FILL_2_DFFPOSX1_524 ( );
FILL FILL_3_DFFPOSX1_524 ( );
FILL FILL_4_DFFPOSX1_524 ( );
FILL FILL_5_DFFPOSX1_524 ( );
FILL FILL_0_NOR2X1_25 ( );
FILL FILL_0_INVX2_43 ( );
FILL FILL_0_INVX2_25 ( );
FILL FILL_0_DFFPOSX1_523 ( );
FILL FILL_1_DFFPOSX1_523 ( );
FILL FILL_2_DFFPOSX1_523 ( );
FILL FILL_3_DFFPOSX1_523 ( );
FILL FILL_4_DFFPOSX1_523 ( );
FILL FILL_5_DFFPOSX1_523 ( );
FILL FILL_6_DFFPOSX1_523 ( );
FILL FILL_0_OAI21X1_604 ( );
FILL FILL_1_OAI21X1_604 ( );
FILL FILL_2_OAI21X1_604 ( );
FILL FILL_0_CLKBUF1_44 ( );
FILL FILL_1_CLKBUF1_44 ( );
FILL FILL_2_CLKBUF1_44 ( );
FILL FILL_3_CLKBUF1_44 ( );
FILL FILL_4_CLKBUF1_44 ( );
FILL FILL_0_NAND2X1_109 ( );
FILL FILL_0_OAI21X1_365 ( );
FILL FILL_1_OAI21X1_365 ( );
FILL FILL_0_OAI21X1_423 ( );
FILL FILL_1_OAI21X1_423 ( );
FILL FILL_0_DFFPOSX1_569 ( );
FILL FILL_1_DFFPOSX1_569 ( );
FILL FILL_2_DFFPOSX1_569 ( );
FILL FILL_3_DFFPOSX1_569 ( );
FILL FILL_4_DFFPOSX1_569 ( );
FILL FILL_5_DFFPOSX1_569 ( );
FILL FILL_0_NOR2X1_12 ( );
FILL FILL_1_NOR2X1_12 ( );
FILL FILL_0_NAND3X1_4 ( );
FILL FILL_1_NAND3X1_4 ( );
FILL FILL_0_NAND2X1_174 ( );
FILL FILL_1_NAND2X1_174 ( );
FILL FILL_0_NAND2X1_182 ( );
FILL FILL_0_NOR2X1_27 ( );
FILL FILL_1_NOR2X1_27 ( );
FILL FILL_0_OR2X2_3 ( );
FILL FILL_1_OR2X2_3 ( );
FILL FILL_0_NOR2X1_68 ( );
FILL FILL_1_NOR2X1_68 ( );
FILL FILL_0_CLKBUF1_18 ( );
FILL FILL_1_CLKBUF1_18 ( );
FILL FILL_2_CLKBUF1_18 ( );
FILL FILL_3_CLKBUF1_18 ( );
FILL FILL_4_CLKBUF1_18 ( );
FILL FILL_0_NAND3X1_3 ( );
FILL FILL_1_NAND3X1_3 ( );
FILL FILL_0_NAND2X1_281 ( );
FILL FILL_1_NAND2X1_281 ( );
FILL FILL_0_NAND2X1_199 ( );
FILL FILL_1_NAND2X1_199 ( );
FILL FILL_0_AOI21X1_1 ( );
FILL FILL_1_AOI21X1_1 ( );
FILL FILL_0_NAND2X1_283 ( );
FILL FILL_1_NAND2X1_283 ( );
FILL FILL_0_INVX2_42 ( );
FILL FILL_0_INVX4_10 ( );
FILL FILL_1_INVX4_10 ( );
FILL FILL_0_NOR2X1_17 ( );
FILL FILL_0_OAI21X1_447 ( );
FILL FILL_1_OAI21X1_447 ( );
FILL FILL_0_OAI21X1_358 ( );
FILL FILL_1_OAI21X1_358 ( );
FILL FILL_0_OAI21X1_552 ( );
FILL FILL_1_OAI21X1_552 ( );
FILL FILL_0_DFFPOSX1_502 ( );
FILL FILL_1_DFFPOSX1_502 ( );
FILL FILL_2_DFFPOSX1_502 ( );
FILL FILL_3_DFFPOSX1_502 ( );
FILL FILL_4_DFFPOSX1_502 ( );
FILL FILL_5_DFFPOSX1_502 ( );
FILL FILL_0_DFFPOSX1_451 ( );
FILL FILL_1_DFFPOSX1_451 ( );
FILL FILL_2_DFFPOSX1_451 ( );
FILL FILL_3_DFFPOSX1_451 ( );
FILL FILL_4_DFFPOSX1_451 ( );
FILL FILL_5_DFFPOSX1_451 ( );
FILL FILL_6_DFFPOSX1_451 ( );
FILL FILL_0_DFFPOSX1_734 ( );
FILL FILL_1_DFFPOSX1_734 ( );
FILL FILL_2_DFFPOSX1_734 ( );
FILL FILL_3_DFFPOSX1_734 ( );
FILL FILL_4_DFFPOSX1_734 ( );
FILL FILL_5_DFFPOSX1_734 ( );
FILL FILL_0_DFFPOSX1_302 ( );
FILL FILL_1_DFFPOSX1_302 ( );
FILL FILL_2_DFFPOSX1_302 ( );
FILL FILL_3_DFFPOSX1_302 ( );
FILL FILL_4_DFFPOSX1_302 ( );
FILL FILL_5_DFFPOSX1_302 ( );
FILL FILL_6_DFFPOSX1_302 ( );
FILL FILL_0_OAI21X1_221 ( );
FILL FILL_1_OAI21X1_221 ( );
FILL FILL_0_OAI21X1_1443 ( );
FILL FILL_1_OAI21X1_1443 ( );
FILL FILL_0_OAI21X1_1444 ( );
FILL FILL_1_OAI21X1_1444 ( );
FILL FILL_2_OAI21X1_1444 ( );
FILL FILL_0_OAI21X1_1445 ( );
FILL FILL_1_OAI21X1_1445 ( );
FILL FILL_0_NAND2X1_629 ( );
FILL FILL_0_INVX1_222 ( );
FILL FILL_0_XNOR2X1_94 ( );
FILL FILL_1_XNOR2X1_94 ( );
FILL FILL_2_XNOR2X1_94 ( );
FILL FILL_0_OAI21X1_1448 ( );
FILL FILL_1_OAI21X1_1448 ( );
FILL FILL_0_INVX4_36 ( );
FILL FILL_1_INVX4_36 ( );
FILL FILL_0_DFFPOSX1_895 ( );
FILL FILL_1_DFFPOSX1_895 ( );
FILL FILL_2_DFFPOSX1_895 ( );
FILL FILL_3_DFFPOSX1_895 ( );
FILL FILL_4_DFFPOSX1_895 ( );
FILL FILL_5_DFFPOSX1_895 ( );
FILL FILL_6_DFFPOSX1_895 ( );
FILL FILL_0_DFFPOSX1_959 ( );
FILL FILL_1_DFFPOSX1_959 ( );
FILL FILL_2_DFFPOSX1_959 ( );
FILL FILL_3_DFFPOSX1_959 ( );
FILL FILL_4_DFFPOSX1_959 ( );
FILL FILL_5_DFFPOSX1_959 ( );
FILL FILL_0_DFFPOSX1_733 ( );
FILL FILL_1_DFFPOSX1_733 ( );
FILL FILL_2_DFFPOSX1_733 ( );
FILL FILL_3_DFFPOSX1_733 ( );
FILL FILL_4_DFFPOSX1_733 ( );
FILL FILL_5_DFFPOSX1_733 ( );
FILL FILL_6_DFFPOSX1_733 ( );
FILL FILL_0_OAI21X1_1266 ( );
FILL FILL_1_OAI21X1_1266 ( );
FILL FILL_2_OAI21X1_1266 ( );
FILL FILL_0_BUFX4_370 ( );
FILL FILL_1_BUFX4_370 ( );
FILL FILL_0_OAI21X1_1310 ( );
FILL FILL_1_OAI21X1_1310 ( );
FILL FILL_0_OAI21X1_1312 ( );
FILL FILL_1_OAI21X1_1312 ( );
FILL FILL_0_OAI21X1_1313 ( );
FILL FILL_1_OAI21X1_1313 ( );
FILL FILL_0_NAND2X1_611 ( );
FILL FILL_1_NAND2X1_611 ( );
FILL FILL_0_XNOR2X1_69 ( );
FILL FILL_1_XNOR2X1_69 ( );
FILL FILL_2_XNOR2X1_69 ( );
FILL FILL_0_NOR2X1_156 ( );
FILL FILL_1_NOR2X1_156 ( );
FILL FILL_0_NOR2X1_199 ( );
FILL FILL_0_OAI21X1_1497 ( );
FILL FILL_1_OAI21X1_1497 ( );
FILL FILL_0_OAI21X1_1489 ( );
FILL FILL_1_OAI21X1_1489 ( );
FILL FILL_0_NOR2X1_154 ( );
FILL FILL_1_NOR2X1_154 ( );
FILL FILL_0_NOR2X1_155 ( );
FILL FILL_0_OAI21X1_1486 ( );
FILL FILL_1_OAI21X1_1486 ( );
FILL FILL_0_NOR2X1_159 ( );
FILL FILL_1_NOR2X1_159 ( );
FILL FILL_0_NAND3X1_44 ( );
FILL FILL_1_NAND3X1_44 ( );
FILL FILL_0_NAND2X1_612 ( );
FILL FILL_1_NAND2X1_612 ( );
FILL FILL_0_AOI21X1_50 ( );
FILL FILL_1_AOI21X1_50 ( );
FILL FILL_0_INVX2_101 ( );
FILL FILL_0_BUFX4_6 ( );
FILL FILL_1_BUFX4_6 ( );
FILL FILL_0_DFFPOSX1_987 ( );
FILL FILL_1_DFFPOSX1_987 ( );
FILL FILL_2_DFFPOSX1_987 ( );
FILL FILL_3_DFFPOSX1_987 ( );
FILL FILL_4_DFFPOSX1_987 ( );
FILL FILL_5_DFFPOSX1_987 ( );
FILL FILL_0_OAI21X1_1539 ( );
FILL FILL_1_OAI21X1_1539 ( );
FILL FILL_0_OAI21X1_1543 ( );
FILL FILL_1_OAI21X1_1543 ( );
FILL FILL_0_OAI21X1_1537 ( );
FILL FILL_1_OAI21X1_1537 ( );
FILL FILL_2_OAI21X1_1537 ( );
FILL FILL_0_NAND2X1_571 ( );
FILL FILL_0_OAI21X1_1536 ( );
FILL FILL_1_OAI21X1_1536 ( );
FILL FILL_0_INVX2_84 ( );
FILL FILL_0_OAI21X1_1182 ( );
FILL FILL_1_OAI21X1_1182 ( );
FILL FILL_0_NOR3X1_13 ( );
FILL FILL_1_NOR3X1_13 ( );
FILL FILL_2_NOR3X1_13 ( );
FILL FILL_3_NOR3X1_13 ( );
FILL FILL_0_NAND2X1_568 ( );
FILL FILL_0_NOR2X1_169 ( );
FILL FILL_1_NOR2X1_169 ( );
FILL FILL_0_AOI21X1_56 ( );
FILL FILL_1_AOI21X1_56 ( );
FILL FILL_0_NOR2X1_172 ( );
FILL FILL_1_NOR2X1_172 ( );
FILL FILL_0_NOR2X1_229 ( );
FILL FILL_0_NOR3X1_14 ( );
FILL FILL_1_NOR3X1_14 ( );
FILL FILL_2_NOR3X1_14 ( );
FILL FILL_3_NOR3X1_14 ( );
FILL FILL_4_NOR3X1_14 ( );
FILL FILL_0_NAND2X1_643 ( );
FILL FILL_1_NAND2X1_643 ( );
FILL FILL_0_INVX2_87 ( );
FILL FILL_1_INVX2_87 ( );
FILL FILL_0_INVX2_86 ( );
FILL FILL_0_OAI21X1_1557 ( );
FILL FILL_1_OAI21X1_1557 ( );
FILL FILL_2_OAI21X1_1557 ( );
FILL FILL_0_INVX1_227 ( );
FILL FILL_0_DFFPOSX1_993 ( );
FILL FILL_1_DFFPOSX1_993 ( );
FILL FILL_2_DFFPOSX1_993 ( );
FILL FILL_3_DFFPOSX1_993 ( );
FILL FILL_4_DFFPOSX1_993 ( );
FILL FILL_5_DFFPOSX1_993 ( );
FILL FILL_6_DFFPOSX1_993 ( );
FILL FILL_0_OAI21X1_1091 ( );
FILL FILL_1_OAI21X1_1091 ( );
FILL FILL_0_NAND2X1_457 ( );
FILL FILL_1_NAND2X1_457 ( );
FILL FILL_0_OAI21X1_1097 ( );
FILL FILL_1_OAI21X1_1097 ( );
FILL FILL_0_NAND2X1_463 ( );
FILL FILL_1_NAND2X1_463 ( );
FILL FILL_0_DFFPOSX1_805 ( );
FILL FILL_1_DFFPOSX1_805 ( );
FILL FILL_2_DFFPOSX1_805 ( );
FILL FILL_3_DFFPOSX1_805 ( );
FILL FILL_4_DFFPOSX1_805 ( );
FILL FILL_5_DFFPOSX1_805 ( );
FILL FILL_0_BUFX4_331 ( );
FILL FILL_1_BUFX4_331 ( );
FILL FILL_0_BUFX4_144 ( );
FILL FILL_1_BUFX4_144 ( );
FILL FILL_2_BUFX4_144 ( );
FILL FILL_0_OAI21X1_1089 ( );
FILL FILL_1_OAI21X1_1089 ( );
FILL FILL_0_NAND2X1_455 ( );
FILL FILL_0_DFFPOSX1_797 ( );
FILL FILL_1_DFFPOSX1_797 ( );
FILL FILL_2_DFFPOSX1_797 ( );
FILL FILL_3_DFFPOSX1_797 ( );
FILL FILL_4_DFFPOSX1_797 ( );
FILL FILL_5_DFFPOSX1_797 ( );
FILL FILL_0_OAI21X1_1643 ( );
FILL FILL_1_OAI21X1_1643 ( );
FILL FILL_0_DFFPOSX1_33 ( );
FILL FILL_1_DFFPOSX1_33 ( );
FILL FILL_2_DFFPOSX1_33 ( );
FILL FILL_3_DFFPOSX1_33 ( );
FILL FILL_4_DFFPOSX1_33 ( );
FILL FILL_5_DFFPOSX1_33 ( );
FILL FILL_6_DFFPOSX1_33 ( );
FILL FILL_0_INVX1_125 ( );
FILL FILL_0_OAI21X1_1003 ( );
FILL FILL_1_OAI21X1_1003 ( );
FILL FILL_0_BUFX2_43 ( );
FILL FILL_0_INVX1_83 ( );
FILL FILL_0_BUFX2_964 ( );
FILL FILL_1_BUFX2_964 ( );
FILL FILL_0_BUFX2_946 ( );
FILL FILL_1_BUFX2_946 ( );
FILL FILL_0_BUFX2_480 ( );
FILL FILL_0_DFFPOSX1_354 ( );
FILL FILL_1_DFFPOSX1_354 ( );
FILL FILL_2_DFFPOSX1_354 ( );
FILL FILL_3_DFFPOSX1_354 ( );
FILL FILL_4_DFFPOSX1_354 ( );
FILL FILL_5_DFFPOSX1_354 ( );
FILL FILL_6_DFFPOSX1_354 ( );
FILL FILL_0_OAI21X1_325 ( );
FILL FILL_1_OAI21X1_325 ( );
FILL FILL_0_OAI21X1_324 ( );
FILL FILL_1_OAI21X1_324 ( );
FILL FILL_2_OAI21X1_324 ( );
FILL FILL_0_OAI21X1_292 ( );
FILL FILL_1_OAI21X1_292 ( );
FILL FILL_2_OAI21X1_292 ( );
FILL FILL_0_OAI21X1_293 ( );
FILL FILL_1_OAI21X1_293 ( );
FILL FILL_0_DFFPOSX1_338 ( );
FILL FILL_1_DFFPOSX1_338 ( );
FILL FILL_2_DFFPOSX1_338 ( );
FILL FILL_3_DFFPOSX1_338 ( );
FILL FILL_4_DFFPOSX1_338 ( );
FILL FILL_5_DFFPOSX1_338 ( );
FILL FILL_6_DFFPOSX1_338 ( );
FILL FILL_0_DFFPOSX1_300 ( );
FILL FILL_1_DFFPOSX1_300 ( );
FILL FILL_2_DFFPOSX1_300 ( );
FILL FILL_3_DFFPOSX1_300 ( );
FILL FILL_4_DFFPOSX1_300 ( );
FILL FILL_5_DFFPOSX1_300 ( );
FILL FILL_0_OAI21X1_217 ( );
FILL FILL_1_OAI21X1_217 ( );
FILL FILL_0_OAI21X1_216 ( );
FILL FILL_1_OAI21X1_216 ( );
FILL FILL_0_NAND2X1_142 ( );
FILL FILL_0_OAI21X1_399 ( );
FILL FILL_1_OAI21X1_399 ( );
FILL FILL_0_NAND2X1_141 ( );
FILL FILL_0_BUFX2_432 ( );
FILL FILL_1_BUFX2_432 ( );
FILL FILL_0_OAI21X1_670 ( );
FILL FILL_1_OAI21X1_670 ( );
FILL FILL_0_DFFPOSX1_552 ( );
FILL FILL_1_DFFPOSX1_552 ( );
FILL FILL_2_DFFPOSX1_552 ( );
FILL FILL_3_DFFPOSX1_552 ( );
FILL FILL_4_DFFPOSX1_552 ( );
FILL FILL_5_DFFPOSX1_552 ( );
FILL FILL_0_OAI21X1_671 ( );
FILL FILL_1_OAI21X1_671 ( );
FILL FILL_0_INVX2_10 ( );
FILL FILL_0_OAI21X1_509 ( );
FILL FILL_1_OAI21X1_509 ( );
FILL FILL_0_CLKBUF1_94 ( );
FILL FILL_1_CLKBUF1_94 ( );
FILL FILL_2_CLKBUF1_94 ( );
FILL FILL_3_CLKBUF1_94 ( );
FILL FILL_4_CLKBUF1_94 ( );
FILL FILL_0_DFFPOSX1_421 ( );
FILL FILL_1_DFFPOSX1_421 ( );
FILL FILL_2_DFFPOSX1_421 ( );
FILL FILL_3_DFFPOSX1_421 ( );
FILL FILL_4_DFFPOSX1_421 ( );
FILL FILL_5_DFFPOSX1_421 ( );
FILL FILL_6_DFFPOSX1_421 ( );
FILL FILL_0_INVX1_6 ( );
FILL FILL_1_INVX1_6 ( );
FILL FILL_0_OAI21X1_393 ( );
FILL FILL_1_OAI21X1_393 ( );
FILL FILL_0_BUFX2_441 ( );
FILL FILL_0_NAND2X1_138 ( );
FILL FILL_1_NAND2X1_138 ( );
FILL FILL_0_OAI21X1_547 ( );
FILL FILL_1_OAI21X1_547 ( );
FILL FILL_2_OAI21X1_547 ( );
FILL FILL_0_OAI21X1_548 ( );
FILL FILL_1_OAI21X1_548 ( );
FILL FILL_0_NAND2X1_118 ( );
FILL FILL_1_NAND2X1_118 ( );
FILL FILL_0_DFFPOSX1_495 ( );
FILL FILL_1_DFFPOSX1_495 ( );
FILL FILL_2_DFFPOSX1_495 ( );
FILL FILL_3_DFFPOSX1_495 ( );
FILL FILL_4_DFFPOSX1_495 ( );
FILL FILL_5_DFFPOSX1_495 ( );
FILL FILL_0_OAI21X1_533 ( );
FILL FILL_1_OAI21X1_533 ( );
FILL FILL_0_OAI21X1_534 ( );
FILL FILL_1_OAI21X1_534 ( );
FILL FILL_0_OAI21X1_695 ( );
FILL FILL_1_OAI21X1_695 ( );
FILL FILL_2_OAI21X1_695 ( );
FILL FILL_0_OAI21X1_694 ( );
FILL FILL_1_OAI21X1_694 ( );
FILL FILL_0_OAI21X1_593 ( );
FILL FILL_1_OAI21X1_593 ( );
FILL FILL_0_BUFX2_563 ( );
FILL FILL_0_DFFPOSX1_499 ( );
FILL FILL_1_DFFPOSX1_499 ( );
FILL FILL_2_DFFPOSX1_499 ( );
FILL FILL_3_DFFPOSX1_499 ( );
FILL FILL_4_DFFPOSX1_499 ( );
FILL FILL_5_DFFPOSX1_499 ( );
FILL FILL_6_DFFPOSX1_499 ( );
FILL FILL_0_BUFX2_433 ( );
FILL FILL_0_DFFPOSX1_401 ( );
FILL FILL_1_DFFPOSX1_401 ( );
FILL FILL_2_DFFPOSX1_401 ( );
FILL FILL_3_DFFPOSX1_401 ( );
FILL FILL_4_DFFPOSX1_401 ( );
FILL FILL_5_DFFPOSX1_401 ( );
FILL FILL_6_DFFPOSX1_401 ( );
FILL FILL_0_OAI21X1_535 ( );
FILL FILL_1_OAI21X1_535 ( );
FILL FILL_0_NAND2X1_117 ( );
FILL FILL_1_NAND2X1_117 ( );
FILL FILL_0_OAI21X1_373 ( );
FILL FILL_1_OAI21X1_373 ( );
FILL FILL_0_INVX1_33 ( );
FILL FILL_0_OAI21X1_619 ( );
FILL FILL_1_OAI21X1_619 ( );
FILL FILL_0_NOR2X1_88 ( );
FILL FILL_1_NOR2X1_88 ( );
FILL FILL_0_INVX2_50 ( );
FILL FILL_0_OAI21X1_616 ( );
FILL FILL_1_OAI21X1_616 ( );
FILL FILL_0_OAI21X1_617 ( );
FILL FILL_1_OAI21X1_617 ( );
FILL FILL_0_OAI21X1_615 ( );
FILL FILL_1_OAI21X1_615 ( );
FILL FILL_0_NOR2X1_48 ( );
FILL FILL_1_NOR2X1_48 ( );
FILL FILL_0_INVX1_3 ( );
FILL FILL_0_INVX2_46 ( );
FILL FILL_0_DFFPOSX1_529 ( );
FILL FILL_1_DFFPOSX1_529 ( );
FILL FILL_2_DFFPOSX1_529 ( );
FILL FILL_3_DFFPOSX1_529 ( );
FILL FILL_4_DFFPOSX1_529 ( );
FILL FILL_5_DFFPOSX1_529 ( );
FILL FILL_6_DFFPOSX1_529 ( );
FILL FILL_0_BUFX4_244 ( );
FILL FILL_1_BUFX4_244 ( );
FILL FILL_0_OAI21X1_382 ( );
FILL FILL_1_OAI21X1_382 ( );
FILL FILL_0_NAND2X1_126 ( );
FILL FILL_0_OAI21X1_599 ( );
FILL FILL_1_OAI21X1_599 ( );
FILL FILL_0_OAI21X1_391 ( );
FILL FILL_1_OAI21X1_391 ( );
FILL FILL_0_CLKBUF1_79 ( );
FILL FILL_1_CLKBUF1_79 ( );
FILL FILL_2_CLKBUF1_79 ( );
FILL FILL_3_CLKBUF1_79 ( );
FILL FILL_4_CLKBUF1_79 ( );
FILL FILL_0_AOI21X1_12 ( );
FILL FILL_1_AOI21X1_12 ( );
FILL FILL_0_NOR2X1_81 ( );
FILL FILL_0_NAND2X1_315 ( );
FILL FILL_0_NOR2X1_77 ( );
FILL FILL_0_NAND2X1_290 ( );
FILL FILL_1_NAND2X1_290 ( );
FILL FILL_0_NAND2X1_291 ( );
FILL FILL_1_NAND2X1_291 ( );
FILL FILL_0_NOR3X1_5 ( );
FILL FILL_1_NOR3X1_5 ( );
FILL FILL_2_NOR3X1_5 ( );
FILL FILL_3_NOR3X1_5 ( );
FILL FILL_0_OAI21X1_603 ( );
FILL FILL_1_OAI21X1_603 ( );
FILL FILL_0_NAND2X1_209 ( );
FILL FILL_1_NAND2X1_209 ( );
FILL FILL_0_DFFPOSX1_601 ( );
FILL FILL_1_DFFPOSX1_601 ( );
FILL FILL_2_DFFPOSX1_601 ( );
FILL FILL_3_DFFPOSX1_601 ( );
FILL FILL_4_DFFPOSX1_601 ( );
FILL FILL_5_DFFPOSX1_601 ( );
FILL FILL_6_DFFPOSX1_601 ( );
FILL FILL_0_NOR2X1_79 ( );
FILL FILL_0_OAI21X1_719 ( );
FILL FILL_1_OAI21X1_719 ( );
FILL FILL_0_OAI21X1_720 ( );
FILL FILL_1_OAI21X1_720 ( );
FILL FILL_2_OAI21X1_720 ( );
FILL FILL_0_OAI21X1_721 ( );
FILL FILL_1_OAI21X1_721 ( );
FILL FILL_0_NAND2X1_171 ( );
FILL FILL_0_XNOR2X1_35 ( );
FILL FILL_1_XNOR2X1_35 ( );
FILL FILL_2_XNOR2X1_35 ( );
FILL FILL_3_XNOR2X1_35 ( );
FILL FILL_0_NAND2X1_175 ( );
FILL FILL_1_NAND2X1_175 ( );
FILL FILL_0_NAND2X1_168 ( );
FILL FILL_1_NAND2X1_168 ( );
FILL FILL_0_XNOR2X1_44 ( );
FILL FILL_1_XNOR2X1_44 ( );
FILL FILL_2_XNOR2X1_44 ( );
FILL FILL_3_XNOR2X1_44 ( );
FILL FILL_0_OAI21X1_550 ( );
FILL FILL_1_OAI21X1_550 ( );
FILL FILL_0_OAI21X1_557 ( );
FILL FILL_1_OAI21X1_557 ( );
FILL FILL_0_BUFX2_606 ( );
FILL FILL_1_BUFX2_606 ( );
FILL FILL_0_NOR2X1_69 ( );
FILL FILL_1_NOR2X1_69 ( );
FILL FILL_0_NAND2X1_319 ( );
FILL FILL_0_NAND2X1_187 ( );
FILL FILL_1_NAND2X1_187 ( );
FILL FILL_0_OAI21X1_575 ( );
FILL FILL_1_OAI21X1_575 ( );
FILL FILL_0_XNOR2X1_46 ( );
FILL FILL_1_XNOR2X1_46 ( );
FILL FILL_2_XNOR2X1_46 ( );
FILL FILL_3_XNOR2X1_46 ( );
FILL FILL_0_OAI21X1_739 ( );
FILL FILL_1_OAI21X1_739 ( );
FILL FILL_0_NAND2X1_321 ( );
FILL FILL_0_INVX1_11 ( );
FILL FILL_0_NAND3X1_2 ( );
FILL FILL_1_NAND3X1_2 ( );
FILL FILL_2_NAND3X1_2 ( );
FILL FILL_0_NAND2X1_323 ( );
FILL FILL_1_NAND2X1_323 ( );
FILL FILL_0_NAND2X1_322 ( );
FILL FILL_0_NOR2X1_108 ( );
FILL FILL_1_NOR2X1_108 ( );
FILL FILL_0_OAI21X1_730 ( );
FILL FILL_1_OAI21X1_730 ( );
FILL FILL_0_NAND2X1_192 ( );
FILL FILL_1_NAND2X1_192 ( );
FILL FILL_0_INVX4_11 ( );
FILL FILL_0_OAI21X1_729 ( );
FILL FILL_1_OAI21X1_729 ( );
FILL FILL_0_OAI21X1_728 ( );
FILL FILL_1_OAI21X1_728 ( );
FILL FILL_0_XNOR2X1_47 ( );
FILL FILL_1_XNOR2X1_47 ( );
FILL FILL_2_XNOR2X1_47 ( );
FILL FILL_3_XNOR2X1_47 ( );
FILL FILL_0_OAI21X1_743 ( );
FILL FILL_1_OAI21X1_743 ( );
FILL FILL_0_OAI21X1_742 ( );
FILL FILL_1_OAI21X1_742 ( );
FILL FILL_0_DFFPOSX1_577 ( );
FILL FILL_1_DFFPOSX1_577 ( );
FILL FILL_2_DFFPOSX1_577 ( );
FILL FILL_3_DFFPOSX1_577 ( );
FILL FILL_4_DFFPOSX1_577 ( );
FILL FILL_5_DFFPOSX1_577 ( );
FILL FILL_6_DFFPOSX1_577 ( );
FILL FILL_0_BUFX2_1025 ( );
FILL FILL_1_BUFX2_1025 ( );
FILL FILL_0_BUFX2_603 ( );
FILL FILL_1_BUFX2_603 ( );
FILL FILL_0_DFFPOSX1_956 ( );
FILL FILL_1_DFFPOSX1_956 ( );
FILL FILL_2_DFFPOSX1_956 ( );
FILL FILL_3_DFFPOSX1_956 ( );
FILL FILL_4_DFFPOSX1_956 ( );
FILL FILL_5_DFFPOSX1_956 ( );
FILL FILL_6_DFFPOSX1_956 ( );
FILL FILL_0_OAI21X1_1264 ( );
FILL FILL_1_OAI21X1_1264 ( );
FILL FILL_0_BUFX2_1026 ( );
FILL FILL_0_NAND2X1_502 ( );
FILL FILL_0_NAND2X1_512 ( );
FILL FILL_0_NAND2X1_509 ( );
FILL FILL_0_OR2X2_17 ( );
FILL FILL_1_OR2X2_17 ( );
FILL FILL_0_NOR2X1_189 ( );
FILL FILL_0_MUX2X1_2 ( );
FILL FILL_1_MUX2X1_2 ( );
FILL FILL_2_MUX2X1_2 ( );
FILL FILL_0_OAI21X1_1132 ( );
FILL FILL_1_OAI21X1_1132 ( );
FILL FILL_2_OAI21X1_1132 ( );
FILL FILL_0_OAI21X1_1453 ( );
FILL FILL_1_OAI21X1_1453 ( );
FILL FILL_0_OAI21X1_1265 ( );
FILL FILL_1_OAI21X1_1265 ( );
FILL FILL_0_BUFX2_20 ( );
FILL FILL_0_OAI21X1_1267 ( );
FILL FILL_1_OAI21X1_1267 ( );
FILL FILL_0_DFFPOSX1_892 ( );
FILL FILL_1_DFFPOSX1_892 ( );
FILL FILL_2_DFFPOSX1_892 ( );
FILL FILL_3_DFFPOSX1_892 ( );
FILL FILL_4_DFFPOSX1_892 ( );
FILL FILL_5_DFFPOSX1_892 ( );
FILL FILL_0_OAI21X1_1014 ( );
FILL FILL_1_OAI21X1_1014 ( );
FILL FILL_0_DFFPOSX1_845 ( );
FILL FILL_1_DFFPOSX1_845 ( );
FILL FILL_2_DFFPOSX1_845 ( );
FILL FILL_3_DFFPOSX1_845 ( );
FILL FILL_4_DFFPOSX1_845 ( );
FILL FILL_5_DFFPOSX1_845 ( );
FILL FILL_6_DFFPOSX1_845 ( );
FILL FILL_0_OAI21X1_1161 ( );
FILL FILL_1_OAI21X1_1161 ( );
FILL FILL_0_NAND2X1_538 ( );
FILL FILL_1_NAND2X1_538 ( );
FILL FILL_0_NOR2X1_198 ( );
FILL FILL_1_NOR2X1_198 ( );
FILL FILL_0_OAI21X1_1485 ( );
FILL FILL_1_OAI21X1_1485 ( );
FILL FILL_2_OAI21X1_1485 ( );
FILL FILL_0_OAI21X1_1490 ( );
FILL FILL_1_OAI21X1_1490 ( );
FILL FILL_0_NOR2X1_200 ( );
FILL FILL_1_NOR2X1_200 ( );
FILL FILL_0_INVX2_100 ( );
FILL FILL_0_NOR2X1_153 ( );
FILL FILL_1_NOR2X1_153 ( );
FILL FILL_0_AND2X2_31 ( );
FILL FILL_1_AND2X2_31 ( );
FILL FILL_0_OAI21X1_1492 ( );
FILL FILL_1_OAI21X1_1492 ( );
FILL FILL_0_DFFPOSX1_842 ( );
FILL FILL_1_DFFPOSX1_842 ( );
FILL FILL_2_DFFPOSX1_842 ( );
FILL FILL_3_DFFPOSX1_842 ( );
FILL FILL_4_DFFPOSX1_842 ( );
FILL FILL_5_DFFPOSX1_842 ( );
FILL FILL_0_OAI21X1_1491 ( );
FILL FILL_1_OAI21X1_1491 ( );
FILL FILL_0_BUFX2_93 ( );
FILL FILL_1_BUFX2_93 ( );
FILL FILL_0_OAI21X1_1538 ( );
FILL FILL_1_OAI21X1_1538 ( );
FILL FILL_0_OAI21X1_1371 ( );
FILL FILL_1_OAI21X1_1371 ( );
FILL FILL_0_DFFPOSX1_930 ( );
FILL FILL_1_DFFPOSX1_930 ( );
FILL FILL_2_DFFPOSX1_930 ( );
FILL FILL_3_DFFPOSX1_930 ( );
FILL FILL_4_DFFPOSX1_930 ( );
FILL FILL_5_DFFPOSX1_930 ( );
FILL FILL_6_DFFPOSX1_930 ( );
FILL FILL_0_AOI21X1_63 ( );
FILL FILL_1_AOI21X1_63 ( );
FILL FILL_0_BUFX4_66 ( );
FILL FILL_1_BUFX4_66 ( );
FILL FILL_2_BUFX4_66 ( );
FILL FILL_0_NOR2X1_168 ( );
FILL FILL_0_INVX2_85 ( );
FILL FILL_0_BUFX4_242 ( );
FILL FILL_1_BUFX4_242 ( );
FILL FILL_0_NAND3X1_47 ( );
FILL FILL_1_NAND3X1_47 ( );
FILL FILL_0_BUFX4_12 ( );
FILL FILL_1_BUFX4_12 ( );
FILL FILL_0_OAI21X1_1356 ( );
FILL FILL_1_OAI21X1_1356 ( );
FILL FILL_0_NAND2X1_621 ( );
FILL FILL_1_NAND2X1_621 ( );
FILL FILL_0_INVX1_196 ( );
FILL FILL_0_INVX1_214 ( );
FILL FILL_0_NAND2X1_622 ( );
FILL FILL_0_OAI21X1_1194 ( );
FILL FILL_1_OAI21X1_1194 ( );
FILL FILL_0_NAND2X1_580 ( );
FILL FILL_0_AOI21X1_57 ( );
FILL FILL_1_AOI21X1_57 ( );
FILL FILL_0_NAND3X1_68 ( );
FILL FILL_1_NAND3X1_68 ( );
FILL FILL_0_INVX1_215 ( );
FILL FILL_0_NOR2X1_209 ( );
FILL FILL_1_NOR2X1_209 ( );
FILL FILL_0_OAI21X1_1359 ( );
FILL FILL_1_OAI21X1_1359 ( );
FILL FILL_0_AOI21X1_55 ( );
FILL FILL_1_AOI21X1_55 ( );
FILL FILL_0_OAI21X1_1360 ( );
FILL FILL_1_OAI21X1_1360 ( );
FILL FILL_0_OAI21X1_1358 ( );
FILL FILL_1_OAI21X1_1358 ( );
FILL FILL_2_OAI21X1_1358 ( );
FILL FILL_0_DFFPOSX1_927 ( );
FILL FILL_1_DFFPOSX1_927 ( );
FILL FILL_2_DFFPOSX1_927 ( );
FILL FILL_3_DFFPOSX1_927 ( );
FILL FILL_4_DFFPOSX1_927 ( );
FILL FILL_5_DFFPOSX1_927 ( );
FILL FILL_0_BUFX2_182 ( );
FILL FILL_1_BUFX2_182 ( );
FILL FILL_0_CLKBUF1_69 ( );
FILL FILL_1_CLKBUF1_69 ( );
FILL FILL_2_CLKBUF1_69 ( );
FILL FILL_3_CLKBUF1_69 ( );
FILL FILL_0_OAI21X1_302 ( );
FILL FILL_1_OAI21X1_302 ( );
FILL FILL_0_OAI21X1_303 ( );
FILL FILL_1_OAI21X1_303 ( );
FILL FILL_0_DFFPOSX1_343 ( );
FILL FILL_1_DFFPOSX1_343 ( );
FILL FILL_2_DFFPOSX1_343 ( );
FILL FILL_3_DFFPOSX1_343 ( );
FILL FILL_4_DFFPOSX1_343 ( );
FILL FILL_5_DFFPOSX1_343 ( );
FILL FILL_6_DFFPOSX1_343 ( );
FILL FILL_0_BUFX2_965 ( );
FILL FILL_1_BUFX2_965 ( );
FILL FILL_0_OAI21X1_940 ( );
FILL FILL_1_OAI21X1_940 ( );
FILL FILL_0_OAI21X1_941 ( );
FILL FILL_1_OAI21X1_941 ( );
FILL FILL_0_DFFPOSX1_696 ( );
FILL FILL_1_DFFPOSX1_696 ( );
FILL FILL_2_DFFPOSX1_696 ( );
FILL FILL_3_DFFPOSX1_696 ( );
FILL FILL_4_DFFPOSX1_696 ( );
FILL FILL_5_DFFPOSX1_696 ( );
FILL FILL_6_DFFPOSX1_696 ( );
FILL FILL_0_OAI21X1_1002 ( );
FILL FILL_1_OAI21X1_1002 ( );
FILL FILL_0_BUFX2_177 ( );
FILL FILL_1_BUFX2_177 ( );
FILL FILL_0_BUFX2_1016 ( );
FILL FILL_1_BUFX2_1016 ( );
FILL FILL_0_INVX1_77 ( );
FILL FILL_1_INVX1_77 ( );
FILL FILL_0_BUFX2_675 ( );
FILL FILL_0_DFFPOSX1_290 ( );
FILL FILL_1_DFFPOSX1_290 ( );
FILL FILL_2_DFFPOSX1_290 ( );
FILL FILL_3_DFFPOSX1_290 ( );
FILL FILL_4_DFFPOSX1_290 ( );
FILL FILL_5_DFFPOSX1_290 ( );
FILL FILL_0_OAI21X1_196 ( );
FILL FILL_1_OAI21X1_196 ( );
FILL FILL_0_OAI21X1_197 ( );
FILL FILL_1_OAI21X1_197 ( );
FILL FILL_0_DFFPOSX1_274 ( );
FILL FILL_1_DFFPOSX1_274 ( );
FILL FILL_2_DFFPOSX1_274 ( );
FILL FILL_3_DFFPOSX1_274 ( );
FILL FILL_4_DFFPOSX1_274 ( );
FILL FILL_5_DFFPOSX1_274 ( );
FILL FILL_0_OAI21X1_165 ( );
FILL FILL_1_OAI21X1_165 ( );
FILL FILL_0_OAI21X1_164 ( );
FILL FILL_1_OAI21X1_164 ( );
FILL FILL_0_BUFX2_405 ( );
FILL FILL_1_BUFX2_405 ( );
FILL FILL_0_BUFX2_928 ( );
FILL FILL_1_BUFX2_928 ( );
FILL FILL_0_BUFX4_134 ( );
FILL FILL_1_BUFX4_134 ( );
FILL FILL_0_DFFPOSX1_423 ( );
FILL FILL_1_DFFPOSX1_423 ( );
FILL FILL_2_DFFPOSX1_423 ( );
FILL FILL_3_DFFPOSX1_423 ( );
FILL FILL_4_DFFPOSX1_423 ( );
FILL FILL_5_DFFPOSX1_423 ( );
FILL FILL_6_DFFPOSX1_423 ( );
FILL FILL_0_NAND2X1_137 ( );
FILL FILL_1_NAND2X1_137 ( );
FILL FILL_0_OAI21X1_398 ( );
FILL FILL_1_OAI21X1_398 ( );
FILL FILL_2_OAI21X1_398 ( );
FILL FILL_0_DFFPOSX1_485 ( );
FILL FILL_1_DFFPOSX1_485 ( );
FILL FILL_2_DFFPOSX1_485 ( );
FILL FILL_3_DFFPOSX1_485 ( );
FILL FILL_4_DFFPOSX1_485 ( );
FILL FILL_5_DFFPOSX1_485 ( );
FILL FILL_0_OAI21X1_503 ( );
FILL FILL_1_OAI21X1_503 ( );
FILL FILL_0_OAI21X1_502 ( );
FILL FILL_1_OAI21X1_502 ( );
FILL FILL_0_NOR2X1_1 ( );
FILL FILL_1_NOR2X1_1 ( );
FILL FILL_0_NOR2X1_3 ( );
FILL FILL_1_NOR2X1_3 ( );
FILL FILL_0_DFFPOSX1_498 ( );
FILL FILL_1_DFFPOSX1_498 ( );
FILL FILL_2_DFFPOSX1_498 ( );
FILL FILL_3_DFFPOSX1_498 ( );
FILL FILL_4_DFFPOSX1_498 ( );
FILL FILL_5_DFFPOSX1_498 ( );
FILL FILL_0_OAI21X1_541 ( );
FILL FILL_1_OAI21X1_541 ( );
FILL FILL_0_INVX1_7 ( );
FILL FILL_0_NOR2X1_2 ( );
FILL FILL_0_DFFPOSX1_501 ( );
FILL FILL_1_DFFPOSX1_501 ( );
FILL FILL_2_DFFPOSX1_501 ( );
FILL FILL_3_DFFPOSX1_501 ( );
FILL FILL_4_DFFPOSX1_501 ( );
FILL FILL_5_DFFPOSX1_501 ( );
FILL FILL_6_DFFPOSX1_501 ( );
FILL FILL_0_DFFPOSX1_402 ( );
FILL FILL_1_DFFPOSX1_402 ( );
FILL FILL_2_DFFPOSX1_402 ( );
FILL FILL_3_DFFPOSX1_402 ( );
FILL FILL_4_DFFPOSX1_402 ( );
FILL FILL_5_DFFPOSX1_402 ( );
FILL FILL_0_BUFX4_372 ( );
FILL FILL_1_BUFX4_372 ( );
FILL FILL_0_OAI21X1_374 ( );
FILL FILL_1_OAI21X1_374 ( );
FILL FILL_0_DFFPOSX1_560 ( );
FILL FILL_1_DFFPOSX1_560 ( );
FILL FILL_2_DFFPOSX1_560 ( );
FILL FILL_3_DFFPOSX1_560 ( );
FILL FILL_4_DFFPOSX1_560 ( );
FILL FILL_5_DFFPOSX1_560 ( );
FILL FILL_0_DFFPOSX1_519 ( );
FILL FILL_1_DFFPOSX1_519 ( );
FILL FILL_2_DFFPOSX1_519 ( );
FILL FILL_3_DFFPOSX1_519 ( );
FILL FILL_4_DFFPOSX1_519 ( );
FILL FILL_5_DFFPOSX1_519 ( );
FILL FILL_0_INVX2_31 ( );
FILL FILL_0_OAI21X1_618 ( );
FILL FILL_1_OAI21X1_618 ( );
FILL FILL_0_OAI21X1_594 ( );
FILL FILL_1_OAI21X1_594 ( );
FILL FILL_0_DFFPOSX1_530 ( );
FILL FILL_1_DFFPOSX1_530 ( );
FILL FILL_2_DFFPOSX1_530 ( );
FILL FILL_3_DFFPOSX1_530 ( );
FILL FILL_4_DFFPOSX1_530 ( );
FILL FILL_5_DFFPOSX1_530 ( );
FILL FILL_0_OAI21X1_620 ( );
FILL FILL_1_OAI21X1_620 ( );
FILL FILL_0_AOI21X1_15 ( );
FILL FILL_1_AOI21X1_15 ( );
FILL FILL_2_AOI21X1_15 ( );
FILL FILL_0_NOR2X1_39 ( );
FILL FILL_1_NOR2X1_39 ( );
FILL FILL_0_INVX2_30 ( );
FILL FILL_0_XNOR2X1_28 ( );
FILL FILL_1_XNOR2X1_28 ( );
FILL FILL_2_XNOR2X1_28 ( );
FILL FILL_0_NAND3X1_9 ( );
FILL FILL_1_NAND3X1_9 ( );
FILL FILL_0_BUFX4_114 ( );
FILL FILL_1_BUFX4_114 ( );
FILL FILL_0_DFFPOSX1_532 ( );
FILL FILL_1_DFFPOSX1_532 ( );
FILL FILL_2_DFFPOSX1_532 ( );
FILL FILL_3_DFFPOSX1_532 ( );
FILL FILL_4_DFFPOSX1_532 ( );
FILL FILL_5_DFFPOSX1_532 ( );
FILL FILL_0_NOR2X1_50 ( );
FILL FILL_0_AND2X2_10 ( );
FILL FILL_1_AND2X2_10 ( );
FILL FILL_0_OAI21X1_479 ( );
FILL FILL_1_OAI21X1_479 ( );
FILL FILL_0_OAI21X1_482 ( );
FILL FILL_1_OAI21X1_482 ( );
FILL FILL_2_OAI21X1_482 ( );
FILL FILL_0_DFFPOSX1_602 ( );
FILL FILL_1_DFFPOSX1_602 ( );
FILL FILL_2_DFFPOSX1_602 ( );
FILL FILL_3_DFFPOSX1_602 ( );
FILL FILL_4_DFFPOSX1_602 ( );
FILL FILL_5_DFFPOSX1_602 ( );
FILL FILL_0_BUFX4_240 ( );
FILL FILL_1_BUFX4_240 ( );
FILL FILL_0_DFFPOSX1_388 ( );
FILL FILL_1_DFFPOSX1_388 ( );
FILL FILL_2_DFFPOSX1_388 ( );
FILL FILL_3_DFFPOSX1_388 ( );
FILL FILL_4_DFFPOSX1_388 ( );
FILL FILL_5_DFFPOSX1_388 ( );
FILL FILL_6_DFFPOSX1_388 ( );
FILL FILL_0_NAND2X1_104 ( );
FILL FILL_0_OAI21X1_360 ( );
FILL FILL_1_OAI21X1_360 ( );
FILL FILL_0_OAI21X1_592 ( );
FILL FILL_1_OAI21X1_592 ( );
FILL FILL_0_OAI21X1_591 ( );
FILL FILL_1_OAI21X1_591 ( );
FILL FILL_0_OR2X2_8 ( );
FILL FILL_1_OR2X2_8 ( );
FILL FILL_2_OR2X2_8 ( );
FILL FILL_0_NOR2X1_110 ( );
FILL FILL_1_NOR2X1_110 ( );
FILL FILL_0_BUFX4_74 ( );
FILL FILL_1_BUFX4_74 ( );
FILL FILL_0_NOR2X1_31 ( );
FILL FILL_0_OAI21X1_788 ( );
FILL FILL_1_OAI21X1_788 ( );
FILL FILL_0_NOR2X1_75 ( );
FILL FILL_1_NOR2X1_75 ( );
FILL FILL_0_OAI21X1_815 ( );
FILL FILL_1_OAI21X1_815 ( );
FILL FILL_0_OAI21X1_814 ( );
FILL FILL_1_OAI21X1_814 ( );
FILL FILL_0_DFFPOSX1_570 ( );
FILL FILL_1_DFFPOSX1_570 ( );
FILL FILL_2_DFFPOSX1_570 ( );
FILL FILL_3_DFFPOSX1_570 ( );
FILL FILL_4_DFFPOSX1_570 ( );
FILL FILL_5_DFFPOSX1_570 ( );
FILL FILL_6_DFFPOSX1_570 ( );
FILL FILL_0_OAI21X1_724 ( );
FILL FILL_1_OAI21X1_724 ( );
FILL FILL_0_INVX2_26 ( );
FILL FILL_1_INVX2_26 ( );
FILL FILL_0_OAI21X1_426 ( );
FILL FILL_1_OAI21X1_426 ( );
FILL FILL_0_NAND2X1_172 ( );
FILL FILL_1_NAND2X1_172 ( );
FILL FILL_0_INVX2_19 ( );
FILL FILL_0_OAI21X1_722 ( );
FILL FILL_1_OAI21X1_722 ( );
FILL FILL_0_OAI21X1_549 ( );
FILL FILL_1_OAI21X1_549 ( );
FILL FILL_0_NAND2X1_202 ( );
FILL FILL_1_NAND2X1_202 ( );
FILL FILL_0_OAI21X1_428 ( );
FILL FILL_1_OAI21X1_428 ( );
FILL FILL_0_NAND2X1_178 ( );
FILL FILL_1_NAND2X1_178 ( );
FILL FILL_0_OR2X2_2 ( );
FILL FILL_1_OR2X2_2 ( );
FILL FILL_0_BUFX4_245 ( );
FILL FILL_1_BUFX4_245 ( );
FILL FILL_0_NOR2X1_109 ( );
FILL FILL_0_OAI21X1_727 ( );
FILL FILL_1_OAI21X1_727 ( );
FILL FILL_0_OAI21X1_741 ( );
FILL FILL_1_OAI21X1_741 ( );
FILL FILL_0_NOR2X1_22 ( );
FILL FILL_1_NOR2X1_22 ( );
FILL FILL_0_OR2X2_4 ( );
FILL FILL_1_OR2X2_4 ( );
FILL FILL_0_NOR2X1_28 ( );
FILL FILL_1_NOR2X1_28 ( );
FILL FILL_0_NOR3X1_1 ( );
FILL FILL_1_NOR3X1_1 ( );
FILL FILL_2_NOR3X1_1 ( );
FILL FILL_3_NOR3X1_1 ( );
FILL FILL_4_NOR3X1_1 ( );
FILL FILL_0_BUFX2_543 ( );
FILL FILL_1_BUFX2_543 ( );
FILL FILL_0_OAI21X1_438 ( );
FILL FILL_1_OAI21X1_438 ( );
FILL FILL_0_INVX2_22 ( );
FILL FILL_0_INVX1_12 ( );
FILL FILL_0_NOR2X1_18 ( );
FILL FILL_0_AOI21X1_32 ( );
FILL FILL_1_AOI21X1_32 ( );
FILL FILL_0_NAND2X1_320 ( );
FILL FILL_1_NAND2X1_320 ( );
FILL FILL_0_INVX1_38 ( );
FILL FILL_0_DFFPOSX1_572 ( );
FILL FILL_1_DFFPOSX1_572 ( );
FILL FILL_2_DFFPOSX1_572 ( );
FILL FILL_3_DFFPOSX1_572 ( );
FILL FILL_4_DFFPOSX1_572 ( );
FILL FILL_5_DFFPOSX1_572 ( );
FILL FILL_6_DFFPOSX1_572 ( );
FILL FILL_0_BUFX2_636 ( );
FILL FILL_0_DFFPOSX1_352 ( );
FILL FILL_1_DFFPOSX1_352 ( );
FILL FILL_2_DFFPOSX1_352 ( );
FILL FILL_3_DFFPOSX1_352 ( );
FILL FILL_4_DFFPOSX1_352 ( );
FILL FILL_5_DFFPOSX1_352 ( );
FILL FILL_0_OAI21X1_321 ( );
FILL FILL_1_OAI21X1_321 ( );
FILL FILL_0_DFFPOSX1_894 ( );
FILL FILL_1_DFFPOSX1_894 ( );
FILL FILL_2_DFFPOSX1_894 ( );
FILL FILL_3_DFFPOSX1_894 ( );
FILL FILL_4_DFFPOSX1_894 ( );
FILL FILL_5_DFFPOSX1_894 ( );
FILL FILL_0_OAI21X1_1273 ( );
FILL FILL_1_OAI21X1_1273 ( );
FILL FILL_0_OAI21X1_1274 ( );
FILL FILL_1_OAI21X1_1274 ( );
FILL FILL_0_OAI21X1_1272 ( );
FILL FILL_1_OAI21X1_1272 ( );
FILL FILL_0_CLKBUF1_34 ( );
FILL FILL_1_CLKBUF1_34 ( );
FILL FILL_2_CLKBUF1_34 ( );
FILL FILL_3_CLKBUF1_34 ( );
FILL FILL_4_CLKBUF1_34 ( );
FILL FILL_0_NOR2X1_188 ( );
FILL FILL_1_NOR2X1_188 ( );
FILL FILL_0_NOR2X1_187 ( );
FILL FILL_1_NOR2X1_187 ( );
FILL FILL_0_NAND2X1_599 ( );
FILL FILL_1_NAND2X1_599 ( );
FILL FILL_0_NOR2X1_140 ( );
FILL FILL_1_NOR2X1_140 ( );
FILL FILL_0_OR2X2_18 ( );
FILL FILL_1_OR2X2_18 ( );
FILL FILL_0_OAI21X1_1268 ( );
FILL FILL_1_OAI21X1_1268 ( );
FILL FILL_0_XNOR2X1_95 ( );
FILL FILL_1_XNOR2X1_95 ( );
FILL FILL_2_XNOR2X1_95 ( );
FILL FILL_3_XNOR2X1_95 ( );
FILL FILL_0_DFFPOSX1_958 ( );
FILL FILL_1_DFFPOSX1_958 ( );
FILL FILL_2_DFFPOSX1_958 ( );
FILL FILL_3_DFFPOSX1_958 ( );
FILL FILL_4_DFFPOSX1_958 ( );
FILL FILL_5_DFFPOSX1_958 ( );
FILL FILL_6_DFFPOSX1_958 ( );
FILL FILL_0_BUFX4_120 ( );
FILL FILL_1_BUFX4_120 ( );
FILL FILL_0_BUFX4_80 ( );
FILL FILL_1_BUFX4_80 ( );
FILL FILL_0_BUFX4_280 ( );
FILL FILL_1_BUFX4_280 ( );
FILL FILL_2_BUFX4_280 ( );
FILL FILL_0_DFFPOSX1_909 ( );
FILL FILL_1_DFFPOSX1_909 ( );
FILL FILL_2_DFFPOSX1_909 ( );
FILL FILL_3_DFFPOSX1_909 ( );
FILL FILL_4_DFFPOSX1_909 ( );
FILL FILL_5_DFFPOSX1_909 ( );
FILL FILL_0_OAI21X1_1311 ( );
FILL FILL_1_OAI21X1_1311 ( );
FILL FILL_0_XNOR2X1_83 ( );
FILL FILL_1_XNOR2X1_83 ( );
FILL FILL_2_XNOR2X1_83 ( );
FILL FILL_3_XNOR2X1_83 ( );
FILL FILL_0_BUFX2_979 ( );
FILL FILL_0_INVX8_1 ( );
FILL FILL_1_INVX8_1 ( );
FILL FILL_0_OAI21X1_1494 ( );
FILL FILL_1_OAI21X1_1494 ( );
FILL FILL_2_OAI21X1_1494 ( );
FILL FILL_0_OAI21X1_1493 ( );
FILL FILL_1_OAI21X1_1493 ( );
FILL FILL_0_NAND2X1_637 ( );
FILL FILL_1_NAND2X1_637 ( );
FILL FILL_0_NAND2X1_608 ( );
FILL FILL_1_NAND2X1_608 ( );
FILL FILL_0_INVX1_208 ( );
FILL FILL_0_NAND2X1_610 ( );
FILL FILL_0_OAI21X1_1158 ( );
FILL FILL_1_OAI21X1_1158 ( );
FILL FILL_0_NAND2X1_534 ( );
FILL FILL_1_NAND2X1_534 ( );
FILL FILL_0_DFFPOSX1_972 ( );
FILL FILL_1_DFFPOSX1_972 ( );
FILL FILL_2_DFFPOSX1_972 ( );
FILL FILL_3_DFFPOSX1_972 ( );
FILL FILL_4_DFFPOSX1_972 ( );
FILL FILL_5_DFFPOSX1_972 ( );
FILL FILL_0_BUFX4_276 ( );
FILL FILL_1_BUFX4_276 ( );
FILL FILL_0_DFFPOSX1_988 ( );
FILL FILL_1_DFFPOSX1_988 ( );
FILL FILL_2_DFFPOSX1_988 ( );
FILL FILL_3_DFFPOSX1_988 ( );
FILL FILL_4_DFFPOSX1_988 ( );
FILL FILL_5_DFFPOSX1_988 ( );
FILL FILL_6_DFFPOSX1_988 ( );
FILL FILL_0_OAI21X1_1542 ( );
FILL FILL_1_OAI21X1_1542 ( );
FILL FILL_0_OAI21X1_1541 ( );
FILL FILL_1_OAI21X1_1541 ( );
FILL FILL_0_BUFX4_39 ( );
FILL FILL_1_BUFX4_39 ( );
FILL FILL_0_NOR2X1_228 ( );
FILL FILL_1_NOR2X1_228 ( );
FILL FILL_0_NOR3X1_12 ( );
FILL FILL_1_NOR3X1_12 ( );
FILL FILL_2_NOR3X1_12 ( );
FILL FILL_3_NOR3X1_12 ( );
FILL FILL_0_NAND2X1_574 ( );
FILL FILL_0_INVX2_103 ( );
FILL FILL_1_INVX2_103 ( );
FILL FILL_0_OAI21X1_1351 ( );
FILL FILL_1_OAI21X1_1351 ( );
FILL FILL_0_NOR2X1_208 ( );
FILL FILL_0_XNOR2X1_87 ( );
FILL FILL_1_XNOR2X1_87 ( );
FILL FILL_2_XNOR2X1_87 ( );
FILL FILL_3_XNOR2X1_87 ( );
FILL FILL_0_NAND3X1_60 ( );
FILL FILL_1_NAND3X1_60 ( );
FILL FILL_2_NAND3X1_60 ( );
FILL FILL_0_NAND3X1_49 ( );
FILL FILL_1_NAND3X1_49 ( );
FILL FILL_0_INVX1_197 ( );
FILL FILL_0_OAI21X1_1366 ( );
FILL FILL_1_OAI21X1_1366 ( );
FILL FILL_0_OAI21X1_1367 ( );
FILL FILL_1_OAI21X1_1367 ( );
FILL FILL_0_DFFPOSX1_929 ( );
FILL FILL_1_DFFPOSX1_929 ( );
FILL FILL_2_DFFPOSX1_929 ( );
FILL FILL_3_DFFPOSX1_929 ( );
FILL FILL_4_DFFPOSX1_929 ( );
FILL FILL_5_DFFPOSX1_929 ( );
FILL FILL_0_OAI21X1_1365 ( );
FILL FILL_1_OAI21X1_1365 ( );
FILL FILL_0_BUFX4_277 ( );
FILL FILL_1_BUFX4_277 ( );
FILL FILL_0_BUFX4_58 ( );
FILL FILL_1_BUFX4_58 ( );
FILL FILL_0_OAI21X1_1352 ( );
FILL FILL_1_OAI21X1_1352 ( );
FILL FILL_0_DFFPOSX1_924 ( );
FILL FILL_1_DFFPOSX1_924 ( );
FILL FILL_2_DFFPOSX1_924 ( );
FILL FILL_3_DFFPOSX1_924 ( );
FILL FILL_4_DFFPOSX1_924 ( );
FILL FILL_5_DFFPOSX1_924 ( );
FILL FILL_0_OAI21X1_1350 ( );
FILL FILL_1_OAI21X1_1350 ( );
FILL FILL_0_BUFX2_229 ( );
FILL FILL_1_BUFX2_229 ( );
FILL FILL_0_OAI21X1_198 ( );
FILL FILL_1_OAI21X1_198 ( );
FILL FILL_0_OAI21X1_199 ( );
FILL FILL_1_OAI21X1_199 ( );
FILL FILL_0_DFFPOSX1_291 ( );
FILL FILL_1_DFFPOSX1_291 ( );
FILL FILL_2_DFFPOSX1_291 ( );
FILL FILL_3_DFFPOSX1_291 ( );
FILL FILL_4_DFFPOSX1_291 ( );
FILL FILL_5_DFFPOSX1_291 ( );
FILL FILL_6_DFFPOSX1_291 ( );
FILL FILL_0_CLKBUF1_40 ( );
FILL FILL_1_CLKBUF1_40 ( );
FILL FILL_2_CLKBUF1_40 ( );
FILL FILL_3_CLKBUF1_40 ( );
FILL FILL_4_CLKBUF1_40 ( );
FILL FILL_0_OAI21X1_1704 ( );
FILL FILL_1_OAI21X1_1704 ( );
FILL FILL_0_OAI21X1_1705 ( );
FILL FILL_1_OAI21X1_1705 ( );
FILL FILL_2_OAI21X1_1705 ( );
FILL FILL_0_OAI21X1_1750 ( );
FILL FILL_1_OAI21X1_1750 ( );
FILL FILL_0_INVX2_185 ( );
FILL FILL_0_OAI21X1_953 ( );
FILL FILL_1_OAI21X1_953 ( );
FILL FILL_0_DFFPOSX1_702 ( );
FILL FILL_1_DFFPOSX1_702 ( );
FILL FILL_2_DFFPOSX1_702 ( );
FILL FILL_3_DFFPOSX1_702 ( );
FILL FILL_4_DFFPOSX1_702 ( );
FILL FILL_5_DFFPOSX1_702 ( );
FILL FILL_6_DFFPOSX1_702 ( );
FILL FILL_0_BUFX2_293 ( );
FILL FILL_0_BUFX2_1020 ( );
FILL FILL_1_BUFX2_1020 ( );
FILL FILL_0_OAI21X1_876 ( );
FILL FILL_1_OAI21X1_876 ( );
FILL FILL_0_NAND2X1_370 ( );
FILL FILL_0_NAND2X1_654 ( );
FILL FILL_0_DFFPOSX1_648 ( );
FILL FILL_1_DFFPOSX1_648 ( );
FILL FILL_2_DFFPOSX1_648 ( );
FILL FILL_3_DFFPOSX1_648 ( );
FILL FILL_4_DFFPOSX1_648 ( );
FILL FILL_5_DFFPOSX1_648 ( );
FILL FILL_6_DFFPOSX1_648 ( );
FILL FILL_0_BUFX2_416 ( );
FILL FILL_1_BUFX2_416 ( );
FILL FILL_0_BUFX2_469 ( );
FILL FILL_0_BUFX4_102 ( );
FILL FILL_1_BUFX4_102 ( );
FILL FILL_0_BUFX2_565 ( );
FILL FILL_1_BUFX2_565 ( );
FILL FILL_0_DFFPOSX1_359 ( );
FILL FILL_1_DFFPOSX1_359 ( );
FILL FILL_2_DFFPOSX1_359 ( );
FILL FILL_3_DFFPOSX1_359 ( );
FILL FILL_4_DFFPOSX1_359 ( );
FILL FILL_5_DFFPOSX1_359 ( );
FILL FILL_0_NAND2X1_75 ( );
FILL FILL_1_NAND2X1_75 ( );
FILL FILL_0_OAI21X1_331 ( );
FILL FILL_1_OAI21X1_331 ( );
FILL FILL_0_BUFX2_533 ( );
FILL FILL_1_BUFX2_533 ( );
FILL FILL_0_BUFX2_588 ( );
FILL FILL_1_BUFX2_588 ( );
FILL FILL_0_NAND2X1_139 ( );
FILL FILL_1_NAND2X1_139 ( );
FILL FILL_0_OAI21X1_397 ( );
FILL FILL_1_OAI21X1_397 ( );
FILL FILL_0_OAI21X1_662 ( );
FILL FILL_1_OAI21X1_662 ( );
FILL FILL_2_OAI21X1_662 ( );
FILL FILL_0_INVX2_9 ( );
FILL FILL_0_INVX2_8 ( );
FILL FILL_0_AOI21X1_29 ( );
FILL FILL_1_AOI21X1_29 ( );
FILL FILL_0_NAND2X1_266 ( );
FILL FILL_1_NAND2X1_266 ( );
FILL FILL_0_OAI21X1_663 ( );
FILL FILL_1_OAI21X1_663 ( );
FILL FILL_0_OAI21X1_540 ( );
FILL FILL_1_OAI21X1_540 ( );
FILL FILL_0_OAI21X1_667 ( );
FILL FILL_1_OAI21X1_667 ( );
FILL FILL_0_OAI21X1_666 ( );
FILL FILL_1_OAI21X1_666 ( );
FILL FILL_0_OAI21X1_330 ( );
FILL FILL_1_OAI21X1_330 ( );
FILL FILL_0_BUFX4_365 ( );
FILL FILL_1_BUFX4_365 ( );
FILL FILL_0_BUFX2_428 ( );
FILL FILL_0_DFFPOSX1_396 ( );
FILL FILL_1_DFFPOSX1_396 ( );
FILL FILL_2_DFFPOSX1_396 ( );
FILL FILL_3_DFFPOSX1_396 ( );
FILL FILL_4_DFFPOSX1_396 ( );
FILL FILL_5_DFFPOSX1_396 ( );
FILL FILL_0_OAI21X1_368 ( );
FILL FILL_1_OAI21X1_368 ( );
FILL FILL_0_BUFX4_358 ( );
FILL FILL_1_BUFX4_358 ( );
FILL FILL_0_DFFPOSX1_408 ( );
FILL FILL_1_DFFPOSX1_408 ( );
FILL FILL_2_DFFPOSX1_408 ( );
FILL FILL_3_DFFPOSX1_408 ( );
FILL FILL_4_DFFPOSX1_408 ( );
FILL FILL_5_DFFPOSX1_408 ( );
FILL FILL_6_DFFPOSX1_408 ( );
FILL FILL_0_NAND2X1_124 ( );
FILL FILL_1_NAND2X1_124 ( );
FILL FILL_0_OAI21X1_380 ( );
FILL FILL_1_OAI21X1_380 ( );
FILL FILL_0_DFFPOSX1_400 ( );
FILL FILL_1_DFFPOSX1_400 ( );
FILL FILL_2_DFFPOSX1_400 ( );
FILL FILL_3_DFFPOSX1_400 ( );
FILL FILL_4_DFFPOSX1_400 ( );
FILL FILL_5_DFFPOSX1_400 ( );
FILL FILL_0_OAI21X1_790 ( );
FILL FILL_1_OAI21X1_790 ( );
FILL FILL_0_DFFPOSX1_594 ( );
FILL FILL_1_DFFPOSX1_594 ( );
FILL FILL_2_DFFPOSX1_594 ( );
FILL FILL_3_DFFPOSX1_594 ( );
FILL FILL_4_DFFPOSX1_594 ( );
FILL FILL_5_DFFPOSX1_594 ( );
FILL FILL_6_DFFPOSX1_594 ( );
FILL FILL_0_OAI21X1_792 ( );
FILL FILL_1_OAI21X1_792 ( );
FILL FILL_2_OAI21X1_792 ( );
FILL FILL_0_AND2X2_22 ( );
FILL FILL_1_AND2X2_22 ( );
FILL FILL_2_AND2X2_22 ( );
FILL FILL_0_OAI21X1_621 ( );
FILL FILL_1_OAI21X1_621 ( );
FILL FILL_0_OAI21X1_791 ( );
FILL FILL_1_OAI21X1_791 ( );
FILL FILL_0_OAI21X1_623 ( );
FILL FILL_1_OAI21X1_623 ( );
FILL FILL_2_OAI21X1_623 ( );
FILL FILL_0_AND2X2_13 ( );
FILL FILL_1_AND2X2_13 ( );
FILL FILL_0_AOI21X1_16 ( );
FILL FILL_1_AOI21X1_16 ( );
FILL FILL_0_OAI21X1_787 ( );
FILL FILL_1_OAI21X1_787 ( );
FILL FILL_0_NAND2X1_329 ( );
FILL FILL_1_NAND2X1_329 ( );
FILL FILL_0_OAI21X1_622 ( );
FILL FILL_1_OAI21X1_622 ( );
FILL FILL_0_INVX1_18 ( );
FILL FILL_0_NAND2X1_298 ( );
FILL FILL_1_NAND2X1_298 ( );
FILL FILL_0_AOI21X1_18 ( );
FILL FILL_1_AOI21X1_18 ( );
FILL FILL_0_NOR2X1_89 ( );
FILL FILL_0_DFFPOSX1_597 ( );
FILL FILL_1_DFFPOSX1_597 ( );
FILL FILL_2_DFFPOSX1_597 ( );
FILL FILL_3_DFFPOSX1_597 ( );
FILL FILL_4_DFFPOSX1_597 ( );
FILL FILL_5_DFFPOSX1_597 ( );
FILL FILL_0_AOI21X1_34 ( );
FILL FILL_1_AOI21X1_34 ( );
FILL FILL_2_AOI21X1_34 ( );
FILL FILL_0_OAI21X1_818 ( );
FILL FILL_1_OAI21X1_818 ( );
FILL FILL_0_OAI21X1_817 ( );
FILL FILL_1_OAI21X1_817 ( );
FILL FILL_0_OAI21X1_816 ( );
FILL FILL_1_OAI21X1_816 ( );
FILL FILL_0_DFFPOSX1_521 ( );
FILL FILL_1_DFFPOSX1_521 ( );
FILL FILL_2_DFFPOSX1_521 ( );
FILL FILL_3_DFFPOSX1_521 ( );
FILL FILL_4_DFFPOSX1_521 ( );
FILL FILL_5_DFFPOSX1_521 ( );
FILL FILL_0_OAI21X1_600 ( );
FILL FILL_1_OAI21X1_600 ( );
FILL FILL_0_NAND3X1_19 ( );
FILL FILL_1_NAND3X1_19 ( );
FILL FILL_2_NAND3X1_19 ( );
FILL FILL_0_NAND2X1_293 ( );
FILL FILL_0_OAI21X1_598 ( );
FILL FILL_1_OAI21X1_598 ( );
FILL FILL_2_OAI21X1_598 ( );
FILL FILL_0_NOR2X1_83 ( );
FILL FILL_1_NOR2X1_83 ( );
FILL FILL_0_NAND2X1_294 ( );
FILL FILL_1_NAND2X1_294 ( );
FILL FILL_0_INVX2_48 ( );
FILL FILL_1_INVX2_48 ( );
FILL FILL_0_OAI21X1_597 ( );
FILL FILL_1_OAI21X1_597 ( );
FILL FILL_0_NAND2X1_326 ( );
FILL FILL_0_OAI21X1_755 ( );
FILL FILL_1_OAI21X1_755 ( );
FILL FILL_0_OAI21X1_789 ( );
FILL FILL_1_OAI21X1_789 ( );
FILL FILL_0_DFFPOSX1_593 ( );
FILL FILL_1_DFFPOSX1_593 ( );
FILL FILL_2_DFFPOSX1_593 ( );
FILL FILL_3_DFFPOSX1_593 ( );
FILL FILL_4_DFFPOSX1_593 ( );
FILL FILL_5_DFFPOSX1_593 ( );
FILL FILL_0_OAI21X1_723 ( );
FILL FILL_1_OAI21X1_723 ( );
FILL FILL_0_CLKBUF1_24 ( );
FILL FILL_1_CLKBUF1_24 ( );
FILL FILL_2_CLKBUF1_24 ( );
FILL FILL_3_CLKBUF1_24 ( );
FILL FILL_4_CLKBUF1_24 ( );
FILL FILL_0_INVX2_18 ( );
FILL FILL_0_DFFPOSX1_565 ( );
FILL FILL_1_DFFPOSX1_565 ( );
FILL FILL_2_DFFPOSX1_565 ( );
FILL FILL_3_DFFPOSX1_565 ( );
FILL FILL_4_DFFPOSX1_565 ( );
FILL FILL_5_DFFPOSX1_565 ( );
FILL FILL_0_INVX1_36 ( );
FILL FILL_0_AOI21X1_31 ( );
FILL FILL_1_AOI21X1_31 ( );
FILL FILL_2_AOI21X1_31 ( );
FILL FILL_0_INVX4_7 ( );
FILL FILL_0_NOR2X1_30 ( );
FILL FILL_0_OAI21X1_558 ( );
FILL FILL_1_OAI21X1_558 ( );
FILL FILL_2_OAI21X1_558 ( );
FILL FILL_0_NOR2X1_64 ( );
FILL FILL_0_OAI21X1_559 ( );
FILL FILL_1_OAI21X1_559 ( );
FILL FILL_0_NOR2X1_67 ( );
FILL FILL_0_OAI21X1_740 ( );
FILL FILL_1_OAI21X1_740 ( );
FILL FILL_0_DFFPOSX1_576 ( );
FILL FILL_1_DFFPOSX1_576 ( );
FILL FILL_2_DFFPOSX1_576 ( );
FILL FILL_3_DFFPOSX1_576 ( );
FILL FILL_4_DFFPOSX1_576 ( );
FILL FILL_5_DFFPOSX1_576 ( );
FILL FILL_0_NAND3X1_5 ( );
FILL FILL_1_NAND3X1_5 ( );
FILL FILL_2_NAND3X1_5 ( );
FILL FILL_0_NOR2X1_29 ( );
FILL FILL_0_NAND3X1_28 ( );
FILL FILL_1_NAND3X1_28 ( );
FILL FILL_2_NAND3X1_28 ( );
FILL FILL_0_INVX1_13 ( );
FILL FILL_0_NOR2X1_20 ( );
FILL FILL_0_NOR2X1_21 ( );
FILL FILL_1_NOR2X1_21 ( );
FILL FILL_0_OAI21X1_446 ( );
FILL FILL_1_OAI21X1_446 ( );
FILL FILL_0_OAI21X1_731 ( );
FILL FILL_1_OAI21X1_731 ( );
FILL FILL_0_INVX2_23 ( );
FILL FILL_0_INVX1_40 ( );
FILL FILL_0_AOI21X1_33 ( );
FILL FILL_1_AOI21X1_33 ( );
FILL FILL_0_INVX4_14 ( );
FILL FILL_0_BUFX2_604 ( );
FILL FILL_1_BUFX2_604 ( );
FILL FILL_0_OAI21X1_735 ( );
FILL FILL_1_OAI21X1_735 ( );
FILL FILL_0_OAI21X1_736 ( );
FILL FILL_1_OAI21X1_736 ( );
FILL FILL_0_OAI21X1_733 ( );
FILL FILL_1_OAI21X1_733 ( );
FILL FILL_2_OAI21X1_733 ( );
FILL FILL_0_DFFPOSX1_573 ( );
FILL FILL_1_DFFPOSX1_573 ( );
FILL FILL_2_DFFPOSX1_573 ( );
FILL FILL_3_DFFPOSX1_573 ( );
FILL FILL_4_DFFPOSX1_573 ( );
FILL FILL_5_DFFPOSX1_573 ( );
FILL FILL_0_OAI21X1_320 ( );
FILL FILL_1_OAI21X1_320 ( );
FILL FILL_0_OAI21X1_732 ( );
FILL FILL_1_OAI21X1_732 ( );
FILL FILL_0_BUFX2_12 ( );
FILL FILL_0_DFFPOSX1_579 ( );
FILL FILL_1_DFFPOSX1_579 ( );
FILL FILL_2_DFFPOSX1_579 ( );
FILL FILL_3_DFFPOSX1_579 ( );
FILL FILL_4_DFFPOSX1_579 ( );
FILL FILL_5_DFFPOSX1_579 ( );
FILL FILL_6_DFFPOSX1_579 ( );
FILL FILL_0_BUFX2_19 ( );
FILL FILL_1_BUFX2_19 ( );
FILL FILL_0_OAI21X1_1276 ( );
FILL FILL_1_OAI21X1_1276 ( );
FILL FILL_0_OAI21X1_1277 ( );
FILL FILL_1_OAI21X1_1277 ( );
FILL FILL_0_NAND2X1_601 ( );
FILL FILL_0_NAND3X1_53 ( );
FILL FILL_1_NAND3X1_53 ( );
FILL FILL_2_NAND3X1_53 ( );
FILL FILL_0_INVX1_202 ( );
FILL FILL_0_NAND2X1_514 ( );
FILL FILL_1_NAND2X1_514 ( );
FILL FILL_0_NOR2X1_186 ( );
FILL FILL_0_BUFX2_146 ( );
FILL FILL_1_BUFX2_146 ( );
FILL FILL_0_OAI21X1_1269 ( );
FILL FILL_1_OAI21X1_1269 ( );
FILL FILL_0_OAI21X1_1449 ( );
FILL FILL_1_OAI21X1_1449 ( );
FILL FILL_0_NOR2X1_222 ( );
FILL FILL_1_NOR2X1_222 ( );
FILL FILL_0_OAI21X1_1451 ( );
FILL FILL_1_OAI21X1_1451 ( );
FILL FILL_0_OAI21X1_1450 ( );
FILL FILL_1_OAI21X1_1450 ( );
FILL FILL_0_OAI21X1_1579 ( );
FILL FILL_1_OAI21X1_1579 ( );
FILL FILL_2_OAI21X1_1579 ( );
FILL FILL_0_OAI21X1_1271 ( );
FILL FILL_1_OAI21X1_1271 ( );
FILL FILL_2_OAI21X1_1271 ( );
FILL FILL_0_OAI21X1_1270 ( );
FILL FILL_1_OAI21X1_1270 ( );
FILL FILL_0_DFFPOSX1_893 ( );
FILL FILL_1_DFFPOSX1_893 ( );
FILL FILL_2_DFFPOSX1_893 ( );
FILL FILL_3_DFFPOSX1_893 ( );
FILL FILL_4_DFFPOSX1_893 ( );
FILL FILL_5_DFFPOSX1_893 ( );
FILL FILL_6_DFFPOSX1_893 ( );
FILL FILL_0_BUFX2_169 ( );
FILL FILL_1_BUFX2_169 ( );
FILL FILL_0_CLKBUF1_77 ( );
FILL FILL_1_CLKBUF1_77 ( );
FILL FILL_2_CLKBUF1_77 ( );
FILL FILL_3_CLKBUF1_77 ( );
FILL FILL_4_CLKBUF1_77 ( );
FILL FILL_0_OAI21X1_1495 ( );
FILL FILL_1_OAI21X1_1495 ( );
FILL FILL_0_OAI21X1_1496 ( );
FILL FILL_1_OAI21X1_1496 ( );
FILL FILL_0_DFFPOSX1_973 ( );
FILL FILL_1_DFFPOSX1_973 ( );
FILL FILL_2_DFFPOSX1_973 ( );
FILL FILL_3_DFFPOSX1_973 ( );
FILL FILL_4_DFFPOSX1_973 ( );
FILL FILL_5_DFFPOSX1_973 ( );
FILL FILL_6_DFFPOSX1_973 ( );
FILL FILL_0_INVX4_40 ( );
FILL FILL_1_INVX4_40 ( );
FILL FILL_0_INVX1_223 ( );
FILL FILL_0_NAND3X1_65 ( );
FILL FILL_1_NAND3X1_65 ( );
FILL FILL_0_OAI21X1_1157 ( );
FILL FILL_1_OAI21X1_1157 ( );
FILL FILL_0_NOR3X1_16 ( );
FILL FILL_1_NOR3X1_16 ( );
FILL FILL_2_NOR3X1_16 ( );
FILL FILL_3_NOR3X1_16 ( );
FILL FILL_4_NOR3X1_16 ( );
FILL FILL_0_OAI21X1_1507 ( );
FILL FILL_1_OAI21X1_1507 ( );
FILL FILL_0_OAI21X1_1506 ( );
FILL FILL_1_OAI21X1_1506 ( );
FILL FILL_0_BUFX4_239 ( );
FILL FILL_1_BUFX4_239 ( );
FILL FILL_0_OAI21X1_1540 ( );
FILL FILL_1_OAI21X1_1540 ( );
FILL FILL_0_DFFPOSX1_858 ( );
FILL FILL_1_DFFPOSX1_858 ( );
FILL FILL_2_DFFPOSX1_858 ( );
FILL FILL_3_DFFPOSX1_858 ( );
FILL FILL_4_DFFPOSX1_858 ( );
FILL FILL_5_DFFPOSX1_858 ( );
FILL FILL_6_DFFPOSX1_858 ( );
FILL FILL_0_NAND2X1_567 ( );
FILL FILL_0_OAI21X1_1180 ( );
FILL FILL_1_OAI21X1_1180 ( );
FILL FILL_0_INVX4_44 ( );
FILL FILL_0_OAI21X1_1509 ( );
FILL FILL_1_OAI21X1_1509 ( );
FILL FILL_2_OAI21X1_1509 ( );
FILL FILL_0_DFFPOSX1_977 ( );
FILL FILL_1_DFFPOSX1_977 ( );
FILL FILL_2_DFFPOSX1_977 ( );
FILL FILL_3_DFFPOSX1_977 ( );
FILL FILL_4_DFFPOSX1_977 ( );
FILL FILL_5_DFFPOSX1_977 ( );
FILL FILL_0_OAI21X1_1508 ( );
FILL FILL_1_OAI21X1_1508 ( );
FILL FILL_0_OAI21X1_1354 ( );
FILL FILL_1_OAI21X1_1354 ( );
FILL FILL_0_OAI21X1_1353 ( );
FILL FILL_1_OAI21X1_1353 ( );
FILL FILL_2_OAI21X1_1353 ( );
FILL FILL_0_NOR2X1_210 ( );
FILL FILL_0_NAND2X1_566 ( );
FILL FILL_1_NAND2X1_566 ( );
FILL FILL_0_OAI21X1_1179 ( );
FILL FILL_1_OAI21X1_1179 ( );
FILL FILL_0_DFFPOSX1_857 ( );
FILL FILL_1_DFFPOSX1_857 ( );
FILL FILL_2_DFFPOSX1_857 ( );
FILL FILL_3_DFFPOSX1_857 ( );
FILL FILL_4_DFFPOSX1_857 ( );
FILL FILL_5_DFFPOSX1_857 ( );
FILL FILL_0_BUFX2_178 ( );
FILL FILL_0_BUFX2_231 ( );
FILL FILL_1_BUFX2_231 ( );
FILL FILL_0_BUFX2_109 ( );
FILL FILL_1_BUFX2_109 ( );
FILL FILL_0_BUFX2_111 ( );
FILL FILL_0_OAI21X1_1377 ( );
FILL FILL_1_OAI21X1_1377 ( );
FILL FILL_0_OAI21X1_1378 ( );
FILL FILL_1_OAI21X1_1378 ( );
FILL FILL_0_OAI21X1_1376 ( );
FILL FILL_1_OAI21X1_1376 ( );
FILL FILL_0_DFFPOSX1_933 ( );
FILL FILL_1_DFFPOSX1_933 ( );
FILL FILL_2_DFFPOSX1_933 ( );
FILL FILL_3_DFFPOSX1_933 ( );
FILL FILL_4_DFFPOSX1_933 ( );
FILL FILL_5_DFFPOSX1_933 ( );
FILL FILL_0_BUFX4_188 ( );
FILL FILL_1_BUFX4_188 ( );
FILL FILL_0_DFFPOSX1_804 ( );
FILL FILL_1_DFFPOSX1_804 ( );
FILL FILL_2_DFFPOSX1_804 ( );
FILL FILL_3_DFFPOSX1_804 ( );
FILL FILL_4_DFFPOSX1_804 ( );
FILL FILL_5_DFFPOSX1_804 ( );
FILL FILL_6_DFFPOSX1_804 ( );
FILL FILL_0_BUFX2_58 ( );
FILL FILL_1_BUFX2_58 ( );
FILL FILL_0_BUFX2_122 ( );
FILL FILL_1_BUFX2_122 ( );
FILL FILL_0_DFFPOSX1_65 ( );
FILL FILL_1_DFFPOSX1_65 ( );
FILL FILL_2_DFFPOSX1_65 ( );
FILL FILL_3_DFFPOSX1_65 ( );
FILL FILL_4_DFFPOSX1_65 ( );
FILL FILL_5_DFFPOSX1_65 ( );
FILL FILL_6_DFFPOSX1_65 ( );
FILL FILL_0_OAI21X1_1751 ( );
FILL FILL_1_OAI21X1_1751 ( );
FILL FILL_0_DFFPOSX1_88 ( );
FILL FILL_1_DFFPOSX1_88 ( );
FILL FILL_2_DFFPOSX1_88 ( );
FILL FILL_3_DFFPOSX1_88 ( );
FILL FILL_4_DFFPOSX1_88 ( );
FILL FILL_5_DFFPOSX1_88 ( );
FILL FILL_0_OAI21X1_952 ( );
FILL FILL_1_OAI21X1_952 ( );
FILL FILL_0_NAND2X1_47 ( );
FILL FILL_1_NAND2X1_47 ( );
FILL FILL_0_BUFX2_938 ( );
FILL FILL_1_BUFX2_938 ( );
FILL FILL_0_BUFX2_248 ( );
FILL FILL_0_BUFX2_874 ( );
FILL FILL_1_BUFX2_874 ( );
FILL FILL_0_INVX2_121 ( );
FILL FILL_0_BUFX2_956 ( );
FILL FILL_0_INVX2_201 ( );
FILL FILL_0_DFFPOSX1_1008 ( );
FILL FILL_1_DFFPOSX1_1008 ( );
FILL FILL_2_DFFPOSX1_1008 ( );
FILL FILL_3_DFFPOSX1_1008 ( );
FILL FILL_4_DFFPOSX1_1008 ( );
FILL FILL_5_DFFPOSX1_1008 ( );
FILL FILL_6_DFFPOSX1_1008 ( );
FILL FILL_0_OAI21X1_1585 ( );
FILL FILL_1_OAI21X1_1585 ( );
FILL FILL_2_OAI21X1_1585 ( );
FILL FILL_0_DFFPOSX1_347 ( );
FILL FILL_1_DFFPOSX1_347 ( );
FILL FILL_2_DFFPOSX1_347 ( );
FILL FILL_3_DFFPOSX1_347 ( );
FILL FILL_4_DFFPOSX1_347 ( );
FILL FILL_5_DFFPOSX1_347 ( );
FILL FILL_6_DFFPOSX1_347 ( );
FILL FILL_0_OAI21X1_311 ( );
FILL FILL_1_OAI21X1_311 ( );
FILL FILL_2_OAI21X1_311 ( );
FILL FILL_0_OAI21X1_310 ( );
FILL FILL_1_OAI21X1_310 ( );
FILL FILL_0_INVX2_5 ( );
FILL FILL_0_OAI21X1_624 ( );
FILL FILL_1_OAI21X1_624 ( );
FILL FILL_0_DFFPOSX1_422 ( );
FILL FILL_1_DFFPOSX1_422 ( );
FILL FILL_2_DFFPOSX1_422 ( );
FILL FILL_3_DFFPOSX1_422 ( );
FILL FILL_4_DFFPOSX1_422 ( );
FILL FILL_5_DFFPOSX1_422 ( );
FILL FILL_0_NAND2X1_140 ( );
FILL FILL_0_OAI21X1_396 ( );
FILL FILL_1_OAI21X1_396 ( );
FILL FILL_2_OAI21X1_396 ( );
FILL FILL_0_OAI21X1_78 ( );
FILL FILL_1_OAI21X1_78 ( );
FILL FILL_0_OAI21X1_79 ( );
FILL FILL_1_OAI21X1_79 ( );
FILL FILL_0_OAI21X1_395 ( );
FILL FILL_1_OAI21X1_395 ( );
FILL FILL_0_OAI21X1_394 ( );
FILL FILL_1_OAI21X1_394 ( );
FILL FILL_0_DFFPOSX1_486 ( );
FILL FILL_1_DFFPOSX1_486 ( );
FILL FILL_2_DFFPOSX1_486 ( );
FILL FILL_3_DFFPOSX1_486 ( );
FILL FILL_4_DFFPOSX1_486 ( );
FILL FILL_5_DFFPOSX1_486 ( );
FILL FILL_6_DFFPOSX1_486 ( );
FILL FILL_0_NAND2X1_267 ( );
FILL FILL_1_NAND2X1_267 ( );
FILL FILL_0_OAI21X1_505 ( );
FILL FILL_1_OAI21X1_505 ( );
FILL FILL_0_NAND2X1_74 ( );
FILL FILL_1_NAND2X1_74 ( );
FILL FILL_0_OAI21X1_504 ( );
FILL FILL_1_OAI21X1_504 ( );
FILL FILL_0_DFFPOSX1_358 ( );
FILL FILL_1_DFFPOSX1_358 ( );
FILL FILL_2_DFFPOSX1_358 ( );
FILL FILL_3_DFFPOSX1_358 ( );
FILL FILL_4_DFFPOSX1_358 ( );
FILL FILL_5_DFFPOSX1_358 ( );
FILL FILL_6_DFFPOSX1_358 ( );
FILL FILL_0_NAND2X1_112 ( );
FILL FILL_1_NAND2X1_112 ( );
FILL FILL_0_BUFX2_622 ( );
FILL FILL_1_BUFX2_622 ( );
FILL FILL_0_BUFX4_7 ( );
FILL FILL_1_BUFX4_7 ( );
FILL FILL_2_BUFX4_7 ( );
FILL FILL_0_OAI21X1_777 ( );
FILL FILL_1_OAI21X1_777 ( );
FILL FILL_0_BUFX4_69 ( );
FILL FILL_1_BUFX4_69 ( );
FILL FILL_0_BUFX4_135 ( );
FILL FILL_1_BUFX4_135 ( );
FILL FILL_0_BUFX2_621 ( );
FILL FILL_1_BUFX2_621 ( );
FILL FILL_0_DFFPOSX1_589 ( );
FILL FILL_1_DFFPOSX1_589 ( );
FILL FILL_2_DFFPOSX1_589 ( );
FILL FILL_3_DFFPOSX1_589 ( );
FILL FILL_4_DFFPOSX1_589 ( );
FILL FILL_5_DFFPOSX1_589 ( );
FILL FILL_0_OAI21X1_773 ( );
FILL FILL_1_OAI21X1_773 ( );
FILL FILL_0_OAI21X1_774 ( );
FILL FILL_1_OAI21X1_774 ( );
FILL FILL_0_NAND2X1_116 ( );
FILL FILL_0_OAI21X1_372 ( );
FILL FILL_1_OAI21X1_372 ( );
FILL FILL_0_INVX2_29 ( );
FILL FILL_0_XNOR2X1_25 ( );
FILL FILL_1_XNOR2X1_25 ( );
FILL FILL_2_XNOR2X1_25 ( );
FILL FILL_3_XNOR2X1_25 ( );
FILL FILL_0_XNOR2X1_52 ( );
FILL FILL_1_XNOR2X1_52 ( );
FILL FILL_2_XNOR2X1_52 ( );
FILL FILL_3_XNOR2X1_52 ( );
FILL FILL_0_DFFPOSX1_531 ( );
FILL FILL_1_DFFPOSX1_531 ( );
FILL FILL_2_DFFPOSX1_531 ( );
FILL FILL_3_DFFPOSX1_531 ( );
FILL FILL_4_DFFPOSX1_531 ( );
FILL FILL_5_DFFPOSX1_531 ( );
FILL FILL_6_DFFPOSX1_531 ( );
FILL FILL_0_NAND3X1_31 ( );
FILL FILL_1_NAND3X1_31 ( );
FILL FILL_0_NOR2X1_87 ( );
FILL FILL_0_INVX2_32 ( );
FILL FILL_0_NOR3X1_2 ( );
FILL FILL_1_NOR3X1_2 ( );
FILL FILL_2_NOR3X1_2 ( );
FILL FILL_3_NOR3X1_2 ( );
FILL FILL_4_NOR3X1_2 ( );
FILL FILL_0_OAI21X1_465 ( );
FILL FILL_1_OAI21X1_465 ( );
FILL FILL_0_BUFX4_20 ( );
FILL FILL_1_BUFX4_20 ( );
FILL FILL_2_BUFX4_20 ( );
FILL FILL_0_OR2X2_11 ( );
FILL FILL_1_OR2X2_11 ( );
FILL FILL_0_AOI21X1_17 ( );
FILL FILL_1_AOI21X1_17 ( );
FILL FILL_0_BUFX4_122 ( );
FILL FILL_1_BUFX4_122 ( );
FILL FILL_0_BUFX4_13 ( );
FILL FILL_1_BUFX4_13 ( );
FILL FILL_0_INVX4_24 ( );
FILL FILL_1_INVX4_24 ( );
FILL FILL_0_NAND3X1_34 ( );
FILL FILL_1_NAND3X1_34 ( );
FILL FILL_0_NAND2X1_332 ( );
FILL FILL_1_NAND2X1_332 ( );
FILL FILL_0_OAI21X1_820 ( );
FILL FILL_1_OAI21X1_820 ( );
FILL FILL_0_XNOR2X1_54 ( );
FILL FILL_1_XNOR2X1_54 ( );
FILL FILL_2_XNOR2X1_54 ( );
FILL FILL_3_XNOR2X1_54 ( );
FILL FILL_0_DFFPOSX1_538 ( );
FILL FILL_1_DFFPOSX1_538 ( );
FILL FILL_2_DFFPOSX1_538 ( );
FILL FILL_3_DFFPOSX1_538 ( );
FILL FILL_4_DFFPOSX1_538 ( );
FILL FILL_5_DFFPOSX1_538 ( );
FILL FILL_6_DFFPOSX1_538 ( );
FILL FILL_0_OAI21X1_636 ( );
FILL FILL_1_OAI21X1_636 ( );
FILL FILL_0_NAND2X1_324 ( );
FILL FILL_1_NAND2X1_324 ( );
FILL FILL_0_NOR3X1_6 ( );
FILL FILL_1_NOR3X1_6 ( );
FILL FILL_2_NOR3X1_6 ( );
FILL FILL_3_NOR3X1_6 ( );
FILL FILL_0_NOR2X1_78 ( );
FILL FILL_0_OR2X2_9 ( );
FILL FILL_1_OR2X2_9 ( );
FILL FILL_0_AOI21X1_11 ( );
FILL FILL_1_AOI21X1_11 ( );
FILL FILL_0_NAND3X1_20 ( );
FILL FILL_1_NAND3X1_20 ( );
FILL FILL_0_INVX1_30 ( );
FILL FILL_0_AOI21X1_10 ( );
FILL FILL_1_AOI21X1_10 ( );
FILL FILL_0_NOR2X1_80 ( );
FILL FILL_1_NOR2X1_80 ( );
FILL FILL_0_NAND2X1_292 ( );
FILL FILL_1_NAND2X1_292 ( );
FILL FILL_0_OR2X2_10 ( );
FILL FILL_1_OR2X2_10 ( );
FILL FILL_0_BUFX4_84 ( );
FILL FILL_1_BUFX4_84 ( );
FILL FILL_0_BUFX4_177 ( );
FILL FILL_1_BUFX4_177 ( );
FILL FILL_0_NOR2X1_113 ( );
FILL FILL_1_NOR2X1_113 ( );
FILL FILL_0_AND2X2_21 ( );
FILL FILL_1_AND2X2_21 ( );
FILL FILL_0_OAI21X1_766 ( );
FILL FILL_1_OAI21X1_766 ( );
FILL FILL_0_OAI21X1_767 ( );
FILL FILL_1_OAI21X1_767 ( );
FILL FILL_0_INVX1_42 ( );
FILL FILL_0_OAI21X1_707 ( );
FILL FILL_1_OAI21X1_707 ( );
FILL FILL_0_OAI21X1_708 ( );
FILL FILL_1_OAI21X1_708 ( );
FILL FILL_0_XNOR2X1_43 ( );
FILL FILL_1_XNOR2X1_43 ( );
FILL FILL_2_XNOR2X1_43 ( );
FILL FILL_3_XNOR2X1_43 ( );
FILL FILL_0_OAI21X1_207 ( );
FILL FILL_1_OAI21X1_207 ( );
FILL FILL_2_OAI21X1_207 ( );
FILL FILL_0_DFFPOSX1_504 ( );
FILL FILL_1_DFFPOSX1_504 ( );
FILL FILL_2_DFFPOSX1_504 ( );
FILL FILL_3_DFFPOSX1_504 ( );
FILL FILL_4_DFFPOSX1_504 ( );
FILL FILL_5_DFFPOSX1_504 ( );
FILL FILL_0_OAI21X1_206 ( );
FILL FILL_1_OAI21X1_206 ( );
FILL FILL_0_NOR2X1_82 ( );
FILL FILL_1_NOR2X1_82 ( );
FILL FILL_0_NAND3X1_18 ( );
FILL FILL_1_NAND3X1_18 ( );
FILL FILL_0_NAND3X1_21 ( );
FILL FILL_1_NAND3X1_21 ( );
FILL FILL_0_AND2X2_14 ( );
FILL FILL_1_AND2X2_14 ( );
FILL FILL_0_NAND2X1_284 ( );
FILL FILL_1_NAND2X1_284 ( );
FILL FILL_0_NAND2X1_282 ( );
FILL FILL_0_INVX1_27 ( );
FILL FILL_0_NAND2X1_201 ( );
FILL FILL_1_NAND2X1_201 ( );
FILL FILL_0_AOI21X1_2 ( );
FILL FILL_1_AOI21X1_2 ( );
FILL FILL_0_AND2X2_6 ( );
FILL FILL_1_AND2X2_6 ( );
FILL FILL_0_XNOR2X1_48 ( );
FILL FILL_1_XNOR2X1_48 ( );
FILL FILL_2_XNOR2X1_48 ( );
FILL FILL_0_NOR3X1_7 ( );
FILL FILL_1_NOR3X1_7 ( );
FILL FILL_2_NOR3X1_7 ( );
FILL FILL_3_NOR3X1_7 ( );
FILL FILL_0_OAI21X1_746 ( );
FILL FILL_1_OAI21X1_746 ( );
FILL FILL_0_OAI21X1_734 ( );
FILL FILL_1_OAI21X1_734 ( );
FILL FILL_2_OAI21X1_734 ( );
FILL FILL_0_DFFPOSX1_574 ( );
FILL FILL_1_DFFPOSX1_574 ( );
FILL FILL_2_DFFPOSX1_574 ( );
FILL FILL_3_DFFPOSX1_574 ( );
FILL FILL_4_DFFPOSX1_574 ( );
FILL FILL_5_DFFPOSX1_574 ( );
FILL FILL_0_OAI21X1_819 ( );
FILL FILL_1_OAI21X1_819 ( );
FILL FILL_2_OAI21X1_819 ( );
FILL FILL_0_OAI21X1_821 ( );
FILL FILL_1_OAI21X1_821 ( );
FILL FILL_0_BUFX4_275 ( );
FILL FILL_1_BUFX4_275 ( );
FILL FILL_0_DFFPOSX1_603 ( );
FILL FILL_1_DFFPOSX1_603 ( );
FILL FILL_2_DFFPOSX1_603 ( );
FILL FILL_3_DFFPOSX1_603 ( );
FILL FILL_4_DFFPOSX1_603 ( );
FILL FILL_5_DFFPOSX1_603 ( );
FILL FILL_6_DFFPOSX1_603 ( );
FILL FILL_0_INVX1_39 ( );
FILL FILL_0_OAI21X1_747 ( );
FILL FILL_1_OAI21X1_747 ( );
FILL FILL_0_DFFPOSX1_161 ( );
FILL FILL_1_DFFPOSX1_161 ( );
FILL FILL_2_DFFPOSX1_161 ( );
FILL FILL_3_DFFPOSX1_161 ( );
FILL FILL_4_DFFPOSX1_161 ( );
FILL FILL_5_DFFPOSX1_161 ( );
FILL FILL_6_DFFPOSX1_161 ( );
FILL FILL_0_OAI21X1_5 ( );
FILL FILL_1_OAI21X1_5 ( );
FILL FILL_0_NAND2X1_5 ( );
FILL FILL_1_NAND2X1_5 ( );
FILL FILL_0_DFFPOSX1_896 ( );
FILL FILL_1_DFFPOSX1_896 ( );
FILL FILL_2_DFFPOSX1_896 ( );
FILL FILL_3_DFFPOSX1_896 ( );
FILL FILL_4_DFFPOSX1_896 ( );
FILL FILL_5_DFFPOSX1_896 ( );
FILL FILL_0_BUFX4_324 ( );
FILL FILL_1_BUFX4_324 ( );
FILL FILL_2_BUFX4_324 ( );
FILL FILL_0_BUFX4_16 ( );
FILL FILL_1_BUFX4_16 ( );
FILL FILL_0_OAI21X1_1278 ( );
FILL FILL_1_OAI21X1_1278 ( );
FILL FILL_2_OAI21X1_1278 ( );
FILL FILL_0_OAI21X1_1580 ( );
FILL FILL_1_OAI21X1_1580 ( );
FILL FILL_0_BUFX4_88 ( );
FILL FILL_1_BUFX4_88 ( );
FILL FILL_0_BUFX2_210 ( );
FILL FILL_1_BUFX2_210 ( );
FILL FILL_0_OAI21X1_1331 ( );
FILL FILL_1_OAI21X1_1331 ( );
FILL FILL_0_DFFPOSX1_917 ( );
FILL FILL_1_DFFPOSX1_917 ( );
FILL FILL_2_DFFPOSX1_917 ( );
FILL FILL_3_DFFPOSX1_917 ( );
FILL FILL_4_DFFPOSX1_917 ( );
FILL FILL_5_DFFPOSX1_917 ( );
FILL FILL_6_DFFPOSX1_917 ( );
FILL FILL_0_OAI21X1_1332 ( );
FILL FILL_1_OAI21X1_1332 ( );
FILL FILL_0_DFFPOSX1_49 ( );
FILL FILL_1_DFFPOSX1_49 ( );
FILL FILL_2_DFFPOSX1_49 ( );
FILL FILL_3_DFFPOSX1_49 ( );
FILL FILL_4_DFFPOSX1_49 ( );
FILL FILL_5_DFFPOSX1_49 ( );
FILL FILL_0_NAND2X1_436 ( );
FILL FILL_0_BUFX4_286 ( );
FILL FILL_1_BUFX4_286 ( );
FILL FILL_0_CLKBUF1_85 ( );
FILL FILL_1_CLKBUF1_85 ( );
FILL FILL_2_CLKBUF1_85 ( );
FILL FILL_3_CLKBUF1_85 ( );
FILL FILL_4_CLKBUF1_85 ( );
FILL FILL_0_INVX2_106 ( );
FILL FILL_0_BUFX2_29 ( );
FILL FILL_1_BUFX2_29 ( );
FILL FILL_0_NAND2X1_614 ( );
FILL FILL_0_OAI21X1_1483 ( );
FILL FILL_1_OAI21X1_1483 ( );
FILL FILL_0_NOR2X1_201 ( );
FILL FILL_1_NOR2X1_201 ( );
FILL FILL_0_NAND2X1_613 ( );
FILL FILL_0_BUFX4_21 ( );
FILL FILL_1_BUFX4_21 ( );
FILL FILL_0_BUFX4_212 ( );
FILL FILL_1_BUFX4_212 ( );
FILL FILL_0_BUFX4_89 ( );
FILL FILL_1_BUFX4_89 ( );
FILL FILL_0_DFFPOSX1_850 ( );
FILL FILL_1_DFFPOSX1_850 ( );
FILL FILL_2_DFFPOSX1_850 ( );
FILL FILL_3_DFFPOSX1_850 ( );
FILL FILL_4_DFFPOSX1_850 ( );
FILL FILL_5_DFFPOSX1_850 ( );
FILL FILL_6_DFFPOSX1_850 ( );
FILL FILL_0_NAND2X1_550 ( );
FILL FILL_0_BUFX2_166 ( );
FILL FILL_1_BUFX2_166 ( );
FILL FILL_0_OAI21X1_1181 ( );
FILL FILL_1_OAI21X1_1181 ( );
FILL FILL_2_OAI21X1_1181 ( );
FILL FILL_0_BUFX4_303 ( );
FILL FILL_1_BUFX4_303 ( );
FILL FILL_0_NOR2X1_167 ( );
FILL FILL_1_NOR2X1_167 ( );
FILL FILL_0_OAI21X1_1345 ( );
FILL FILL_1_OAI21X1_1345 ( );
FILL FILL_0_BUFX2_175 ( );
FILL FILL_1_BUFX2_175 ( );
FILL FILL_0_NAND2X1_581 ( );
FILL FILL_1_NAND2X1_581 ( );
FILL FILL_0_OAI21X1_1196 ( );
FILL FILL_1_OAI21X1_1196 ( );
FILL FILL_0_DFFPOSX1_925 ( );
FILL FILL_1_DFFPOSX1_925 ( );
FILL FILL_2_DFFPOSX1_925 ( );
FILL FILL_3_DFFPOSX1_925 ( );
FILL FILL_4_DFFPOSX1_925 ( );
FILL FILL_5_DFFPOSX1_925 ( );
FILL FILL_0_OAI21X1_1369 ( );
FILL FILL_1_OAI21X1_1369 ( );
FILL FILL_2_OAI21X1_1369 ( );
FILL FILL_0_INVX1_216 ( );
FILL FILL_0_OAI21X1_1368 ( );
FILL FILL_1_OAI21X1_1368 ( );
FILL FILL_0_NAND2X1_562 ( );
FILL FILL_1_NAND2X1_562 ( );
FILL FILL_0_BUFX4_187 ( );
FILL FILL_1_BUFX4_187 ( );
FILL FILL_0_OAI21X1_1513 ( );
FILL FILL_1_OAI21X1_1513 ( );
FILL FILL_0_BUFX4_357 ( );
FILL FILL_1_BUFX4_357 ( );
FILL FILL_0_DFFPOSX1_868 ( );
FILL FILL_1_DFFPOSX1_868 ( );
FILL FILL_2_DFFPOSX1_868 ( );
FILL FILL_3_DFFPOSX1_868 ( );
FILL FILL_4_DFFPOSX1_868 ( );
FILL FILL_5_DFFPOSX1_868 ( );
FILL FILL_0_NAND2X1_584 ( );
FILL FILL_1_NAND2X1_584 ( );
FILL FILL_0_DFFPOSX1_867 ( );
FILL FILL_1_DFFPOSX1_867 ( );
FILL FILL_2_DFFPOSX1_867 ( );
FILL FILL_3_DFFPOSX1_867 ( );
FILL FILL_4_DFFPOSX1_867 ( );
FILL FILL_5_DFFPOSX1_867 ( );
FILL FILL_6_DFFPOSX1_867 ( );
FILL FILL_0_NAND2X1_583 ( );
FILL FILL_0_OAI21X1_1096 ( );
FILL FILL_1_OAI21X1_1096 ( );
FILL FILL_0_NAND2X1_462 ( );
FILL FILL_1_NAND2X1_462 ( );
FILL FILL_0_DFFPOSX1_995 ( );
FILL FILL_1_DFFPOSX1_995 ( );
FILL FILL_2_DFFPOSX1_995 ( );
FILL FILL_3_DFFPOSX1_995 ( );
FILL FILL_4_DFFPOSX1_995 ( );
FILL FILL_5_DFFPOSX1_995 ( );
FILL FILL_6_DFFPOSX1_995 ( );
FILL FILL_0_OAI21X1_1561 ( );
FILL FILL_1_OAI21X1_1561 ( );
FILL FILL_0_BUFX4_141 ( );
FILL FILL_1_BUFX4_141 ( );
FILL FILL_0_DFFPOSX1_267 ( );
FILL FILL_1_DFFPOSX1_267 ( );
FILL FILL_2_DFFPOSX1_267 ( );
FILL FILL_3_DFFPOSX1_267 ( );
FILL FILL_4_DFFPOSX1_267 ( );
FILL FILL_5_DFFPOSX1_267 ( );
FILL FILL_6_DFFPOSX1_267 ( );
FILL FILL_0_OAI21X1_151 ( );
FILL FILL_1_OAI21X1_151 ( );
FILL FILL_0_OAI21X1_150 ( );
FILL FILL_1_OAI21X1_150 ( );
FILL FILL_0_OAI21X1_47 ( );
FILL FILL_1_OAI21X1_47 ( );
FILL FILL_0_DFFPOSX1_203 ( );
FILL FILL_1_DFFPOSX1_203 ( );
FILL FILL_2_DFFPOSX1_203 ( );
FILL FILL_3_DFFPOSX1_203 ( );
FILL FILL_4_DFFPOSX1_203 ( );
FILL FILL_5_DFFPOSX1_203 ( );
FILL FILL_0_INVX1_124 ( );
FILL FILL_0_BUFX2_332 ( );
FILL FILL_0_BUFX2_262 ( );
FILL FILL_1_BUFX2_262 ( );
FILL FILL_0_INVX1_46 ( );
FILL FILL_0_OAI21X1_845 ( );
FILL FILL_1_OAI21X1_845 ( );
FILL FILL_0_BUFX2_771 ( );
FILL FILL_0_BUFX2_707 ( );
FILL FILL_1_BUFX2_707 ( );
FILL FILL_0_OAI21X1_182 ( );
FILL FILL_1_OAI21X1_182 ( );
FILL FILL_0_OAI21X1_183 ( );
FILL FILL_1_OAI21X1_183 ( );
FILL FILL_0_DFFPOSX1_283 ( );
FILL FILL_1_DFFPOSX1_283 ( );
FILL FILL_2_DFFPOSX1_283 ( );
FILL FILL_3_DFFPOSX1_283 ( );
FILL FILL_4_DFFPOSX1_283 ( );
FILL FILL_5_DFFPOSX1_283 ( );
FILL FILL_0_OAI21X1_1718 ( );
FILL FILL_1_OAI21X1_1718 ( );
FILL FILL_0_DFFPOSX1_533 ( );
FILL FILL_1_DFFPOSX1_533 ( );
FILL FILL_2_DFFPOSX1_533 ( );
FILL FILL_3_DFFPOSX1_533 ( );
FILL FILL_4_DFFPOSX1_533 ( );
FILL FILL_5_DFFPOSX1_533 ( );
FILL FILL_6_DFFPOSX1_533 ( );
FILL FILL_0_OAI21X1_625 ( );
FILL FILL_1_OAI21X1_625 ( );
FILL FILL_0_BUFX4_176 ( );
FILL FILL_1_BUFX4_176 ( );
FILL FILL_2_BUFX4_176 ( );
FILL FILL_0_CLKBUF1_4 ( );
FILL FILL_1_CLKBUF1_4 ( );
FILL FILL_2_CLKBUF1_4 ( );
FILL FILL_3_CLKBUF1_4 ( );
FILL FILL_0_DFFPOSX1_231 ( );
FILL FILL_1_DFFPOSX1_231 ( );
FILL FILL_2_DFFPOSX1_231 ( );
FILL FILL_3_DFFPOSX1_231 ( );
FILL FILL_4_DFFPOSX1_231 ( );
FILL FILL_5_DFFPOSX1_231 ( );
FILL FILL_0_BUFX2_521 ( );
FILL FILL_0_OAI21X1_691 ( );
FILL FILL_1_OAI21X1_691 ( );
FILL FILL_0_DFFPOSX1_559 ( );
FILL FILL_1_DFFPOSX1_559 ( );
FILL FILL_2_DFFPOSX1_559 ( );
FILL FILL_3_DFFPOSX1_559 ( );
FILL FILL_4_DFFPOSX1_559 ( );
FILL FILL_5_DFFPOSX1_559 ( );
FILL FILL_6_DFFPOSX1_559 ( );
FILL FILL_0_OAI21X1_692 ( );
FILL FILL_1_OAI21X1_692 ( );
FILL FILL_0_BUFX2_597 ( );
FILL FILL_0_OAI21X1_664 ( );
FILL FILL_1_OAI21X1_664 ( );
FILL FILL_0_OAI21X1_665 ( );
FILL FILL_1_OAI21X1_665 ( );
FILL FILL_0_DFFPOSX1_550 ( );
FILL FILL_1_DFFPOSX1_550 ( );
FILL FILL_2_DFFPOSX1_550 ( );
FILL FILL_3_DFFPOSX1_550 ( );
FILL FILL_4_DFFPOSX1_550 ( );
FILL FILL_5_DFFPOSX1_550 ( );
FILL FILL_0_BUFX2_494 ( );
FILL FILL_1_BUFX2_494 ( );
FILL FILL_0_BUFX2_560 ( );
FILL FILL_0_DFFPOSX1_590 ( );
FILL FILL_1_DFFPOSX1_590 ( );
FILL FILL_2_DFFPOSX1_590 ( );
FILL FILL_3_DFFPOSX1_590 ( );
FILL FILL_4_DFFPOSX1_590 ( );
FILL FILL_5_DFFPOSX1_590 ( );
FILL FILL_6_DFFPOSX1_590 ( );
FILL FILL_0_OAI21X1_778 ( );
FILL FILL_1_OAI21X1_778 ( );
FILL FILL_0_CLKBUF1_90 ( );
FILL FILL_1_CLKBUF1_90 ( );
FILL FILL_2_CLKBUF1_90 ( );
FILL FILL_3_CLKBUF1_90 ( );
FILL FILL_4_CLKBUF1_90 ( );
FILL FILL_0_DFFPOSX1_462 ( );
FILL FILL_1_DFFPOSX1_462 ( );
FILL FILL_2_DFFPOSX1_462 ( );
FILL FILL_3_DFFPOSX1_462 ( );
FILL FILL_4_DFFPOSX1_462 ( );
FILL FILL_5_DFFPOSX1_462 ( );
FILL FILL_6_DFFPOSX1_462 ( );
FILL FILL_0_BUFX4_76 ( );
FILL FILL_1_BUFX4_76 ( );
FILL FILL_0_NAND2X1_230 ( );
FILL FILL_0_BUFX4_37 ( );
FILL FILL_1_BUFX4_37 ( );
FILL FILL_0_NAND2X1_295 ( );
FILL FILL_1_NAND2X1_295 ( );
FILL FILL_0_NOR2X1_86 ( );
FILL FILL_0_NAND2X1_221 ( );
FILL FILL_1_NAND2X1_221 ( );
FILL FILL_0_NAND3X1_8 ( );
FILL FILL_1_NAND3X1_8 ( );
FILL FILL_2_NAND3X1_8 ( );
FILL FILL_0_OAI21X1_776 ( );
FILL FILL_1_OAI21X1_776 ( );
FILL FILL_2_OAI21X1_776 ( );
FILL FILL_0_OAI21X1_783 ( );
FILL FILL_1_OAI21X1_783 ( );
FILL FILL_2_OAI21X1_783 ( );
FILL FILL_0_INVX4_31 ( );
FILL FILL_1_INVX4_31 ( );
FILL FILL_0_NOR2X1_114 ( );
FILL FILL_0_NAND2X1_330 ( );
FILL FILL_0_INVX2_49 ( );
FILL FILL_0_NOR2X1_90 ( );
FILL FILL_1_NOR2X1_90 ( );
FILL FILL_0_NAND3X1_23 ( );
FILL FILL_1_NAND3X1_23 ( );
FILL FILL_0_NOR3X1_3 ( );
FILL FILL_1_NOR3X1_3 ( );
FILL FILL_2_NOR3X1_3 ( );
FILL FILL_3_NOR3X1_3 ( );
FILL FILL_4_NOR3X1_3 ( );
FILL FILL_0_BUFX2_442 ( );
FILL FILL_1_BUFX2_442 ( );
FILL FILL_0_NOR2X1_41 ( );
FILL FILL_1_NOR2X1_41 ( );
FILL FILL_0_NAND2X1_233 ( );
FILL FILL_1_NAND2X1_233 ( );
FILL FILL_0_OAI21X1_801 ( );
FILL FILL_1_OAI21X1_801 ( );
FILL FILL_0_OAI21X1_800 ( );
FILL FILL_1_OAI21X1_800 ( );
FILL FILL_0_INVX2_35 ( );
FILL FILL_0_NAND2X1_249 ( );
FILL FILL_0_AOI21X1_20 ( );
FILL FILL_1_AOI21X1_20 ( );
FILL FILL_2_AOI21X1_20 ( );
FILL FILL_0_NOR2X1_91 ( );
FILL FILL_1_NOR2X1_91 ( );
FILL FILL_0_NAND3X1_22 ( );
FILL FILL_1_NAND3X1_22 ( );
FILL FILL_0_INVX1_31 ( );
FILL FILL_0_NOR3X1_9 ( );
FILL FILL_1_NOR3X1_9 ( );
FILL FILL_2_NOR3X1_9 ( );
FILL FILL_3_NOR3X1_9 ( );
FILL FILL_0_OAI21X1_637 ( );
FILL FILL_1_OAI21X1_637 ( );
FILL FILL_0_DFFPOSX1_520 ( );
FILL FILL_1_DFFPOSX1_520 ( );
FILL FILL_2_DFFPOSX1_520 ( );
FILL FILL_3_DFFPOSX1_520 ( );
FILL FILL_4_DFFPOSX1_520 ( );
FILL FILL_5_DFFPOSX1_520 ( );
FILL FILL_6_DFFPOSX1_520 ( );
FILL FILL_0_OAI21X1_595 ( );
FILL FILL_1_OAI21X1_595 ( );
FILL FILL_0_OAI21X1_596 ( );
FILL FILL_1_OAI21X1_596 ( );
FILL FILL_0_OAI22X1_2 ( );
FILL FILL_1_OAI22X1_2 ( );
FILL FILL_2_OAI22X1_2 ( );
FILL FILL_0_OR2X2_15 ( );
FILL FILL_1_OR2X2_15 ( );
FILL FILL_0_NAND2X1_325 ( );
FILL FILL_1_NAND2X1_325 ( );
FILL FILL_0_OAI21X1_748 ( );
FILL FILL_1_OAI21X1_748 ( );
FILL FILL_0_XNOR2X1_49 ( );
FILL FILL_1_XNOR2X1_49 ( );
FILL FILL_2_XNOR2X1_49 ( );
FILL FILL_0_NAND2X1_212 ( );
FILL FILL_1_NAND2X1_212 ( );
FILL FILL_0_INVX4_17 ( );
FILL FILL_1_INVX4_17 ( );
FILL FILL_0_BUFX4_304 ( );
FILL FILL_1_BUFX4_304 ( );
FILL FILL_2_BUFX4_304 ( );
FILL FILL_0_BUFX4_285 ( );
FILL FILL_1_BUFX4_285 ( );
FILL FILL_2_BUFX4_285 ( );
FILL FILL_0_DFFPOSX1_586 ( );
FILL FILL_1_DFFPOSX1_586 ( );
FILL FILL_2_DFFPOSX1_586 ( );
FILL FILL_3_DFFPOSX1_586 ( );
FILL FILL_4_DFFPOSX1_586 ( );
FILL FILL_5_DFFPOSX1_586 ( );
FILL FILL_0_OAI21X1_716 ( );
FILL FILL_1_OAI21X1_716 ( );
FILL FILL_0_NOR2X1_106 ( );
FILL FILL_0_NAND2X1_317 ( );
FILL FILL_1_NAND2X1_317 ( );
FILL FILL_0_OR2X2_5 ( );
FILL FILL_1_OR2X2_5 ( );
FILL FILL_0_BUFX4_56 ( );
FILL FILL_1_BUFX4_56 ( );
FILL FILL_0_NOR2X1_63 ( );
FILL FILL_1_NOR2X1_63 ( );
FILL FILL_0_DFFPOSX1_295 ( );
FILL FILL_1_DFFPOSX1_295 ( );
FILL FILL_2_DFFPOSX1_295 ( );
FILL FILL_3_DFFPOSX1_295 ( );
FILL FILL_4_DFFPOSX1_295 ( );
FILL FILL_5_DFFPOSX1_295 ( );
FILL FILL_6_DFFPOSX1_295 ( );
FILL FILL_0_NAND2X1_288 ( );
FILL FILL_1_NAND2X1_288 ( );
FILL FILL_0_NAND2X1_287 ( );
FILL FILL_0_NOR2X1_74 ( );
FILL FILL_1_NOR2X1_74 ( );
FILL FILL_0_OR2X2_6 ( );
FILL FILL_1_OR2X2_6 ( );
FILL FILL_0_OAI21X1_582 ( );
FILL FILL_1_OAI21X1_582 ( );
FILL FILL_2_OAI21X1_582 ( );
FILL FILL_0_NAND3X1_17 ( );
FILL FILL_1_NAND3X1_17 ( );
FILL FILL_0_NAND3X1_16 ( );
FILL FILL_1_NAND3X1_16 ( );
FILL FILL_0_NOR2X1_72 ( );
FILL FILL_0_OAI21X1_580 ( );
FILL FILL_1_OAI21X1_580 ( );
FILL FILL_0_NAND2X1_285 ( );
FILL FILL_0_AOI21X1_7 ( );
FILL FILL_1_AOI21X1_7 ( );
FILL FILL_2_AOI21X1_7 ( );
FILL FILL_0_BUFX2_545 ( );
FILL FILL_0_XNOR2X1_33 ( );
FILL FILL_1_XNOR2X1_33 ( );
FILL FILL_2_XNOR2X1_33 ( );
FILL FILL_3_XNOR2X1_33 ( );
FILL FILL_0_BUFX4_130 ( );
FILL FILL_1_BUFX4_130 ( );
FILL FILL_0_BUFX4_133 ( );
FILL FILL_1_BUFX4_133 ( );
FILL FILL_0_DFFPOSX1_513 ( );
FILL FILL_1_DFFPOSX1_513 ( );
FILL FILL_2_DFFPOSX1_513 ( );
FILL FILL_3_DFFPOSX1_513 ( );
FILL FILL_4_DFFPOSX1_513 ( );
FILL FILL_5_DFFPOSX1_513 ( );
FILL FILL_0_BUFX4_79 ( );
FILL FILL_1_BUFX4_79 ( );
FILL FILL_2_BUFX4_79 ( );
FILL FILL_0_BUFX4_31 ( );
FILL FILL_1_BUFX4_31 ( );
FILL FILL_0_OAI21X1_212 ( );
FILL FILL_1_OAI21X1_212 ( );
FILL FILL_0_BUFX4_27 ( );
FILL FILL_1_BUFX4_27 ( );
FILL FILL_2_BUFX4_27 ( );
FILL FILL_0_NAND2X1_421 ( );
FILL FILL_1_NAND2X1_421 ( );
FILL FILL_0_CLKBUF1_83 ( );
FILL FILL_1_CLKBUF1_83 ( );
FILL FILL_2_CLKBUF1_83 ( );
FILL FILL_3_CLKBUF1_83 ( );
FILL FILL_4_CLKBUF1_83 ( );
FILL FILL_0_DFFPOSX1_769 ( );
FILL FILL_1_DFFPOSX1_769 ( );
FILL FILL_2_DFFPOSX1_769 ( );
FILL FILL_3_DFFPOSX1_769 ( );
FILL FILL_4_DFFPOSX1_769 ( );
FILL FILL_5_DFFPOSX1_769 ( );
FILL FILL_0_NAND2X1_427 ( );
FILL FILL_0_OAI21X1_1061 ( );
FILL FILL_1_OAI21X1_1061 ( );
FILL FILL_0_BUFX4_86 ( );
FILL FILL_1_BUFX4_86 ( );
FILL FILL_0_BUFX4_371 ( );
FILL FILL_1_BUFX4_371 ( );
FILL FILL_0_OAI21X1_1279 ( );
FILL FILL_1_OAI21X1_1279 ( );
FILL FILL_0_AND2X2_27 ( );
FILL FILL_1_AND2X2_27 ( );
FILL FILL_0_DFFPOSX1_891 ( );
FILL FILL_1_DFFPOSX1_891 ( );
FILL FILL_2_DFFPOSX1_891 ( );
FILL FILL_3_DFFPOSX1_891 ( );
FILL FILL_4_DFFPOSX1_891 ( );
FILL FILL_5_DFFPOSX1_891 ( );
FILL FILL_6_DFFPOSX1_891 ( );
FILL FILL_0_OAI21X1_1280 ( );
FILL FILL_1_OAI21X1_1280 ( );
FILL FILL_0_DFFPOSX1_897 ( );
FILL FILL_1_DFFPOSX1_897 ( );
FILL FILL_2_DFFPOSX1_897 ( );
FILL FILL_3_DFFPOSX1_897 ( );
FILL FILL_4_DFFPOSX1_897 ( );
FILL FILL_5_DFFPOSX1_897 ( );
FILL FILL_6_DFFPOSX1_897 ( );
FILL FILL_0_DFFPOSX1_1003 ( );
FILL FILL_1_DFFPOSX1_1003 ( );
FILL FILL_2_DFFPOSX1_1003 ( );
FILL FILL_3_DFFPOSX1_1003 ( );
FILL FILL_4_DFFPOSX1_1003 ( );
FILL FILL_5_DFFPOSX1_1003 ( );
FILL FILL_0_OAI21X1_236 ( );
FILL FILL_1_OAI21X1_236 ( );
FILL FILL_0_DFFPOSX1_310 ( );
FILL FILL_1_DFFPOSX1_310 ( );
FILL FILL_2_DFFPOSX1_310 ( );
FILL FILL_3_DFFPOSX1_310 ( );
FILL FILL_4_DFFPOSX1_310 ( );
FILL FILL_5_DFFPOSX1_310 ( );
FILL FILL_6_DFFPOSX1_310 ( );
FILL FILL_0_OAI21X1_1673 ( );
FILL FILL_1_OAI21X1_1673 ( );
FILL FILL_2_OAI21X1_1673 ( );
FILL FILL_0_OAI21X1_1070 ( );
FILL FILL_1_OAI21X1_1070 ( );
FILL FILL_2_OAI21X1_1070 ( );
FILL FILL_0_OAI21X1_1627 ( );
FILL FILL_1_OAI21X1_1627 ( );
FILL FILL_0_NAND2X1_695 ( );
FILL FILL_0_BUFX4_267 ( );
FILL FILL_1_BUFX4_267 ( );
FILL FILL_2_BUFX4_267 ( );
FILL FILL_0_NOR2X1_197 ( );
FILL FILL_1_NOR2X1_197 ( );
FILL FILL_0_NOR3X1_17 ( );
FILL FILL_1_NOR3X1_17 ( );
FILL FILL_2_NOR3X1_17 ( );
FILL FILL_3_NOR3X1_17 ( );
FILL FILL_4_NOR3X1_17 ( );
FILL FILL_0_BUFX4_308 ( );
FILL FILL_1_BUFX4_308 ( );
FILL FILL_0_BUFX2_215 ( );
FILL FILL_0_DFFPOSX1_970 ( );
FILL FILL_1_DFFPOSX1_970 ( );
FILL FILL_2_DFFPOSX1_970 ( );
FILL FILL_3_DFFPOSX1_970 ( );
FILL FILL_4_DFFPOSX1_970 ( );
FILL FILL_5_DFFPOSX1_970 ( );
FILL FILL_0_OAI21X1_1323 ( );
FILL FILL_1_OAI21X1_1323 ( );
FILL FILL_0_NOR2X1_202 ( );
FILL FILL_0_OAI21X1_1169 ( );
FILL FILL_1_OAI21X1_1169 ( );
FILL FILL_0_OAI21X1_1168 ( );
FILL FILL_1_OAI21X1_1168 ( );
FILL FILL_2_OAI21X1_1168 ( );
FILL FILL_0_OAI21X1_1324 ( );
FILL FILL_1_OAI21X1_1324 ( );
FILL FILL_2_OAI21X1_1324 ( );
FILL FILL_0_INVX1_209 ( );
FILL FILL_0_OAI21X1_1347 ( );
FILL FILL_1_OAI21X1_1347 ( );
FILL FILL_0_DFFPOSX1_922 ( );
FILL FILL_1_DFFPOSX1_922 ( );
FILL FILL_2_DFFPOSX1_922 ( );
FILL FILL_3_DFFPOSX1_922 ( );
FILL FILL_4_DFFPOSX1_922 ( );
FILL FILL_5_DFFPOSX1_922 ( );
FILL FILL_0_DFFPOSX1_786 ( );
FILL FILL_1_DFFPOSX1_786 ( );
FILL FILL_2_DFFPOSX1_786 ( );
FILL FILL_3_DFFPOSX1_786 ( );
FILL FILL_4_DFFPOSX1_786 ( );
FILL FILL_5_DFFPOSX1_786 ( );
FILL FILL_0_NAND3X1_51 ( );
FILL FILL_1_NAND3X1_51 ( );
FILL FILL_0_BUFX4_99 ( );
FILL FILL_1_BUFX4_99 ( );
FILL FILL_0_NOR2X1_211 ( );
FILL FILL_1_NOR2X1_211 ( );
FILL FILL_0_BUFX4_96 ( );
FILL FILL_1_BUFX4_96 ( );
FILL FILL_0_OAI21X1_1514 ( );
FILL FILL_1_OAI21X1_1514 ( );
FILL FILL_2_OAI21X1_1514 ( );
FILL FILL_0_DFFPOSX1_979 ( );
FILL FILL_1_DFFPOSX1_979 ( );
FILL FILL_2_DFFPOSX1_979 ( );
FILL FILL_3_DFFPOSX1_979 ( );
FILL FILL_4_DFFPOSX1_979 ( );
FILL FILL_5_DFFPOSX1_979 ( );
FILL FILL_0_INVX2_89 ( );
FILL FILL_0_NAND3X1_61 ( );
FILL FILL_1_NAND3X1_61 ( );
FILL FILL_0_INVX1_199 ( );
FILL FILL_0_OAI21X1_1200 ( );
FILL FILL_1_OAI21X1_1200 ( );
FILL FILL_0_OAI21X1_1201 ( );
FILL FILL_1_OAI21X1_1201 ( );
FILL FILL_0_INVX1_217 ( );
FILL FILL_0_NOR2X1_212 ( );
FILL FILL_1_NOR2X1_212 ( );
FILL FILL_0_OAI21X1_1198 ( );
FILL FILL_1_OAI21X1_1198 ( );
FILL FILL_0_OAI21X1_1199 ( );
FILL FILL_1_OAI21X1_1199 ( );
FILL FILL_0_NOR2X1_175 ( );
FILL FILL_1_NOR2X1_175 ( );
FILL FILL_0_INVX1_181 ( );
FILL FILL_0_AOI21X1_58 ( );
FILL FILL_1_AOI21X1_58 ( );
FILL FILL_0_OAI21X1_1563 ( );
FILL FILL_1_OAI21X1_1563 ( );
FILL FILL_0_XNOR2X1_88 ( );
FILL FILL_1_XNOR2X1_88 ( );
FILL FILL_2_XNOR2X1_88 ( );
FILL FILL_0_BUFX4_1 ( );
FILL FILL_1_BUFX4_1 ( );
FILL FILL_2_BUFX4_1 ( );
FILL FILL_0_BUFX2_38 ( );
FILL FILL_0_OAI21X1_1373 ( );
FILL FILL_1_OAI21X1_1373 ( );
FILL FILL_2_OAI21X1_1373 ( );
FILL FILL_0_OAI21X1_1372 ( );
FILL FILL_1_OAI21X1_1372 ( );
FILL FILL_0_DFFPOSX1_931 ( );
FILL FILL_1_DFFPOSX1_931 ( );
FILL FILL_2_DFFPOSX1_931 ( );
FILL FILL_3_DFFPOSX1_931 ( );
FILL FILL_4_DFFPOSX1_931 ( );
FILL FILL_5_DFFPOSX1_931 ( );
FILL FILL_0_BUFX2_184 ( );
FILL FILL_1_BUFX2_184 ( );
FILL FILL_0_OAI21X1_938 ( );
FILL FILL_1_OAI21X1_938 ( );
FILL FILL_2_OAI21X1_938 ( );
FILL FILL_0_OAI21X1_939 ( );
FILL FILL_1_OAI21X1_939 ( );
FILL FILL_0_DFFPOSX1_695 ( );
FILL FILL_1_DFFPOSX1_695 ( );
FILL FILL_2_DFFPOSX1_695 ( );
FILL FILL_3_DFFPOSX1_695 ( );
FILL FILL_4_DFFPOSX1_695 ( );
FILL FILL_5_DFFPOSX1_695 ( );
FILL FILL_0_DFFPOSX1_617 ( );
FILL FILL_1_DFFPOSX1_617 ( );
FILL FILL_2_DFFPOSX1_617 ( );
FILL FILL_3_DFFPOSX1_617 ( );
FILL FILL_4_DFFPOSX1_617 ( );
FILL FILL_5_DFFPOSX1_617 ( );
FILL FILL_0_BUFX2_739 ( );
FILL FILL_1_BUFX2_739 ( );
FILL FILL_0_NAND2X1_686 ( );
FILL FILL_1_NAND2X1_686 ( );
FILL FILL_0_OAI21X1_1618 ( );
FILL FILL_1_OAI21X1_1618 ( );
FILL FILL_0_DFFPOSX1_8 ( );
FILL FILL_1_DFFPOSX1_8 ( );
FILL FILL_2_DFFPOSX1_8 ( );
FILL FILL_3_DFFPOSX1_8 ( );
FILL FILL_4_DFFPOSX1_8 ( );
FILL FILL_5_DFFPOSX1_8 ( );
FILL FILL_0_OAI21X1_1719 ( );
FILL FILL_1_OAI21X1_1719 ( );
FILL FILL_0_DFFPOSX1_72 ( );
FILL FILL_1_DFFPOSX1_72 ( );
FILL FILL_2_DFFPOSX1_72 ( );
FILL FILL_3_DFFPOSX1_72 ( );
FILL FILL_4_DFFPOSX1_72 ( );
FILL FILL_5_DFFPOSX1_72 ( );
FILL FILL_6_DFFPOSX1_72 ( );
FILL FILL_0_BUFX2_394 ( );
FILL FILL_0_BUFX2_724 ( );
FILL FILL_0_BUFX2_393 ( );
FILL FILL_1_BUFX2_393 ( );
FILL FILL_0_DFFPOSX1_356 ( );
FILL FILL_1_DFFPOSX1_356 ( );
FILL FILL_2_DFFPOSX1_356 ( );
FILL FILL_3_DFFPOSX1_356 ( );
FILL FILL_4_DFFPOSX1_356 ( );
FILL FILL_5_DFFPOSX1_356 ( );
FILL FILL_6_DFFPOSX1_356 ( );
FILL FILL_0_NAND2X1_72 ( );
FILL FILL_0_OAI21X1_328 ( );
FILL FILL_1_OAI21X1_328 ( );
FILL FILL_0_NAND2X1_73 ( );
FILL FILL_1_NAND2X1_73 ( );
FILL FILL_0_OAI21X1_329 ( );
FILL FILL_1_OAI21X1_329 ( );
FILL FILL_0_INVX4_1 ( );
FILL FILL_1_INVX4_1 ( );
FILL FILL_0_DFFPOSX1_484 ( );
FILL FILL_1_DFFPOSX1_484 ( );
FILL FILL_2_DFFPOSX1_484 ( );
FILL FILL_3_DFFPOSX1_484 ( );
FILL FILL_4_DFFPOSX1_484 ( );
FILL FILL_5_DFFPOSX1_484 ( );
FILL FILL_6_DFFPOSX1_484 ( );
FILL FILL_0_OAI21X1_501 ( );
FILL FILL_1_OAI21X1_501 ( );
FILL FILL_0_OAI21X1_500 ( );
FILL FILL_1_OAI21X1_500 ( );
FILL FILL_0_BUFX4_302 ( );
FILL FILL_1_BUFX4_302 ( );
FILL FILL_0_CLKBUF1_80 ( );
FILL FILL_1_CLKBUF1_80 ( );
FILL FILL_2_CLKBUF1_80 ( );
FILL FILL_3_CLKBUF1_80 ( );
FILL FILL_4_CLKBUF1_80 ( );
FILL FILL_0_CLKBUF1_84 ( );
FILL FILL_1_CLKBUF1_84 ( );
FILL FILL_2_CLKBUF1_84 ( );
FILL FILL_3_CLKBUF1_84 ( );
FILL FILL_4_CLKBUF1_84 ( );
FILL FILL_0_BUFX4_90 ( );
FILL FILL_1_BUFX4_90 ( );
FILL FILL_0_BUFX4_254 ( );
FILL FILL_1_BUFX4_254 ( );
FILL FILL_2_BUFX4_254 ( );
FILL FILL_0_DFFPOSX1_528 ( );
FILL FILL_1_DFFPOSX1_528 ( );
FILL FILL_2_DFFPOSX1_528 ( );
FILL FILL_3_DFFPOSX1_528 ( );
FILL FILL_4_DFFPOSX1_528 ( );
FILL FILL_5_DFFPOSX1_528 ( );
FILL FILL_0_OAI21X1_614 ( );
FILL FILL_1_OAI21X1_614 ( );
FILL FILL_2_OAI21X1_614 ( );
FILL FILL_0_NOR2X1_85 ( );
FILL FILL_1_NOR2X1_85 ( );
FILL FILL_0_AOI21X1_14 ( );
FILL FILL_1_AOI21X1_14 ( );
FILL FILL_2_AOI21X1_14 ( );
FILL FILL_0_NAND2X1_222 ( );
FILL FILL_1_NAND2X1_222 ( );
FILL FILL_0_OAI21X1_463 ( );
FILL FILL_1_OAI21X1_463 ( );
FILL FILL_0_NOR2X1_37 ( );
FILL FILL_0_INVX4_21 ( );
FILL FILL_1_INVX4_21 ( );
FILL FILL_0_AND2X2_15 ( );
FILL FILL_1_AND2X2_15 ( );
FILL FILL_0_INVX1_32 ( );
FILL FILL_0_OAI21X1_613 ( );
FILL FILL_1_OAI21X1_613 ( );
FILL FILL_0_NOR2X1_36 ( );
FILL FILL_1_NOR2X1_36 ( );
FILL FILL_0_INVX2_28 ( );
FILL FILL_0_OAI21X1_775 ( );
FILL FILL_1_OAI21X1_775 ( );
FILL FILL_0_OAI21X1_784 ( );
FILL FILL_1_OAI21X1_784 ( );
FILL FILL_0_NOR2X1_38 ( );
FILL FILL_0_INVX2_44 ( );
FILL FILL_0_OAI21X1_779 ( );
FILL FILL_1_OAI21X1_779 ( );
FILL FILL_0_OAI21X1_780 ( );
FILL FILL_1_OAI21X1_780 ( );
FILL FILL_0_OAI21X1_793 ( );
FILL FILL_1_OAI21X1_793 ( );
FILL FILL_0_OAI21X1_794 ( );
FILL FILL_1_OAI21X1_794 ( );
FILL FILL_0_OAI21X1_797 ( );
FILL FILL_1_OAI21X1_797 ( );
FILL FILL_0_NAND2X1_231 ( );
FILL FILL_0_NAND3X1_7 ( );
FILL FILL_1_NAND3X1_7 ( );
FILL FILL_0_NAND3X1_30 ( );
FILL FILL_1_NAND3X1_30 ( );
FILL FILL_0_NAND3X1_32 ( );
FILL FILL_1_NAND3X1_32 ( );
FILL FILL_0_NOR2X1_42 ( );
FILL FILL_0_NAND3X1_10 ( );
FILL FILL_1_NAND3X1_10 ( );
FILL FILL_0_OAI21X1_639 ( );
FILL FILL_1_OAI21X1_639 ( );
FILL FILL_0_NAND2X1_300 ( );
FILL FILL_0_INVX1_21 ( );
FILL FILL_1_INVX1_21 ( );
FILL FILL_0_NAND3X1_24 ( );
FILL FILL_1_NAND3X1_24 ( );
FILL FILL_0_NAND2X1_301 ( );
FILL FILL_1_NAND2X1_301 ( );
FILL FILL_0_OAI21X1_770 ( );
FILL FILL_1_OAI21X1_770 ( );
FILL FILL_0_NAND2X1_328 ( );
FILL FILL_1_NAND2X1_328 ( );
FILL FILL_0_NOR2X1_84 ( );
FILL FILL_1_NOR2X1_84 ( );
FILL FILL_0_NAND2X1_289 ( );
FILL FILL_1_NAND2X1_289 ( );
FILL FILL_0_AND2X2_7 ( );
FILL FILL_1_AND2X2_7 ( );
FILL FILL_2_AND2X2_7 ( );
FILL FILL_0_NAND2X1_232 ( );
FILL FILL_0_BUFX2_611 ( );
FILL FILL_1_BUFX2_611 ( );
FILL FILL_0_INVX4_18 ( );
FILL FILL_1_INVX4_18 ( );
FILL FILL_0_NOR2X1_34 ( );
FILL FILL_0_NAND2X1_216 ( );
FILL FILL_1_NAND2X1_216 ( );
FILL FILL_0_OAI21X1_750 ( );
FILL FILL_1_OAI21X1_750 ( );
FILL FILL_0_NAND3X1_6 ( );
FILL FILL_1_NAND3X1_6 ( );
FILL FILL_2_NAND3X1_6 ( );
FILL FILL_0_OAI21X1_761 ( );
FILL FILL_1_OAI21X1_761 ( );
FILL FILL_0_OAI21X1_760 ( );
FILL FILL_1_OAI21X1_760 ( );
FILL FILL_0_CLKBUF1_9 ( );
FILL FILL_1_CLKBUF1_9 ( );
FILL FILL_2_CLKBUF1_9 ( );
FILL FILL_3_CLKBUF1_9 ( );
FILL FILL_4_CLKBUF1_9 ( );
FILL FILL_0_NAND3X1_29 ( );
FILL FILL_1_NAND3X1_29 ( );
FILL FILL_2_NAND3X1_29 ( );
FILL FILL_0_INVX1_41 ( );
FILL FILL_0_OAI21X1_757 ( );
FILL FILL_1_OAI21X1_757 ( );
FILL FILL_0_DFFPOSX1_582 ( );
FILL FILL_1_DFFPOSX1_582 ( );
FILL FILL_2_DFFPOSX1_582 ( );
FILL FILL_3_DFFPOSX1_582 ( );
FILL FILL_4_DFFPOSX1_582 ( );
FILL FILL_5_DFFPOSX1_582 ( );
FILL FILL_0_BUFX4_300 ( );
FILL FILL_1_BUFX4_300 ( );
FILL FILL_0_OAI21X1_713 ( );
FILL FILL_1_OAI21X1_713 ( );
FILL FILL_0_INVX1_37 ( );
FILL FILL_0_OAI21X1_712 ( );
FILL FILL_1_OAI21X1_712 ( );
FILL FILL_0_OAI21X1_709 ( );
FILL FILL_1_OAI21X1_709 ( );
FILL FILL_0_BUFX2_547 ( );
FILL FILL_0_OAI21X1_554 ( );
FILL FILL_1_OAI21X1_554 ( );
FILL FILL_0_OAI21X1_553 ( );
FILL FILL_1_OAI21X1_553 ( );
FILL FILL_2_OAI21X1_553 ( );
FILL FILL_0_BUFX2_445 ( );
FILL FILL_1_BUFX2_445 ( );
FILL FILL_0_BUFX4_271 ( );
FILL FILL_1_BUFX4_271 ( );
FILL FILL_0_NAND2X1_279 ( );
FILL FILL_1_NAND2X1_279 ( );
FILL FILL_0_NOR2X1_76 ( );
FILL FILL_0_AOI21X1_8 ( );
FILL FILL_1_AOI21X1_8 ( );
FILL FILL_2_AOI21X1_8 ( );
FILL FILL_0_OR2X2_7 ( );
FILL FILL_1_OR2X2_7 ( );
FILL FILL_0_BUFX4_287 ( );
FILL FILL_1_BUFX4_287 ( );
FILL FILL_0_NAND2X1_286 ( );
FILL FILL_0_XNOR2X1_12 ( );
FILL FILL_1_XNOR2X1_12 ( );
FILL FILL_2_XNOR2X1_12 ( );
FILL FILL_0_CLKBUF1_63 ( );
FILL FILL_1_CLKBUF1_63 ( );
FILL FILL_2_CLKBUF1_63 ( );
FILL FILL_3_CLKBUF1_63 ( );
FILL FILL_4_CLKBUF1_63 ( );
FILL FILL_0_OAI21X1_581 ( );
FILL FILL_1_OAI21X1_581 ( );
FILL FILL_0_DFFPOSX1_514 ( );
FILL FILL_1_DFFPOSX1_514 ( );
FILL FILL_2_DFFPOSX1_514 ( );
FILL FILL_3_DFFPOSX1_514 ( );
FILL FILL_4_DFFPOSX1_514 ( );
FILL FILL_5_DFFPOSX1_514 ( );
FILL FILL_6_DFFPOSX1_514 ( );
FILL FILL_0_OAI21X1_578 ( );
FILL FILL_1_OAI21X1_578 ( );
FILL FILL_0_OAI21X1_579 ( );
FILL FILL_1_OAI21X1_579 ( );
FILL FILL_0_DFFPOSX1_763 ( );
FILL FILL_1_DFFPOSX1_763 ( );
FILL FILL_2_DFFPOSX1_763 ( );
FILL FILL_3_DFFPOSX1_763 ( );
FILL FILL_4_DFFPOSX1_763 ( );
FILL FILL_5_DFFPOSX1_763 ( );
FILL FILL_6_DFFPOSX1_763 ( );
FILL FILL_0_DFFPOSX1_298 ( );
FILL FILL_1_DFFPOSX1_298 ( );
FILL FILL_2_DFFPOSX1_298 ( );
FILL FILL_3_DFFPOSX1_298 ( );
FILL FILL_4_DFFPOSX1_298 ( );
FILL FILL_5_DFFPOSX1_298 ( );
FILL FILL_0_OAI21X1_213 ( );
FILL FILL_1_OAI21X1_213 ( );
FILL FILL_0_OAI21X1_1055 ( );
FILL FILL_1_OAI21X1_1055 ( );
FILL FILL_0_NOR2X1_221 ( );
FILL FILL_1_NOR2X1_221 ( );
FILL FILL_0_NOR2X1_137 ( );
FILL FILL_0_INVX1_188 ( );
FILL FILL_0_DFFPOSX1_960 ( );
FILL FILL_1_DFFPOSX1_960 ( );
FILL FILL_2_DFFPOSX1_960 ( );
FILL FILL_3_DFFPOSX1_960 ( );
FILL FILL_4_DFFPOSX1_960 ( );
FILL FILL_5_DFFPOSX1_960 ( );
FILL FILL_6_DFFPOSX1_960 ( );
FILL FILL_0_BUFX4_113 ( );
FILL FILL_1_BUFX4_113 ( );
FILL FILL_0_XNOR2X1_78 ( );
FILL FILL_1_XNOR2X1_78 ( );
FILL FILL_2_XNOR2X1_78 ( );
FILL FILL_3_XNOR2X1_78 ( );
FILL FILL_0_OAI21X1_1263 ( );
FILL FILL_1_OAI21X1_1263 ( );
FILL FILL_0_OAI21X1_1262 ( );
FILL FILL_1_OAI21X1_1262 ( );
FILL FILL_0_OAI21X1_1577 ( );
FILL FILL_1_OAI21X1_1577 ( );
FILL FILL_0_OAI21X1_1578 ( );
FILL FILL_1_OAI21X1_1578 ( );
FILL FILL_0_DFFPOSX1_1002 ( );
FILL FILL_1_DFFPOSX1_1002 ( );
FILL FILL_2_DFFPOSX1_1002 ( );
FILL FILL_3_DFFPOSX1_1002 ( );
FILL FILL_4_DFFPOSX1_1002 ( );
FILL FILL_5_DFFPOSX1_1002 ( );
FILL FILL_0_DFFPOSX1_778 ( );
FILL FILL_1_DFFPOSX1_778 ( );
FILL FILL_2_DFFPOSX1_778 ( );
FILL FILL_3_DFFPOSX1_778 ( );
FILL FILL_4_DFFPOSX1_778 ( );
FILL FILL_5_DFFPOSX1_778 ( );
FILL FILL_6_DFFPOSX1_778 ( );
FILL FILL_0_OAI21X1_1325 ( );
FILL FILL_1_OAI21X1_1325 ( );
FILL FILL_0_DFFPOSX1_17 ( );
FILL FILL_1_DFFPOSX1_17 ( );
FILL FILL_2_DFFPOSX1_17 ( );
FILL FILL_3_DFFPOSX1_17 ( );
FILL FILL_4_DFFPOSX1_17 ( );
FILL FILL_5_DFFPOSX1_17 ( );
FILL FILL_0_OAI21X1_237 ( );
FILL FILL_1_OAI21X1_237 ( );
FILL FILL_0_XNOR2X1_100 ( );
FILL FILL_1_XNOR2X1_100 ( );
FILL FILL_2_XNOR2X1_100 ( );
FILL FILL_3_XNOR2X1_100 ( );
FILL FILL_0_OAI21X1_1672 ( );
FILL FILL_1_OAI21X1_1672 ( );
FILL FILL_0_OAI21X1_1484 ( );
FILL FILL_1_OAI21X1_1484 ( );
FILL FILL_0_NAND2X1_533 ( );
FILL FILL_0_AND2X2_23 ( );
FILL FILL_1_AND2X2_23 ( );
FILL FILL_0_OAI21X1_1346 ( );
FILL FILL_1_OAI21X1_1346 ( );
FILL FILL_0_NOR3X1_18 ( );
FILL FILL_1_NOR3X1_18 ( );
FILL FILL_2_NOR3X1_18 ( );
FILL FILL_3_NOR3X1_18 ( );
FILL FILL_0_NOR2X1_160 ( );
FILL FILL_1_NOR2X1_160 ( );
FILL FILL_0_OAI21X1_1511 ( );
FILL FILL_1_OAI21X1_1511 ( );
FILL FILL_0_DFFPOSX1_978 ( );
FILL FILL_1_DFFPOSX1_978 ( );
FILL FILL_2_DFFPOSX1_978 ( );
FILL FILL_3_DFFPOSX1_978 ( );
FILL FILL_4_DFFPOSX1_978 ( );
FILL FILL_5_DFFPOSX1_978 ( );
FILL FILL_6_DFFPOSX1_978 ( );
FILL FILL_0_NAND2X1_549 ( );
FILL FILL_0_INVX2_80 ( );
FILL FILL_0_INVX1_194 ( );
FILL FILL_0_BUFX4_258 ( );
FILL FILL_1_BUFX4_258 ( );
FILL FILL_0_DFFPOSX1_914 ( );
FILL FILL_1_DFFPOSX1_914 ( );
FILL FILL_2_DFFPOSX1_914 ( );
FILL FILL_3_DFFPOSX1_914 ( );
FILL FILL_4_DFFPOSX1_914 ( );
FILL FILL_5_DFFPOSX1_914 ( );
FILL FILL_0_OAI21X1_1078 ( );
FILL FILL_1_OAI21X1_1078 ( );
FILL FILL_0_NAND2X1_444 ( );
FILL FILL_1_NAND2X1_444 ( );
FILL FILL_0_NAND2X1_565 ( );
FILL FILL_1_NAND2X1_565 ( );
FILL FILL_0_AND2X2_24 ( );
FILL FILL_1_AND2X2_24 ( );
FILL FILL_0_NAND3X1_50 ( );
FILL FILL_1_NAND3X1_50 ( );
FILL FILL_2_NAND3X1_50 ( );
FILL FILL_0_INVX1_198 ( );
FILL FILL_0_OAI21X1_1558 ( );
FILL FILL_1_OAI21X1_1558 ( );
FILL FILL_0_NAND2X1_646 ( );
FILL FILL_1_NAND2X1_646 ( );
FILL FILL_0_OR2X2_21 ( );
FILL FILL_1_OR2X2_21 ( );
FILL FILL_0_NOR2X1_231 ( );
FILL FILL_0_NAND2X1_645 ( );
FILL FILL_1_NAND2X1_645 ( );
FILL FILL_0_NAND3X1_62 ( );
FILL FILL_1_NAND3X1_62 ( );
FILL FILL_0_NOR2X1_214 ( );
FILL FILL_1_NOR2X1_214 ( );
FILL FILL_0_INVX2_112 ( );
FILL FILL_0_INVX1_218 ( );
FILL FILL_0_NOR2X1_213 ( );
FILL FILL_1_NOR2X1_213 ( );
FILL FILL_0_INVX2_91 ( );
FILL FILL_0_NOR2X1_176 ( );
FILL FILL_0_NAND2X1_586 ( );
FILL FILL_1_NAND2X1_586 ( );
FILL FILL_0_OAI21X1_1565 ( );
FILL FILL_1_OAI21X1_1565 ( );
FILL FILL_0_BUFX4_105 ( );
FILL FILL_1_BUFX4_105 ( );
FILL FILL_2_BUFX4_105 ( );
FILL FILL_0_BUFX2_230 ( );
FILL FILL_0_NOR2X1_174 ( );
FILL FILL_1_NOR2X1_174 ( );
FILL FILL_0_AOI21X1_44 ( );
FILL FILL_1_AOI21X1_44 ( );
FILL FILL_0_OAI21X1_1562 ( );
FILL FILL_1_OAI21X1_1562 ( );
FILL FILL_0_INVX2_90 ( );
FILL FILL_0_AOI21X1_65 ( );
FILL FILL_1_AOI21X1_65 ( );
FILL FILL_0_NOR2X1_232 ( );
FILL FILL_1_NOR2X1_232 ( );
FILL FILL_0_OAI21X1_1566 ( );
FILL FILL_1_OAI21X1_1566 ( );
FILL FILL_2_OAI21X1_1566 ( );
FILL FILL_0_DFFPOSX1_996 ( );
FILL FILL_1_DFFPOSX1_996 ( );
FILL FILL_2_DFFPOSX1_996 ( );
FILL FILL_3_DFFPOSX1_996 ( );
FILL FILL_4_DFFPOSX1_996 ( );
FILL FILL_5_DFFPOSX1_996 ( );
FILL FILL_0_BUFX4_111 ( );
FILL FILL_1_BUFX4_111 ( );
FILL FILL_2_BUFX4_111 ( );
FILL FILL_0_OAI21X1_1564 ( );
FILL FILL_1_OAI21X1_1564 ( );
FILL FILL_0_BUFX2_250 ( );
FILL FILL_1_BUFX2_250 ( );
FILL FILL_0_OAI21X1_170 ( );
FILL FILL_1_OAI21X1_170 ( );
FILL FILL_0_OAI21X1_171 ( );
FILL FILL_1_OAI21X1_171 ( );
FILL FILL_0_DFFPOSX1_277 ( );
FILL FILL_1_DFFPOSX1_277 ( );
FILL FILL_2_DFFPOSX1_277 ( );
FILL FILL_3_DFFPOSX1_277 ( );
FILL FILL_4_DFFPOSX1_277 ( );
FILL FILL_5_DFFPOSX1_277 ( );
FILL FILL_0_OAI21X1_922 ( );
FILL FILL_1_OAI21X1_922 ( );
FILL FILL_0_OAI21X1_923 ( );
FILL FILL_1_OAI21X1_923 ( );
FILL FILL_2_OAI21X1_923 ( );
FILL FILL_0_INVX1_116 ( );
FILL FILL_0_BUFX2_354 ( );
FILL FILL_1_BUFX2_354 ( );
FILL FILL_0_INVX1_80 ( );
FILL FILL_0_BUFX2_340 ( );
FILL FILL_1_BUFX2_340 ( );
FILL FILL_0_BUFX2_316 ( );
FILL FILL_0_BUFX2_892 ( );
FILL FILL_1_BUFX2_892 ( );
FILL FILL_0_BUFX2_828 ( );
FILL FILL_0_DFFPOSX1_219 ( );
FILL FILL_1_DFFPOSX1_219 ( );
FILL FILL_2_DFFPOSX1_219 ( );
FILL FILL_3_DFFPOSX1_219 ( );
FILL FILL_4_DFFPOSX1_219 ( );
FILL FILL_5_DFFPOSX1_219 ( );
FILL FILL_6_DFFPOSX1_219 ( );
FILL FILL_0_NAND2X1_63 ( );
FILL FILL_0_OAI21X1_63 ( );
FILL FILL_1_OAI21X1_63 ( );
FILL FILL_0_NAND2X1_770 ( );
FILL FILL_1_NAND2X1_770 ( );
FILL FILL_0_OAI21X1_1829 ( );
FILL FILL_1_OAI21X1_1829 ( );
FILL FILL_0_OAI21X1_1654 ( );
FILL FILL_1_OAI21X1_1654 ( );
FILL FILL_0_OAI21X1_1655 ( );
FILL FILL_1_OAI21X1_1655 ( );
FILL FILL_0_DFFPOSX1_40 ( );
FILL FILL_1_DFFPOSX1_40 ( );
FILL FILL_2_DFFPOSX1_40 ( );
FILL FILL_3_DFFPOSX1_40 ( );
FILL FILL_4_DFFPOSX1_40 ( );
FILL FILL_5_DFFPOSX1_40 ( );
FILL FILL_0_BUFX4_367 ( );
FILL FILL_1_BUFX4_367 ( );
FILL FILL_0_BUFX2_749 ( );
FILL FILL_1_BUFX2_749 ( );
FILL FILL_0_CLKBUF1_87 ( );
FILL FILL_1_CLKBUF1_87 ( );
FILL FILL_2_CLKBUF1_87 ( );
FILL FILL_3_CLKBUF1_87 ( );
FILL FILL_4_CLKBUF1_87 ( );
FILL FILL_0_BUFX2_660 ( );
FILL FILL_1_BUFX2_660 ( );
FILL FILL_0_BUFX4_321 ( );
FILL FILL_1_BUFX4_321 ( );
FILL FILL_0_DFFPOSX1_357 ( );
FILL FILL_1_DFFPOSX1_357 ( );
FILL FILL_2_DFFPOSX1_357 ( );
FILL FILL_3_DFFPOSX1_357 ( );
FILL FILL_4_DFFPOSX1_357 ( );
FILL FILL_5_DFFPOSX1_357 ( );
FILL FILL_0_NAND2X1_669 ( );
FILL FILL_1_NAND2X1_669 ( );
FILL FILL_0_OAI21X1_1600 ( );
FILL FILL_1_OAI21X1_1600 ( );
FILL FILL_0_DFFPOSX1_55 ( );
FILL FILL_1_DFFPOSX1_55 ( );
FILL FILL_2_DFFPOSX1_55 ( );
FILL FILL_3_DFFPOSX1_55 ( );
FILL FILL_4_DFFPOSX1_55 ( );
FILL FILL_5_DFFPOSX1_55 ( );
FILL FILL_6_DFFPOSX1_55 ( );
FILL FILL_0_OAI21X1_1685 ( );
FILL FILL_1_OAI21X1_1685 ( );
FILL FILL_0_OAI21X1_1684 ( );
FILL FILL_1_OAI21X1_1684 ( );
FILL FILL_0_BUFX2_429 ( );
FILL FILL_1_BUFX2_429 ( );
FILL FILL_0_BUFX4_362 ( );
FILL FILL_1_BUFX4_362 ( );
FILL FILL_0_NAND2X1_113 ( );
FILL FILL_0_OAI21X1_369 ( );
FILL FILL_1_OAI21X1_369 ( );
FILL FILL_0_BUFX2_559 ( );
FILL FILL_1_BUFX2_559 ( );
FILL FILL_0_BUFX2_430 ( );
FILL FILL_0_BUFX4_274 ( );
FILL FILL_1_BUFX4_274 ( );
FILL FILL_2_BUFX4_274 ( );
FILL FILL_0_BUFX2_493 ( );
FILL FILL_0_OAI21X1_612 ( );
FILL FILL_1_OAI21X1_612 ( );
FILL FILL_0_DFFPOSX1_461 ( );
FILL FILL_1_DFFPOSX1_461 ( );
FILL FILL_2_DFFPOSX1_461 ( );
FILL FILL_3_DFFPOSX1_461 ( );
FILL FILL_4_DFFPOSX1_461 ( );
FILL FILL_5_DFFPOSX1_461 ( );
FILL FILL_0_NAND2X1_220 ( );
FILL FILL_0_OAI21X1_461 ( );
FILL FILL_1_OAI21X1_461 ( );
FILL FILL_0_NAND2X1_224 ( );
FILL FILL_0_XNOR2X1_36 ( );
FILL FILL_1_XNOR2X1_36 ( );
FILL FILL_2_XNOR2X1_36 ( );
FILL FILL_3_XNOR2X1_36 ( );
FILL FILL_0_AOI21X1_13 ( );
FILL FILL_1_AOI21X1_13 ( );
FILL FILL_0_NAND2X1_296 ( );
FILL FILL_0_NAND2X1_114 ( );
FILL FILL_1_NAND2X1_114 ( );
FILL FILL_0_INVX4_20 ( );
FILL FILL_1_INVX4_20 ( );
FILL FILL_0_NAND2X1_219 ( );
FILL FILL_1_NAND2X1_219 ( );
FILL FILL_0_NAND2X1_218 ( );
FILL FILL_1_NAND2X1_218 ( );
FILL FILL_0_OAI21X1_460 ( );
FILL FILL_1_OAI21X1_460 ( );
FILL FILL_0_NOR2X1_35 ( );
FILL FILL_0_OAI21X1_459 ( );
FILL FILL_1_OAI21X1_459 ( );
FILL FILL_0_NAND2X1_217 ( );
FILL FILL_0_DFFPOSX1_460 ( );
FILL FILL_1_DFFPOSX1_460 ( );
FILL FILL_2_DFFPOSX1_460 ( );
FILL FILL_3_DFFPOSX1_460 ( );
FILL FILL_4_DFFPOSX1_460 ( );
FILL FILL_5_DFFPOSX1_460 ( );
FILL FILL_6_DFFPOSX1_460 ( );
FILL FILL_0_DFFPOSX1_409 ( );
FILL FILL_1_DFFPOSX1_409 ( );
FILL FILL_2_DFFPOSX1_409 ( );
FILL FILL_3_DFFPOSX1_409 ( );
FILL FILL_4_DFFPOSX1_409 ( );
FILL FILL_5_DFFPOSX1_409 ( );
FILL FILL_0_NAND2X1_125 ( );
FILL FILL_0_OAI21X1_381 ( );
FILL FILL_1_OAI21X1_381 ( );
FILL FILL_2_OAI21X1_381 ( );
FILL FILL_0_INVX4_19 ( );
FILL FILL_0_NOR2X1_47 ( );
FILL FILL_1_NOR2X1_47 ( );
FILL FILL_0_NOR3X1_8 ( );
FILL FILL_1_NOR3X1_8 ( );
FILL FILL_2_NOR3X1_8 ( );
FILL FILL_3_NOR3X1_8 ( );
FILL FILL_0_NAND2X1_302 ( );
FILL FILL_1_NAND2X1_302 ( );
FILL FILL_0_DFFPOSX1_540 ( );
FILL FILL_1_DFFPOSX1_540 ( );
FILL FILL_2_DFFPOSX1_540 ( );
FILL FILL_3_DFFPOSX1_540 ( );
FILL FILL_4_DFFPOSX1_540 ( );
FILL FILL_5_DFFPOSX1_540 ( );
FILL FILL_6_DFFPOSX1_540 ( );
FILL FILL_0_NAND2X1_255 ( );
FILL FILL_1_NAND2X1_255 ( );
FILL FILL_0_BUFX4_61 ( );
FILL FILL_1_BUFX4_61 ( );
FILL FILL_0_BUFX4_155 ( );
FILL FILL_1_BUFX4_155 ( );
FILL FILL_0_BUFX4_33 ( );
FILL FILL_1_BUFX4_33 ( );
FILL FILL_2_BUFX4_33 ( );
FILL FILL_0_BUFX4_346 ( );
FILL FILL_1_BUFX4_346 ( );
FILL FILL_0_OAI21X1_749 ( );
FILL FILL_1_OAI21X1_749 ( );
FILL FILL_0_DFFPOSX1_580 ( );
FILL FILL_1_DFFPOSX1_580 ( );
FILL FILL_2_DFFPOSX1_580 ( );
FILL FILL_3_DFFPOSX1_580 ( );
FILL FILL_4_DFFPOSX1_580 ( );
FILL FILL_5_DFFPOSX1_580 ( );
FILL FILL_0_BUFX4_299 ( );
FILL FILL_1_BUFX4_299 ( );
FILL FILL_0_BUFX4_306 ( );
FILL FILL_1_BUFX4_306 ( );
FILL FILL_0_INVX2_27 ( );
FILL FILL_0_XNOR2X1_51 ( );
FILL FILL_1_XNOR2X1_51 ( );
FILL FILL_2_XNOR2X1_51 ( );
FILL FILL_0_NAND2X1_327 ( );
FILL FILL_1_NAND2X1_327 ( );
FILL FILL_0_NOR2X1_112 ( );
FILL FILL_1_NOR2X1_112 ( );
FILL FILL_0_NOR2X1_32 ( );
FILL FILL_1_NOR2X1_32 ( );
FILL FILL_0_BUFX4_288 ( );
FILL FILL_1_BUFX4_288 ( );
FILL FILL_0_BUFX4_142 ( );
FILL FILL_1_BUFX4_142 ( );
FILL FILL_0_OAI21X1_756 ( );
FILL FILL_1_OAI21X1_756 ( );
FILL FILL_2_OAI21X1_756 ( );
FILL FILL_0_NOR2X1_111 ( );
FILL FILL_0_XNOR2X1_50 ( );
FILL FILL_1_XNOR2X1_50 ( );
FILL FILL_2_XNOR2X1_50 ( );
FILL FILL_3_XNOR2X1_50 ( );
FILL FILL_0_BUFX4_119 ( );
FILL FILL_1_BUFX4_119 ( );
FILL FILL_0_OAI21X1_711 ( );
FILL FILL_1_OAI21X1_711 ( );
FILL FILL_0_BUFX4_54 ( );
FILL FILL_1_BUFX4_54 ( );
FILL FILL_0_BUFX4_71 ( );
FILL FILL_1_BUFX4_71 ( );
FILL FILL_0_INVX8_6 ( );
FILL FILL_1_INVX8_6 ( );
FILL FILL_0_BUFX4_41 ( );
FILL FILL_1_BUFX4_41 ( );
FILL FILL_0_NOR2X1_73 ( );
FILL FILL_0_AOI21X1_9 ( );
FILL FILL_1_AOI21X1_9 ( );
FILL FILL_0_DFFPOSX1_512 ( );
FILL FILL_1_DFFPOSX1_512 ( );
FILL FILL_2_DFFPOSX1_512 ( );
FILL FILL_3_DFFPOSX1_512 ( );
FILL FILL_4_DFFPOSX1_512 ( );
FILL FILL_5_DFFPOSX1_512 ( );
FILL FILL_6_DFFPOSX1_512 ( );
FILL FILL_0_OAI21X1_576 ( );
FILL FILL_1_OAI21X1_576 ( );
FILL FILL_2_OAI21X1_576 ( );
FILL FILL_0_BUFX4_309 ( );
FILL FILL_1_BUFX4_309 ( );
FILL FILL_0_BUFX4_266 ( );
FILL FILL_1_BUFX4_266 ( );
FILL FILL_0_BUFX4_260 ( );
FILL FILL_1_BUFX4_260 ( );
FILL FILL_0_CLKBUF1_60 ( );
FILL FILL_1_CLKBUF1_60 ( );
FILL FILL_2_CLKBUF1_60 ( );
FILL FILL_3_CLKBUF1_60 ( );
FILL FILL_4_CLKBUF1_60 ( );
FILL FILL_0_OAI21X1_577 ( );
FILL FILL_1_OAI21X1_577 ( );
FILL FILL_0_BUFX4_378 ( );
FILL FILL_1_BUFX4_378 ( );
FILL FILL_0_OAI21X1_1441 ( );
FILL FILL_1_OAI21X1_1441 ( );
FILL FILL_0_OAI21X1_1442 ( );
FILL FILL_1_OAI21X1_1442 ( );
FILL FILL_0_OAI21X1_1440 ( );
FILL FILL_1_OAI21X1_1440 ( );
FILL FILL_2_OAI21X1_1440 ( );
FILL FILL_0_OAI21X1_1439 ( );
FILL FILL_1_OAI21X1_1439 ( );
FILL FILL_0_NOR2X1_136 ( );
FILL FILL_1_NOR2X1_136 ( );
FILL FILL_0_INVX2_97 ( );
FILL FILL_0_BUFX4_174 ( );
FILL FILL_1_BUFX4_174 ( );
FILL FILL_0_NAND2X1_630 ( );
FILL FILL_1_NAND2X1_630 ( );
FILL FILL_0_OAI21X1_1455 ( );
FILL FILL_1_OAI21X1_1455 ( );
FILL FILL_0_OAI21X1_1454 ( );
FILL FILL_1_OAI21X1_1454 ( );
FILL FILL_0_NAND2X1_513 ( );
FILL FILL_0_NAND2X1_602 ( );
FILL FILL_1_NAND2X1_602 ( );
FILL FILL_0_BUFX4_298 ( );
FILL FILL_1_BUFX4_298 ( );
FILL FILL_2_BUFX4_298 ( );
FILL FILL_0_OAI21X1_1717 ( );
FILL FILL_1_OAI21X1_1717 ( );
FILL FILL_0_INVX8_2 ( );
FILL FILL_1_INVX8_2 ( );
FILL FILL_2_INVX8_2 ( );
FILL FILL_0_OAI21X1_1716 ( );
FILL FILL_1_OAI21X1_1716 ( );
FILL FILL_2_OAI21X1_1716 ( );
FILL FILL_0_BUFX4_129 ( );
FILL FILL_1_BUFX4_129 ( );
FILL FILL_0_OAI21X1_93 ( );
FILL FILL_1_OAI21X1_93 ( );
FILL FILL_0_BUFX4_157 ( );
FILL FILL_1_BUFX4_157 ( );
FILL FILL_2_BUFX4_157 ( );
FILL FILL_0_OAI21X1_92 ( );
FILL FILL_1_OAI21X1_92 ( );
FILL FILL_0_BUFX4_5 ( );
FILL FILL_1_BUFX4_5 ( );
FILL FILL_0_BUFX4_160 ( );
FILL FILL_1_BUFX4_160 ( );
FILL FILL_0_BUFX4_284 ( );
FILL FILL_1_BUFX4_284 ( );
FILL FILL_0_NAND2X1_635 ( );
FILL FILL_0_NAND2X1_616 ( );
FILL FILL_1_NAND2X1_616 ( );
FILL FILL_0_OAI21X1_1327 ( );
FILL FILL_1_OAI21X1_1327 ( );
FILL FILL_0_BUFX4_297 ( );
FILL FILL_1_BUFX4_297 ( );
FILL FILL_0_AND2X2_33 ( );
FILL FILL_1_AND2X2_33 ( );
FILL FILL_0_NAND3X1_59 ( );
FILL FILL_1_NAND3X1_59 ( );
FILL FILL_0_NAND2X1_620 ( );
FILL FILL_1_NAND2X1_620 ( );
FILL FILL_0_INVX2_107 ( );
FILL FILL_0_NAND2X1_615 ( );
FILL FILL_0_OAI21X1_1510 ( );
FILL FILL_1_OAI21X1_1510 ( );
FILL FILL_2_OAI21X1_1510 ( );
FILL FILL_0_NAND2X1_639 ( );
FILL FILL_0_OAI21X1_1512 ( );
FILL FILL_1_OAI21X1_1512 ( );
FILL FILL_2_OAI21X1_1512 ( );
FILL FILL_0_XNOR2X1_102 ( );
FILL FILL_1_XNOR2X1_102 ( );
FILL FILL_2_XNOR2X1_102 ( );
FILL FILL_0_NAND3X1_67 ( );
FILL FILL_1_NAND3X1_67 ( );
FILL FILL_0_NOR2X1_166 ( );
FILL FILL_0_NAND2X1_556 ( );
FILL FILL_1_NAND2X1_556 ( );
FILL FILL_0_INVX1_213 ( );
FILL FILL_0_NOR2X1_206 ( );
FILL FILL_1_NOR2X1_206 ( );
FILL FILL_0_AOI21X1_54 ( );
FILL FILL_1_AOI21X1_54 ( );
FILL FILL_0_NAND2X1_619 ( );
FILL FILL_0_BUFX4_243 ( );
FILL FILL_1_BUFX4_243 ( );
FILL FILL_0_OAI21X1_1344 ( );
FILL FILL_1_OAI21X1_1344 ( );
FILL FILL_2_OAI21X1_1344 ( );
FILL FILL_0_OAI21X1_1342 ( );
FILL FILL_1_OAI21X1_1342 ( );
FILL FILL_0_OAI21X1_1559 ( );
FILL FILL_1_OAI21X1_1559 ( );
FILL FILL_0_OAI21X1_1560 ( );
FILL FILL_1_OAI21X1_1560 ( );
FILL FILL_0_DFFPOSX1_994 ( );
FILL FILL_1_DFFPOSX1_994 ( );
FILL FILL_2_DFFPOSX1_994 ( );
FILL FILL_3_DFFPOSX1_994 ( );
FILL FILL_4_DFFPOSX1_994 ( );
FILL FILL_5_DFFPOSX1_994 ( );
FILL FILL_0_BUFX2_247 ( );
FILL FILL_1_BUFX2_247 ( );
FILL FILL_0_OAI21X1_1567 ( );
FILL FILL_1_OAI21X1_1567 ( );
FILL FILL_0_OAI21X1_1570 ( );
FILL FILL_1_OAI21X1_1570 ( );
FILL FILL_2_OAI21X1_1570 ( );
FILL FILL_0_OAI21X1_1197 ( );
FILL FILL_1_OAI21X1_1197 ( );
FILL FILL_0_AOI21X1_45 ( );
FILL FILL_1_AOI21X1_45 ( );
FILL FILL_0_AOI21X1_66 ( );
FILL FILL_1_AOI21X1_66 ( );
FILL FILL_0_OAI21X1_1202 ( );
FILL FILL_1_OAI21X1_1202 ( );
FILL FILL_0_OAI21X1_1203 ( );
FILL FILL_1_OAI21X1_1203 ( );
FILL FILL_0_NAND2X1_585 ( );
FILL FILL_1_NAND2X1_585 ( );
FILL FILL_0_NOR2X1_173 ( );
FILL FILL_0_DFFPOSX1_869 ( );
FILL FILL_1_DFFPOSX1_869 ( );
FILL FILL_2_DFFPOSX1_869 ( );
FILL FILL_3_DFFPOSX1_869 ( );
FILL FILL_4_DFFPOSX1_869 ( );
FILL FILL_5_DFFPOSX1_869 ( );
FILL FILL_6_DFFPOSX1_869 ( );
FILL FILL_0_AOI21X1_59 ( );
FILL FILL_1_AOI21X1_59 ( );
FILL FILL_0_OAI21X1_1205 ( );
FILL FILL_1_OAI21X1_1205 ( );
FILL FILL_0_NAND2X1_587 ( );
FILL FILL_1_NAND2X1_587 ( );
FILL FILL_0_DFFPOSX1_870 ( );
FILL FILL_1_DFFPOSX1_870 ( );
FILL FILL_2_DFFPOSX1_870 ( );
FILL FILL_3_DFFPOSX1_870 ( );
FILL FILL_4_DFFPOSX1_870 ( );
FILL FILL_5_DFFPOSX1_870 ( );
FILL FILL_0_BUFX2_124 ( );
FILL FILL_0_OAI21X1_1206 ( );
FILL FILL_1_OAI21X1_1206 ( );
FILL FILL_0_AND2X2_25 ( );
FILL FILL_1_AND2X2_25 ( );
FILL FILL_0_OAI21X1_1207 ( );
FILL FILL_1_OAI21X1_1207 ( );
FILL FILL_0_NAND2X1_589 ( );
FILL FILL_1_NAND2X1_589 ( );
FILL FILL_0_DFFPOSX1_871 ( );
FILL FILL_1_DFFPOSX1_871 ( );
FILL FILL_2_DFFPOSX1_871 ( );
FILL FILL_3_DFFPOSX1_871 ( );
FILL FILL_4_DFFPOSX1_871 ( );
FILL FILL_5_DFFPOSX1_871 ( );
FILL FILL_6_DFFPOSX1_871 ( );
FILL FILL_0_BUFX2_55 ( );
FILL FILL_1_BUFX2_55 ( );
FILL FILL_0_BUFX2_123 ( );
FILL FILL_1_BUFX2_123 ( );
FILL FILL_0_BUFX2_125 ( );
FILL FILL_1_BUFX2_125 ( );
FILL FILL_0_BUFX2_173 ( );
FILL FILL_0_DFFPOSX1_687 ( );
FILL FILL_1_DFFPOSX1_687 ( );
FILL FILL_2_DFFPOSX1_687 ( );
FILL FILL_3_DFFPOSX1_687 ( );
FILL FILL_4_DFFPOSX1_687 ( );
FILL FILL_5_DFFPOSX1_687 ( );
FILL FILL_6_DFFPOSX1_687 ( );
FILL FILL_0_BUFX2_683 ( );
FILL FILL_0_DFFPOSX1_661 ( );
FILL FILL_1_DFFPOSX1_661 ( );
FILL FILL_2_DFFPOSX1_661 ( );
FILL FILL_3_DFFPOSX1_661 ( );
FILL FILL_4_DFFPOSX1_661 ( );
FILL FILL_5_DFFPOSX1_661 ( );
FILL FILL_6_DFFPOSX1_661 ( );
FILL FILL_0_BUFX2_187 ( );
FILL FILL_1_BUFX2_187 ( );
FILL FILL_0_BUFX2_382 ( );
FILL FILL_1_BUFX2_382 ( );
FILL FILL_0_BUFX2_349 ( );
FILL FILL_1_BUFX2_349 ( );
FILL FILL_0_DFFPOSX1_651 ( );
FILL FILL_1_DFFPOSX1_651 ( );
FILL FILL_2_DFFPOSX1_651 ( );
FILL FILL_3_DFFPOSX1_651 ( );
FILL FILL_4_DFFPOSX1_651 ( );
FILL FILL_5_DFFPOSX1_651 ( );
FILL FILL_0_BUFX2_297 ( );
FILL FILL_1_BUFX2_297 ( );
FILL FILL_0_BUFX2_671 ( );
FILL FILL_1_BUFX2_671 ( );
FILL FILL_0_OAI21X1_870 ( );
FILL FILL_1_OAI21X1_870 ( );
FILL FILL_0_BUFX2_708 ( );
FILL FILL_1_BUFX2_708 ( );
FILL FILL_0_BUFX2_280 ( );
FILL FILL_0_INVX2_129 ( );
FILL FILL_0_BUFX2_685 ( );
FILL FILL_0_DFFPOSX1_16 ( );
FILL FILL_1_DFFPOSX1_16 ( );
FILL FILL_2_DFFPOSX1_16 ( );
FILL FILL_3_DFFPOSX1_16 ( );
FILL FILL_4_DFFPOSX1_16 ( );
FILL FILL_5_DFFPOSX1_16 ( );
FILL FILL_6_DFFPOSX1_16 ( );
FILL FILL_0_NAND2X1_694 ( );
FILL FILL_0_OAI21X1_1626 ( );
FILL FILL_1_OAI21X1_1626 ( );
FILL FILL_0_DFFPOSX1_155 ( );
FILL FILL_1_DFFPOSX1_155 ( );
FILL FILL_2_DFFPOSX1_155 ( );
FILL FILL_3_DFFPOSX1_155 ( );
FILL FILL_4_DFFPOSX1_155 ( );
FILL FILL_5_DFFPOSX1_155 ( );
FILL FILL_0_BUFX2_717 ( );
FILL FILL_1_BUFX2_717 ( );
FILL FILL_0_DFFPOSX1_48 ( );
FILL FILL_1_DFFPOSX1_48 ( );
FILL FILL_2_DFFPOSX1_48 ( );
FILL FILL_3_DFFPOSX1_48 ( );
FILL FILL_4_DFFPOSX1_48 ( );
FILL FILL_5_DFFPOSX1_48 ( );
FILL FILL_6_DFFPOSX1_48 ( );
FILL FILL_0_OAI21X1_1671 ( );
FILL FILL_1_OAI21X1_1671 ( );
FILL FILL_0_OAI21X1_1735 ( );
FILL FILL_1_OAI21X1_1735 ( );
FILL FILL_0_OAI21X1_1734 ( );
FILL FILL_1_OAI21X1_1734 ( );
FILL FILL_0_DFFPOSX1_80 ( );
FILL FILL_1_DFFPOSX1_80 ( );
FILL FILL_2_DFFPOSX1_80 ( );
FILL FILL_3_DFFPOSX1_80 ( );
FILL FILL_4_DFFPOSX1_80 ( );
FILL FILL_5_DFFPOSX1_80 ( );
FILL FILL_0_CLKBUF1_45 ( );
FILL FILL_1_CLKBUF1_45 ( );
FILL FILL_2_CLKBUF1_45 ( );
FILL FILL_3_CLKBUF1_45 ( );
FILL FILL_4_CLKBUF1_45 ( );
FILL FILL_0_DFFPOSX1_1023 ( );
FILL FILL_1_DFFPOSX1_1023 ( );
FILL FILL_2_DFFPOSX1_1023 ( );
FILL FILL_3_DFFPOSX1_1023 ( );
FILL FILL_4_DFFPOSX1_1023 ( );
FILL FILL_5_DFFPOSX1_1023 ( );
FILL FILL_6_DFFPOSX1_1023 ( );
FILL FILL_0_BUFX2_624 ( );
FILL FILL_1_BUFX2_624 ( );
FILL FILL_0_OAI21X1_669 ( );
FILL FILL_1_OAI21X1_669 ( );
FILL FILL_2_OAI21X1_669 ( );
FILL FILL_0_OAI21X1_668 ( );
FILL FILL_1_OAI21X1_668 ( );
FILL FILL_0_BUFX4_72 ( );
FILL FILL_1_BUFX4_72 ( );
FILL FILL_2_BUFX4_72 ( );
FILL FILL_0_BUFX4_52 ( );
FILL FILL_1_BUFX4_52 ( );
FILL FILL_0_DFFPOSX1_397 ( );
FILL FILL_1_DFFPOSX1_397 ( );
FILL FILL_2_DFFPOSX1_397 ( );
FILL FILL_3_DFFPOSX1_397 ( );
FILL FILL_4_DFFPOSX1_397 ( );
FILL FILL_5_DFFPOSX1_397 ( );
FILL FILL_6_DFFPOSX1_397 ( );
FILL FILL_0_DFFPOSX1_527 ( );
FILL FILL_1_DFFPOSX1_527 ( );
FILL FILL_2_DFFPOSX1_527 ( );
FILL FILL_3_DFFPOSX1_527 ( );
FILL FILL_4_DFFPOSX1_527 ( );
FILL FILL_5_DFFPOSX1_527 ( );
FILL FILL_6_DFFPOSX1_527 ( );
FILL FILL_0_OAI21X1_609 ( );
FILL FILL_1_OAI21X1_609 ( );
FILL FILL_0_OAI21X1_611 ( );
FILL FILL_1_OAI21X1_611 ( );
FILL FILL_0_XNOR2X1_37 ( );
FILL FILL_1_XNOR2X1_37 ( );
FILL FILL_2_XNOR2X1_37 ( );
FILL FILL_3_XNOR2X1_37 ( );
FILL FILL_0_XNOR2X1_19 ( );
FILL FILL_1_XNOR2X1_19 ( );
FILL FILL_2_XNOR2X1_19 ( );
FILL FILL_3_XNOR2X1_19 ( );
FILL FILL_0_OAI21X1_610 ( );
FILL FILL_1_OAI21X1_610 ( );
FILL FILL_0_DFFPOSX1_398 ( );
FILL FILL_1_DFFPOSX1_398 ( );
FILL FILL_2_DFFPOSX1_398 ( );
FILL FILL_3_DFFPOSX1_398 ( );
FILL FILL_4_DFFPOSX1_398 ( );
FILL FILL_5_DFFPOSX1_398 ( );
FILL FILL_0_OAI21X1_370 ( );
FILL FILL_1_OAI21X1_370 ( );
FILL FILL_0_OAI21X1_462 ( );
FILL FILL_1_OAI21X1_462 ( );
FILL FILL_0_BUFX4_256 ( );
FILL FILL_1_BUFX4_256 ( );
FILL FILL_0_INVX4_23 ( );
FILL FILL_1_INVX4_23 ( );
FILL FILL_0_INVX1_17 ( );
FILL FILL_0_OAI21X1_458 ( );
FILL FILL_1_OAI21X1_458 ( );
FILL FILL_2_OAI21X1_458 ( );
FILL FILL_0_XNOR2X1_53 ( );
FILL FILL_1_XNOR2X1_53 ( );
FILL FILL_2_XNOR2X1_53 ( );
FILL FILL_3_XNOR2X1_53 ( );
FILL FILL_0_INVX2_53 ( );
FILL FILL_0_NOR2X1_115 ( );
FILL FILL_1_NOR2X1_115 ( );
FILL FILL_0_BUFX4_116 ( );
FILL FILL_1_BUFX4_116 ( );
FILL FILL_0_OAI21X1_640 ( );
FILL FILL_1_OAI21X1_640 ( );
FILL FILL_2_OAI21X1_640 ( );
FILL FILL_0_AOI21X1_21 ( );
FILL FILL_1_AOI21X1_21 ( );
FILL FILL_0_NAND3X1_25 ( );
FILL FILL_1_NAND3X1_25 ( );
FILL FILL_2_NAND3X1_25 ( );
FILL FILL_0_OR2X2_12 ( );
FILL FILL_1_OR2X2_12 ( );
FILL FILL_0_AOI21X1_22 ( );
FILL FILL_1_AOI21X1_22 ( );
FILL FILL_0_AOI21X1_23 ( );
FILL FILL_1_AOI21X1_23 ( );
FILL FILL_0_NOR2X1_96 ( );
FILL FILL_0_DFFPOSX1_477 ( );
FILL FILL_1_DFFPOSX1_477 ( );
FILL FILL_2_DFFPOSX1_477 ( );
FILL FILL_3_DFFPOSX1_477 ( );
FILL FILL_4_DFFPOSX1_477 ( );
FILL FILL_5_DFFPOSX1_477 ( );
FILL FILL_6_DFFPOSX1_477 ( );
FILL FILL_0_DFFPOSX1_476 ( );
FILL FILL_1_DFFPOSX1_476 ( );
FILL FILL_2_DFFPOSX1_476 ( );
FILL FILL_3_DFFPOSX1_476 ( );
FILL FILL_4_DFFPOSX1_476 ( );
FILL FILL_5_DFFPOSX1_476 ( );
FILL FILL_0_DFFPOSX1_611 ( );
FILL FILL_1_DFFPOSX1_611 ( );
FILL FILL_2_DFFPOSX1_611 ( );
FILL FILL_3_DFFPOSX1_611 ( );
FILL FILL_4_DFFPOSX1_611 ( );
FILL FILL_5_DFFPOSX1_611 ( );
FILL FILL_6_DFFPOSX1_611 ( );
FILL FILL_0_OAI21X1_843 ( );
FILL FILL_1_OAI21X1_843 ( );
FILL FILL_0_OAI21X1_841 ( );
FILL FILL_1_OAI21X1_841 ( );
FILL FILL_0_NAND2X1_259 ( );
FILL FILL_0_DFFPOSX1_587 ( );
FILL FILL_1_DFFPOSX1_587 ( );
FILL FILL_2_DFFPOSX1_587 ( );
FILL FILL_3_DFFPOSX1_587 ( );
FILL FILL_4_DFFPOSX1_587 ( );
FILL FILL_5_DFFPOSX1_587 ( );
FILL FILL_0_NOR2X1_33 ( );
FILL FILL_0_OAI21X1_768 ( );
FILL FILL_1_OAI21X1_768 ( );
FILL FILL_2_OAI21X1_768 ( );
FILL FILL_0_OAI21X1_769 ( );
FILL FILL_1_OAI21X1_769 ( );
FILL FILL_0_INVX8_4 ( );
FILL FILL_1_INVX8_4 ( );
FILL FILL_2_INVX8_4 ( );
FILL FILL_0_XNOR2X1_16 ( );
FILL FILL_1_XNOR2X1_16 ( );
FILL FILL_2_XNOR2X1_16 ( );
FILL FILL_0_DFFPOSX1_503 ( );
FILL FILL_1_DFFPOSX1_503 ( );
FILL FILL_2_DFFPOSX1_503 ( );
FILL FILL_3_DFFPOSX1_503 ( );
FILL FILL_4_DFFPOSX1_503 ( );
FILL FILL_5_DFFPOSX1_503 ( );
FILL FILL_6_DFFPOSX1_503 ( );
FILL FILL_0_OAI21X1_555 ( );
FILL FILL_1_OAI21X1_555 ( );
FILL FILL_0_OAI21X1_556 ( );
FILL FILL_1_OAI21X1_556 ( );
FILL FILL_0_OAI21X1_718 ( );
FILL FILL_1_OAI21X1_718 ( );
FILL FILL_0_BUFX4_22 ( );
FILL FILL_1_BUFX4_22 ( );
FILL FILL_0_OAI21X1_710 ( );
FILL FILL_1_OAI21X1_710 ( );
FILL FILL_0_DFFPOSX1_516 ( );
FILL FILL_1_DFFPOSX1_516 ( );
FILL FILL_2_DFFPOSX1_516 ( );
FILL FILL_3_DFFPOSX1_516 ( );
FILL FILL_4_DFFPOSX1_516 ( );
FILL FILL_5_DFFPOSX1_516 ( );
FILL FILL_6_DFFPOSX1_516 ( );
FILL FILL_0_OAI21X1_772 ( );
FILL FILL_1_OAI21X1_772 ( );
FILL FILL_0_OAI21X1_771 ( );
FILL FILL_1_OAI21X1_771 ( );
FILL FILL_0_BUFX4_175 ( );
FILL FILL_1_BUFX4_175 ( );
FILL FILL_0_INVX1_28 ( );
FILL FILL_0_OAI21X1_354 ( );
FILL FILL_1_OAI21X1_354 ( );
FILL FILL_0_OAI21X1_569 ( );
FILL FILL_1_OAI21X1_569 ( );
FILL FILL_2_OAI21X1_569 ( );
FILL FILL_0_OAI21X1_570 ( );
FILL FILL_1_OAI21X1_570 ( );
FILL FILL_0_XNOR2X1_32 ( );
FILL FILL_1_XNOR2X1_32 ( );
FILL FILL_2_XNOR2X1_32 ( );
FILL FILL_3_XNOR2X1_32 ( );
FILL FILL_0_OAI21X1_567 ( );
FILL FILL_1_OAI21X1_567 ( );
FILL FILL_0_OAI21X1_566 ( );
FILL FILL_1_OAI21X1_566 ( );
FILL FILL_0_DFFPOSX1_509 ( );
FILL FILL_1_DFFPOSX1_509 ( );
FILL FILL_2_DFFPOSX1_509 ( );
FILL FILL_3_DFFPOSX1_509 ( );
FILL FILL_4_DFFPOSX1_509 ( );
FILL FILL_5_DFFPOSX1_509 ( );
FILL FILL_0_BUFX4_19 ( );
FILL FILL_1_BUFX4_19 ( );
FILL FILL_0_DFFPOSX1_955 ( );
FILL FILL_1_DFFPOSX1_955 ( );
FILL FILL_2_DFFPOSX1_955 ( );
FILL FILL_3_DFFPOSX1_955 ( );
FILL FILL_4_DFFPOSX1_955 ( );
FILL FILL_5_DFFPOSX1_955 ( );
FILL FILL_0_BUFX4_15 ( );
FILL FILL_1_BUFX4_15 ( );
FILL FILL_0_NAND2X1_627 ( );
FILL FILL_1_NAND2X1_627 ( );
FILL FILL_0_XNOR2X1_96 ( );
FILL FILL_1_XNOR2X1_96 ( );
FILL FILL_2_XNOR2X1_96 ( );
FILL FILL_3_XNOR2X1_96 ( );
FILL FILL_0_NOR2X1_223 ( );
FILL FILL_0_NOR2X1_142 ( );
FILL FILL_1_NOR2X1_142 ( );
FILL FILL_0_NAND2X1_519 ( );
FILL FILL_0_NOR2X1_141 ( );
FILL FILL_1_NOR2X1_141 ( );
FILL FILL_0_DFFPOSX1_71 ( );
FILL FILL_1_DFFPOSX1_71 ( );
FILL FILL_2_DFFPOSX1_71 ( );
FILL FILL_3_DFFPOSX1_71 ( );
FILL FILL_4_DFFPOSX1_71 ( );
FILL FILL_5_DFFPOSX1_71 ( );
FILL FILL_0_DFFPOSX1_770 ( );
FILL FILL_1_DFFPOSX1_770 ( );
FILL FILL_2_DFFPOSX1_770 ( );
FILL FILL_3_DFFPOSX1_770 ( );
FILL FILL_4_DFFPOSX1_770 ( );
FILL FILL_5_DFFPOSX1_770 ( );
FILL FILL_6_DFFPOSX1_770 ( );
FILL FILL_0_DFFPOSX1_238 ( );
FILL FILL_1_DFFPOSX1_238 ( );
FILL FILL_2_DFFPOSX1_238 ( );
FILL FILL_3_DFFPOSX1_238 ( );
FILL FILL_4_DFFPOSX1_238 ( );
FILL FILL_5_DFFPOSX1_238 ( );
FILL FILL_0_DFFPOSX1_965 ( );
FILL FILL_1_DFFPOSX1_965 ( );
FILL FILL_2_DFFPOSX1_965 ( );
FILL FILL_3_DFFPOSX1_965 ( );
FILL FILL_4_DFFPOSX1_965 ( );
FILL FILL_5_DFFPOSX1_965 ( );
FILL FILL_6_DFFPOSX1_965 ( );
FILL FILL_0_NOR2X1_152 ( );
FILL FILL_1_NOR2X1_152 ( );
FILL FILL_0_BUFX4_307 ( );
FILL FILL_1_BUFX4_307 ( );
FILL FILL_0_DFFPOSX1_915 ( );
FILL FILL_1_DFFPOSX1_915 ( );
FILL FILL_2_DFFPOSX1_915 ( );
FILL FILL_3_DFFPOSX1_915 ( );
FILL FILL_4_DFFPOSX1_915 ( );
FILL FILL_5_DFFPOSX1_915 ( );
FILL FILL_6_DFFPOSX1_915 ( );
FILL FILL_0_BUFX4_259 ( );
FILL FILL_1_BUFX4_259 ( );
FILL FILL_0_NAND3X1_57 ( );
FILL FILL_1_NAND3X1_57 ( );
FILL FILL_0_INVX1_210 ( );
FILL FILL_0_OAI21X1_259 ( );
FILL FILL_1_OAI21X1_259 ( );
FILL FILL_2_OAI21X1_259 ( );
FILL FILL_0_BUFX4_294 ( );
FILL FILL_1_BUFX4_294 ( );
FILL FILL_0_BUFX4_59 ( );
FILL FILL_1_BUFX4_59 ( );
FILL FILL_2_BUFX4_59 ( );
FILL FILL_0_BUFX4_32 ( );
FILL FILL_1_BUFX4_32 ( );
FILL FILL_0_INVX2_110 ( );
FILL FILL_0_INVX4_43 ( );
FILL FILL_1_INVX4_43 ( );
FILL FILL_0_INVX1_224 ( );
FILL FILL_0_NAND3X1_66 ( );
FILL FILL_1_NAND3X1_66 ( );
FILL FILL_0_XNOR2X1_85 ( );
FILL FILL_1_XNOR2X1_85 ( );
FILL FILL_2_XNOR2X1_85 ( );
FILL FILL_3_XNOR2X1_85 ( );
FILL FILL_0_AND2X2_32 ( );
FILL FILL_1_AND2X2_32 ( );
FILL FILL_0_NOR2X1_207 ( );
FILL FILL_1_NOR2X1_207 ( );
FILL FILL_0_NAND2X1_564 ( );
FILL FILL_1_NAND2X1_564 ( );
FILL FILL_0_NOR2X1_165 ( );
FILL FILL_0_NAND2X1_563 ( );
FILL FILL_1_NAND2X1_563 ( );
FILL FILL_0_OAI21X1_1343 ( );
FILL FILL_1_OAI21X1_1343 ( );
FILL FILL_0_DFFPOSX1_921 ( );
FILL FILL_1_DFFPOSX1_921 ( );
FILL FILL_2_DFFPOSX1_921 ( );
FILL FILL_3_DFFPOSX1_921 ( );
FILL FILL_4_DFFPOSX1_921 ( );
FILL FILL_5_DFFPOSX1_921 ( );
FILL FILL_6_DFFPOSX1_921 ( );
FILL FILL_0_INVX2_83 ( );
FILL FILL_0_NAND3X1_58 ( );
FILL FILL_1_NAND3X1_58 ( );
FILL FILL_0_INVX1_195 ( );
FILL FILL_0_AOI21X1_41 ( );
FILL FILL_1_AOI21X1_41 ( );
FILL FILL_0_DFFPOSX1_866 ( );
FILL FILL_1_DFFPOSX1_866 ( );
FILL FILL_2_DFFPOSX1_866 ( );
FILL FILL_3_DFFPOSX1_866 ( );
FILL FILL_4_DFFPOSX1_866 ( );
FILL FILL_5_DFFPOSX1_866 ( );
FILL FILL_0_NAND2X1_582 ( );
FILL FILL_1_NAND2X1_582 ( );
FILL FILL_0_BUFX2_119 ( );
FILL FILL_1_BUFX2_119 ( );
FILL FILL_0_OAI21X1_1569 ( );
FILL FILL_1_OAI21X1_1569 ( );
FILL FILL_0_NOR3X1_15 ( );
FILL FILL_1_NOR3X1_15 ( );
FILL FILL_2_NOR3X1_15 ( );
FILL FILL_3_NOR3X1_15 ( );
FILL FILL_0_OAI21X1_1204 ( );
FILL FILL_1_OAI21X1_1204 ( );
FILL FILL_0_INVX4_49 ( );
FILL FILL_1_INVX4_49 ( );
FILL FILL_0_NAND2X1_588 ( );
FILL FILL_1_NAND2X1_588 ( );
FILL FILL_0_INVX2_92 ( );
FILL FILL_0_NAND3X1_69 ( );
FILL FILL_1_NAND3X1_69 ( );
FILL FILL_0_XNOR2X1_89 ( );
FILL FILL_1_XNOR2X1_89 ( );
FILL FILL_2_XNOR2X1_89 ( );
FILL FILL_3_XNOR2X1_89 ( );
FILL FILL_0_OAI21X1_1383 ( );
FILL FILL_1_OAI21X1_1383 ( );
FILL FILL_0_DFFPOSX1_935 ( );
FILL FILL_1_DFFPOSX1_935 ( );
FILL FILL_2_DFFPOSX1_935 ( );
FILL FILL_3_DFFPOSX1_935 ( );
FILL FILL_4_DFFPOSX1_935 ( );
FILL FILL_5_DFFPOSX1_935 ( );
FILL FILL_0_INVX4_46 ( );
FILL FILL_0_BUFX4_330 ( );
FILL FILL_1_BUFX4_330 ( );
FILL FILL_2_BUFX4_330 ( );
FILL FILL_0_OAI21X1_1094 ( );
FILL FILL_1_OAI21X1_1094 ( );
FILL FILL_0_NAND2X1_460 ( );
FILL FILL_1_NAND2X1_460 ( );
FILL FILL_0_DFFPOSX1_802 ( );
FILL FILL_1_DFFPOSX1_802 ( );
FILL FILL_2_DFFPOSX1_802 ( );
FILL FILL_3_DFFPOSX1_802 ( );
FILL FILL_4_DFFPOSX1_802 ( );
FILL FILL_5_DFFPOSX1_802 ( );
FILL FILL_6_DFFPOSX1_802 ( );
FILL FILL_0_OAI21X1_1768 ( );
FILL FILL_1_OAI21X1_1768 ( );
FILL FILL_2_OAI21X1_1768 ( );
FILL FILL_0_OAI21X1_1769 ( );
FILL FILL_1_OAI21X1_1769 ( );
FILL FILL_0_DFFPOSX1_97 ( );
FILL FILL_1_DFFPOSX1_97 ( );
FILL FILL_2_DFFPOSX1_97 ( );
FILL FILL_3_DFFPOSX1_97 ( );
FILL FILL_4_DFFPOSX1_97 ( );
FILL FILL_5_DFFPOSX1_97 ( );
FILL FILL_0_OAI21X1_976 ( );
FILL FILL_1_OAI21X1_976 ( );
FILL FILL_0_OAI21X1_977 ( );
FILL FILL_1_OAI21X1_977 ( );
FILL FILL_0_DFFPOSX1_714 ( );
FILL FILL_1_DFFPOSX1_714 ( );
FILL FILL_2_DFFPOSX1_714 ( );
FILL FILL_3_DFFPOSX1_714 ( );
FILL FILL_4_DFFPOSX1_714 ( );
FILL FILL_5_DFFPOSX1_714 ( );
FILL FILL_0_INVX1_143 ( );
FILL FILL_0_BUFX2_767 ( );
FILL FILL_1_BUFX2_767 ( );
FILL FILL_0_BUFX2_369 ( );
FILL FILL_1_BUFX2_369 ( );
FILL FILL_0_BUFX2_668 ( );
FILL FILL_1_BUFX2_668 ( );
FILL FILL_0_DFFPOSX1_743 ( );
FILL FILL_1_DFFPOSX1_743 ( );
FILL FILL_2_DFFPOSX1_743 ( );
FILL FILL_3_DFFPOSX1_743 ( );
FILL FILL_4_DFFPOSX1_743 ( );
FILL FILL_5_DFFPOSX1_743 ( );
FILL FILL_0_INVX1_89 ( );
FILL FILL_0_BUFX2_952 ( );
FILL FILL_1_BUFX2_952 ( );
FILL FILL_0_BUFX2_320 ( );
FILL FILL_1_BUFX2_320 ( );
FILL FILL_0_BUFX2_120 ( );
FILL FILL_1_BUFX2_120 ( );
FILL FILL_0_BUFX2_364 ( );
FILL FILL_1_BUFX2_364 ( );
FILL FILL_0_BUFX2_693 ( );
FILL FILL_0_BUFX2_2 ( );
FILL FILL_1_BUFX2_2 ( );
FILL FILL_0_BUFX2_806 ( );
FILL FILL_1_BUFX2_806 ( );
FILL FILL_0_BUFX2_653 ( );
FILL FILL_1_BUFX2_653 ( );
FILL FILL_0_NAND2X1_403 ( );
FILL FILL_1_NAND2X1_403 ( );
FILL FILL_0_OAI21X1_1037 ( );
FILL FILL_1_OAI21X1_1037 ( );
FILL FILL_0_DFFPOSX1_745 ( );
FILL FILL_1_DFFPOSX1_745 ( );
FILL FILL_2_DFFPOSX1_745 ( );
FILL FILL_3_DFFPOSX1_745 ( );
FILL FILL_4_DFFPOSX1_745 ( );
FILL FILL_5_DFFPOSX1_745 ( );
FILL FILL_0_DFFPOSX1_1016 ( );
FILL FILL_1_DFFPOSX1_1016 ( );
FILL FILL_2_DFFPOSX1_1016 ( );
FILL FILL_3_DFFPOSX1_1016 ( );
FILL FILL_4_DFFPOSX1_1016 ( );
FILL FILL_5_DFFPOSX1_1016 ( );
FILL FILL_0_NAND2X1_662 ( );
FILL FILL_1_NAND2X1_662 ( );
FILL FILL_0_OAI21X1_1593 ( );
FILL FILL_1_OAI21X1_1593 ( );
FILL FILL_0_OAI21X1_1670 ( );
FILL FILL_1_OAI21X1_1670 ( );
FILL FILL_0_NAND2X1_750 ( );
FILL FILL_1_NAND2X1_750 ( );
FILL FILL_0_OAI21X1_1809 ( );
FILL FILL_1_OAI21X1_1809 ( );
FILL FILL_0_DFFPOSX1_135 ( );
FILL FILL_1_DFFPOSX1_135 ( );
FILL FILL_2_DFFPOSX1_135 ( );
FILL FILL_3_DFFPOSX1_135 ( );
FILL FILL_4_DFFPOSX1_135 ( );
FILL FILL_5_DFFPOSX1_135 ( );
FILL FILL_6_DFFPOSX1_135 ( );
FILL FILL_0_DFFPOSX1_199 ( );
FILL FILL_1_DFFPOSX1_199 ( );
FILL FILL_2_DFFPOSX1_199 ( );
FILL FILL_3_DFFPOSX1_199 ( );
FILL FILL_4_DFFPOSX1_199 ( );
FILL FILL_5_DFFPOSX1_199 ( );
FILL FILL_0_NAND2X1_43 ( );
FILL FILL_1_NAND2X1_43 ( );
FILL FILL_0_OAI21X1_43 ( );
FILL FILL_1_OAI21X1_43 ( );
FILL FILL_0_BUFX4_81 ( );
FILL FILL_1_BUFX4_81 ( );
FILL FILL_0_BUFX2_495 ( );
FILL FILL_0_NAND2X1_223 ( );
FILL FILL_1_NAND2X1_223 ( );
FILL FILL_0_OAI21X1_464 ( );
FILL FILL_1_OAI21X1_464 ( );
FILL FILL_0_BUFX2_608 ( );
FILL FILL_1_BUFX2_608 ( );
FILL FILL_0_DFFPOSX1_551 ( );
FILL FILL_1_DFFPOSX1_551 ( );
FILL FILL_2_DFFPOSX1_551 ( );
FILL FILL_3_DFFPOSX1_551 ( );
FILL FILL_4_DFFPOSX1_551 ( );
FILL FILL_5_DFFPOSX1_551 ( );
FILL FILL_6_DFFPOSX1_551 ( );
FILL FILL_0_BUFX2_435 ( );
FILL FILL_1_BUFX2_435 ( );
FILL FILL_0_DFFPOSX1_403 ( );
FILL FILL_1_DFFPOSX1_403 ( );
FILL FILL_2_DFFPOSX1_403 ( );
FILL FILL_3_DFFPOSX1_403 ( );
FILL FILL_4_DFFPOSX1_403 ( );
FILL FILL_5_DFFPOSX1_403 ( );
FILL FILL_6_DFFPOSX1_403 ( );
FILL FILL_0_NAND2X1_119 ( );
FILL FILL_1_NAND2X1_119 ( );
FILL FILL_0_OAI21X1_375 ( );
FILL FILL_1_OAI21X1_375 ( );
FILL FILL_0_BUFX2_227 ( );
FILL FILL_1_BUFX2_227 ( );
FILL FILL_0_DFFPOSX1_592 ( );
FILL FILL_1_DFFPOSX1_592 ( );
FILL FILL_2_DFFPOSX1_592 ( );
FILL FILL_3_DFFPOSX1_592 ( );
FILL FILL_4_DFFPOSX1_592 ( );
FILL FILL_5_DFFPOSX1_592 ( );
FILL FILL_6_DFFPOSX1_592 ( );
FILL FILL_0_OAI21X1_785 ( );
FILL FILL_1_OAI21X1_785 ( );
FILL FILL_0_OAI21X1_786 ( );
FILL FILL_1_OAI21X1_786 ( );
FILL FILL_0_NAND2X1_297 ( );
FILL FILL_1_NAND2X1_297 ( );
FILL FILL_0_OAI21X1_1395 ( );
FILL FILL_1_OAI21X1_1395 ( );
FILL FILL_0_OAI21X1_1394 ( );
FILL FILL_1_OAI21X1_1394 ( );
FILL FILL_0_DFFPOSX1_940 ( );
FILL FILL_1_DFFPOSX1_940 ( );
FILL FILL_2_DFFPOSX1_940 ( );
FILL FILL_3_DFFPOSX1_940 ( );
FILL FILL_4_DFFPOSX1_940 ( );
FILL FILL_5_DFFPOSX1_940 ( );
FILL FILL_0_NAND2X1_115 ( );
FILL FILL_0_OAI21X1_371 ( );
FILL FILL_1_OAI21X1_371 ( );
FILL FILL_2_OAI21X1_371 ( );
FILL FILL_0_OAI21X1_474 ( );
FILL FILL_1_OAI21X1_474 ( );
FILL FILL_0_OAI21X1_1119 ( );
FILL FILL_1_OAI21X1_1119 ( );
FILL FILL_0_NAND2X1_331 ( );
FILL FILL_1_NAND2X1_331 ( );
FILL FILL_0_DFFPOSX1_817 ( );
FILL FILL_1_DFFPOSX1_817 ( );
FILL FILL_2_DFFPOSX1_817 ( );
FILL FILL_3_DFFPOSX1_817 ( );
FILL FILL_4_DFFPOSX1_817 ( );
FILL FILL_5_DFFPOSX1_817 ( );
FILL FILL_6_DFFPOSX1_817 ( );
FILL FILL_0_OAI21X1_638 ( );
FILL FILL_1_OAI21X1_638 ( );
FILL FILL_0_BUFX2_572 ( );
FILL FILL_1_BUFX2_572 ( );
FILL FILL_0_DFFPOSX1_539 ( );
FILL FILL_1_DFFPOSX1_539 ( );
FILL FILL_2_DFFPOSX1_539 ( );
FILL FILL_3_DFFPOSX1_539 ( );
FILL FILL_4_DFFPOSX1_539 ( );
FILL FILL_5_DFFPOSX1_539 ( );
FILL FILL_0_INVX4_22 ( );
FILL FILL_1_INVX4_22 ( );
FILL FILL_0_NOR2X1_95 ( );
FILL FILL_0_BUFX4_325 ( );
FILL FILL_1_BUFX4_325 ( );
FILL FILL_0_XNOR2X1_39 ( );
FILL FILL_1_XNOR2X1_39 ( );
FILL FILL_2_XNOR2X1_39 ( );
FILL FILL_3_XNOR2X1_39 ( );
FILL FILL_0_NAND3X1_11 ( );
FILL FILL_1_NAND3X1_11 ( );
FILL FILL_0_NAND3X1_33 ( );
FILL FILL_1_NAND3X1_33 ( );
FILL FILL_0_OAI21X1_489 ( );
FILL FILL_1_OAI21X1_489 ( );
FILL FILL_0_NAND2X1_251 ( );
FILL FILL_0_OAI21X1_367 ( );
FILL FILL_1_OAI21X1_367 ( );
FILL FILL_2_OAI21X1_367 ( );
FILL FILL_0_BUFX4_241 ( );
FILL FILL_1_BUFX4_241 ( );
FILL FILL_2_BUFX4_241 ( );
FILL FILL_0_XNOR2X1_18 ( );
FILL FILL_1_XNOR2X1_18 ( );
FILL FILL_2_XNOR2X1_18 ( );
FILL FILL_3_XNOR2X1_18 ( );
FILL FILL_0_OAI21X1_494 ( );
FILL FILL_1_OAI21X1_494 ( );
FILL FILL_0_NOR3X1_4 ( );
FILL FILL_1_NOR3X1_4 ( );
FILL FILL_2_NOR3X1_4 ( );
FILL FILL_3_NOR3X1_4 ( );
FILL FILL_0_NAND2X1_215 ( );
FILL FILL_0_XNOR2X1_17 ( );
FILL FILL_1_XNOR2X1_17 ( );
FILL FILL_2_XNOR2X1_17 ( );
FILL FILL_3_XNOR2X1_17 ( );
FILL FILL_0_DFFPOSX1_480 ( );
FILL FILL_1_DFFPOSX1_480 ( );
FILL FILL_2_DFFPOSX1_480 ( );
FILL FILL_3_DFFPOSX1_480 ( );
FILL FILL_4_DFFPOSX1_480 ( );
FILL FILL_5_DFFPOSX1_480 ( );
FILL FILL_0_DFFPOSX1_584 ( );
FILL FILL_1_DFFPOSX1_584 ( );
FILL FILL_2_DFFPOSX1_584 ( );
FILL FILL_3_DFFPOSX1_584 ( );
FILL FILL_4_DFFPOSX1_584 ( );
FILL FILL_5_DFFPOSX1_584 ( );
FILL FILL_0_BUFX4_17 ( );
FILL FILL_1_BUFX4_17 ( );
FILL FILL_0_OAI21X1_455 ( );
FILL FILL_1_OAI21X1_455 ( );
FILL FILL_0_NAND2X1_211 ( );
FILL FILL_1_NAND2X1_211 ( );
FILL FILL_0_DFFPOSX1_457 ( );
FILL FILL_1_DFFPOSX1_457 ( );
FILL FILL_2_DFFPOSX1_457 ( );
FILL FILL_3_DFFPOSX1_457 ( );
FILL FILL_4_DFFPOSX1_457 ( );
FILL FILL_5_DFFPOSX1_457 ( );
FILL FILL_0_DFFPOSX1_568 ( );
FILL FILL_1_DFFPOSX1_568 ( );
FILL FILL_2_DFFPOSX1_568 ( );
FILL FILL_3_DFFPOSX1_568 ( );
FILL FILL_4_DFFPOSX1_568 ( );
FILL FILL_5_DFFPOSX1_568 ( );
FILL FILL_6_DFFPOSX1_568 ( );
FILL FILL_0_DFFPOSX1_566 ( );
FILL FILL_1_DFFPOSX1_566 ( );
FILL FILL_2_DFFPOSX1_566 ( );
FILL FILL_3_DFFPOSX1_566 ( );
FILL FILL_4_DFFPOSX1_566 ( );
FILL FILL_5_DFFPOSX1_566 ( );
FILL FILL_6_DFFPOSX1_566 ( );
FILL FILL_0_DFFPOSX1_588 ( );
FILL FILL_1_DFFPOSX1_588 ( );
FILL FILL_2_DFFPOSX1_588 ( );
FILL FILL_3_DFFPOSX1_588 ( );
FILL FILL_4_DFFPOSX1_588 ( );
FILL FILL_5_DFFPOSX1_588 ( );
FILL FILL_6_DFFPOSX1_588 ( );
FILL FILL_0_DFFPOSX1_412 ( );
FILL FILL_1_DFFPOSX1_412 ( );
FILL FILL_2_DFFPOSX1_412 ( );
FILL FILL_3_DFFPOSX1_412 ( );
FILL FILL_4_DFFPOSX1_412 ( );
FILL FILL_5_DFFPOSX1_412 ( );
FILL FILL_6_DFFPOSX1_412 ( );
FILL FILL_0_BUFX4_319 ( );
FILL FILL_1_BUFX4_319 ( );
FILL FILL_0_CLKBUF1_88 ( );
FILL FILL_1_CLKBUF1_88 ( );
FILL FILL_2_CLKBUF1_88 ( );
FILL FILL_3_CLKBUF1_88 ( );
FILL FILL_0_DFFPOSX1_382 ( );
FILL FILL_1_DFFPOSX1_382 ( );
FILL FILL_2_DFFPOSX1_382 ( );
FILL FILL_3_DFFPOSX1_382 ( );
FILL FILL_4_DFFPOSX1_382 ( );
FILL FILL_5_DFFPOSX1_382 ( );
FILL FILL_6_DFFPOSX1_382 ( );
FILL FILL_0_OAI21X1_1760 ( );
FILL FILL_1_OAI21X1_1760 ( );
FILL FILL_0_OAI21X1_1761 ( );
FILL FILL_1_OAI21X1_1761 ( );
FILL FILL_0_OAI21X1_353 ( );
FILL FILL_1_OAI21X1_353 ( );
FILL FILL_0_DFFPOSX1_381 ( );
FILL FILL_1_DFFPOSX1_381 ( );
FILL FILL_2_DFFPOSX1_381 ( );
FILL FILL_3_DFFPOSX1_381 ( );
FILL FILL_4_DFFPOSX1_381 ( );
FILL FILL_5_DFFPOSX1_381 ( );
FILL FILL_0_INVX2_69 ( );
FILL FILL_0_BUFX2_539 ( );
FILL FILL_1_BUFX2_539 ( );
FILL FILL_0_BUFX4_295 ( );
FILL FILL_1_BUFX4_295 ( );
FILL FILL_0_XNOR2X1_63 ( );
FILL FILL_1_XNOR2X1_63 ( );
FILL FILL_2_XNOR2X1_63 ( );
FILL FILL_3_XNOR2X1_63 ( );
FILL FILL_0_NAND2X1_517 ( );
FILL FILL_0_NAND2X1_518 ( );
FILL FILL_1_NAND2X1_518 ( );
FILL FILL_0_INVX4_37 ( );
FILL FILL_1_INVX4_37 ( );
FILL FILL_0_NAND2X1_631 ( );
FILL FILL_1_NAND2X1_631 ( );
FILL FILL_0_OAI21X1_1062 ( );
FILL FILL_1_OAI21X1_1062 ( );
FILL FILL_0_NAND2X1_428 ( );
FILL FILL_1_NAND2X1_428 ( );
FILL FILL_0_XNOR2X1_97 ( );
FILL FILL_1_XNOR2X1_97 ( );
FILL FILL_2_XNOR2X1_97 ( );
FILL FILL_3_XNOR2X1_97 ( );
FILL FILL_0_DFFPOSX1_901 ( );
FILL FILL_1_DFFPOSX1_901 ( );
FILL FILL_2_DFFPOSX1_901 ( );
FILL FILL_3_DFFPOSX1_901 ( );
FILL FILL_4_DFFPOSX1_901 ( );
FILL FILL_5_DFFPOSX1_901 ( );
FILL FILL_0_XNOR2X1_62 ( );
FILL FILL_1_XNOR2X1_62 ( );
FILL FILL_2_XNOR2X1_62 ( );
FILL FILL_0_OAI21X1_144 ( );
FILL FILL_1_OAI21X1_144 ( );
FILL FILL_0_OAI21X1_145 ( );
FILL FILL_1_OAI21X1_145 ( );
FILL FILL_0_DFFPOSX1_264 ( );
FILL FILL_1_DFFPOSX1_264 ( );
FILL FILL_2_DFFPOSX1_264 ( );
FILL FILL_3_DFFPOSX1_264 ( );
FILL FILL_4_DFFPOSX1_264 ( );
FILL FILL_5_DFFPOSX1_264 ( );
FILL FILL_0_OAI21X1_1326 ( );
FILL FILL_1_OAI21X1_1326 ( );
FILL FILL_0_BUFX4_238 ( );
FILL FILL_1_BUFX4_238 ( );
FILL FILL_0_OAI21X1_1470 ( );
FILL FILL_1_OAI21X1_1470 ( );
FILL FILL_0_OAI21X1_258 ( );
FILL FILL_1_OAI21X1_258 ( );
FILL FILL_0_OAI21X1_1469 ( );
FILL FILL_1_OAI21X1_1469 ( );
FILL FILL_2_OAI21X1_1469 ( );
FILL FILL_0_BUFX4_278 ( );
FILL FILL_1_BUFX4_278 ( );
FILL FILL_0_BUFX4_53 ( );
FILL FILL_1_BUFX4_53 ( );
FILL FILL_2_BUFX4_53 ( );
FILL FILL_0_DFFPOSX1_106 ( );
FILL FILL_1_DFFPOSX1_106 ( );
FILL FILL_2_DFFPOSX1_106 ( );
FILL FILL_3_DFFPOSX1_106 ( );
FILL FILL_4_DFFPOSX1_106 ( );
FILL FILL_5_DFFPOSX1_106 ( );
FILL FILL_0_BUFX4_344 ( );
FILL FILL_1_BUFX4_344 ( );
FILL FILL_0_NOR2X1_163 ( );
FILL FILL_0_BUFX4_166 ( );
FILL FILL_1_BUFX4_166 ( );
FILL FILL_0_OAI21X1_1328 ( );
FILL FILL_1_OAI21X1_1328 ( );
FILL FILL_0_OAI21X1_1330 ( );
FILL FILL_1_OAI21X1_1330 ( );
FILL FILL_0_AOI21X1_52 ( );
FILL FILL_1_AOI21X1_52 ( );
FILL FILL_0_NOR2X1_203 ( );
FILL FILL_1_NOR2X1_203 ( );
FILL FILL_0_OAI21X1_1329 ( );
FILL FILL_1_OAI21X1_1329 ( );
FILL FILL_0_NAND2X1_553 ( );
FILL FILL_1_NAND2X1_553 ( );
FILL FILL_0_AOI21X1_61 ( );
FILL FILL_1_AOI21X1_61 ( );
FILL FILL_0_NOR2X1_225 ( );
FILL FILL_0_OAI21X1_1334 ( );
FILL FILL_1_OAI21X1_1334 ( );
FILL FILL_0_INVX1_211 ( );
FILL FILL_1_INVX1_211 ( );
FILL FILL_0_AOI21X1_51 ( );
FILL FILL_1_AOI21X1_51 ( );
FILL FILL_2_AOI21X1_51 ( );
FILL FILL_0_NAND2X1_618 ( );
FILL FILL_1_NAND2X1_618 ( );
FILL FILL_0_BUFX4_342 ( );
FILL FILL_1_BUFX4_342 ( );
FILL FILL_0_OAI21X1_1531 ( );
FILL FILL_1_OAI21X1_1531 ( );
FILL FILL_0_NAND2X1_642 ( );
FILL FILL_1_NAND2X1_642 ( );
FILL FILL_0_OAI21X1_1085 ( );
FILL FILL_1_OAI21X1_1085 ( );
FILL FILL_2_OAI21X1_1085 ( );
FILL FILL_0_NAND2X1_451 ( );
FILL FILL_0_DFFPOSX1_793 ( );
FILL FILL_1_DFFPOSX1_793 ( );
FILL FILL_2_DFFPOSX1_793 ( );
FILL FILL_3_DFFPOSX1_793 ( );
FILL FILL_4_DFFPOSX1_793 ( );
FILL FILL_5_DFFPOSX1_793 ( );
FILL FILL_6_DFFPOSX1_793 ( );
FILL FILL_0_OAI21X1_1568 ( );
FILL FILL_1_OAI21X1_1568 ( );
FILL FILL_0_DFFPOSX1_997 ( );
FILL FILL_1_DFFPOSX1_997 ( );
FILL FILL_2_DFFPOSX1_997 ( );
FILL FILL_3_DFFPOSX1_997 ( );
FILL FILL_4_DFFPOSX1_997 ( );
FILL FILL_5_DFFPOSX1_997 ( );
FILL FILL_6_DFFPOSX1_997 ( );
FILL FILL_0_OAI21X1_1380 ( );
FILL FILL_1_OAI21X1_1380 ( );
FILL FILL_0_NAND2X1_623 ( );
FILL FILL_1_NAND2X1_623 ( );
FILL FILL_0_OAI21X1_1382 ( );
FILL FILL_1_OAI21X1_1382 ( );
FILL FILL_0_NAND2X1_647 ( );
FILL FILL_0_BUFX2_251 ( );
FILL FILL_0_XNOR2X1_104 ( );
FILL FILL_1_XNOR2X1_104 ( );
FILL FILL_2_XNOR2X1_104 ( );
FILL FILL_3_XNOR2X1_104 ( );
FILL FILL_0_OAI21X1_1574 ( );
FILL FILL_1_OAI21X1_1574 ( );
FILL FILL_2_OAI21X1_1574 ( );
FILL FILL_0_OAI21X1_1573 ( );
FILL FILL_1_OAI21X1_1573 ( );
FILL FILL_0_DFFPOSX1_999 ( );
FILL FILL_1_DFFPOSX1_999 ( );
FILL FILL_2_DFFPOSX1_999 ( );
FILL FILL_3_DFFPOSX1_999 ( );
FILL FILL_4_DFFPOSX1_999 ( );
FILL FILL_5_DFFPOSX1_999 ( );
FILL FILL_6_DFFPOSX1_999 ( );
FILL FILL_0_BUFX4_360 ( );
FILL FILL_1_BUFX4_360 ( );
FILL FILL_0_BUFX4_348 ( );
FILL FILL_1_BUFX4_348 ( );
FILL FILL_0_OAI21X1_1095 ( );
FILL FILL_1_OAI21X1_1095 ( );
FILL FILL_0_NAND2X1_461 ( );
FILL FILL_1_NAND2X1_461 ( );
FILL FILL_0_DFFPOSX1_803 ( );
FILL FILL_1_DFFPOSX1_803 ( );
FILL FILL_2_DFFPOSX1_803 ( );
FILL FILL_3_DFFPOSX1_803 ( );
FILL FILL_4_DFFPOSX1_803 ( );
FILL FILL_5_DFFPOSX1_803 ( );
FILL FILL_0_BUFX2_253 ( );
FILL FILL_1_BUFX2_253 ( );
FILL FILL_0_DFFPOSX1_250 ( );
FILL FILL_1_DFFPOSX1_250 ( );
FILL FILL_2_DFFPOSX1_250 ( );
FILL FILL_3_DFFPOSX1_250 ( );
FILL FILL_4_DFFPOSX1_250 ( );
FILL FILL_5_DFFPOSX1_250 ( );
FILL FILL_6_DFFPOSX1_250 ( );
FILL FILL_0_OAI21X1_117 ( );
FILL FILL_1_OAI21X1_117 ( );
FILL FILL_0_OAI21X1_116 ( );
FILL FILL_1_OAI21X1_116 ( );
FILL FILL_2_OAI21X1_116 ( );
FILL FILL_0_OAI21X1_86 ( );
FILL FILL_1_OAI21X1_86 ( );
FILL FILL_0_OAI21X1_87 ( );
FILL FILL_1_OAI21X1_87 ( );
FILL FILL_0_DFFPOSX1_235 ( );
FILL FILL_1_DFFPOSX1_235 ( );
FILL FILL_2_DFFPOSX1_235 ( );
FILL FILL_3_DFFPOSX1_235 ( );
FILL FILL_4_DFFPOSX1_235 ( );
FILL FILL_5_DFFPOSX1_235 ( );
FILL FILL_0_BUFX2_920 ( );
FILL FILL_1_BUFX2_920 ( );
FILL FILL_0_BUFX2_56 ( );
FILL FILL_0_BUFX2_189 ( );
FILL FILL_0_INVX2_181 ( );
FILL FILL_0_BUFX2_934 ( );
FILL FILL_1_BUFX2_934 ( );
FILL FILL_0_DFFPOSX1_263 ( );
FILL FILL_1_DFFPOSX1_263 ( );
FILL FILL_2_DFFPOSX1_263 ( );
FILL FILL_3_DFFPOSX1_263 ( );
FILL FILL_4_DFFPOSX1_263 ( );
FILL FILL_5_DFFPOSX1_263 ( );
FILL FILL_6_DFFPOSX1_263 ( );
FILL FILL_0_OAI21X1_142 ( );
FILL FILL_1_OAI21X1_142 ( );
FILL FILL_2_OAI21X1_142 ( );
FILL FILL_0_OAI21X1_143 ( );
FILL FILL_1_OAI21X1_143 ( );
FILL FILL_0_BUFX2_870 ( );
FILL FILL_0_BUFX2_194 ( );
FILL FILL_0_DFFPOSX1_937 ( );
FILL FILL_1_DFFPOSX1_937 ( );
FILL FILL_2_DFFPOSX1_937 ( );
FILL FILL_3_DFFPOSX1_937 ( );
FILL FILL_4_DFFPOSX1_937 ( );
FILL FILL_5_DFFPOSX1_937 ( );
FILL FILL_0_OAI21X1_1387 ( );
FILL FILL_1_OAI21X1_1387 ( );
FILL FILL_0_OAI21X1_1386 ( );
FILL FILL_1_OAI21X1_1386 ( );
FILL FILL_2_OAI21X1_1386 ( );
FILL FILL_0_BUFX4_376 ( );
FILL FILL_1_BUFX4_376 ( );
FILL FILL_2_BUFX4_376 ( );
FILL FILL_0_BUFX4_180 ( );
FILL FILL_1_BUFX4_180 ( );
FILL FILL_0_BUFX4_46 ( );
FILL FILL_1_BUFX4_46 ( );
FILL FILL_2_BUFX4_46 ( );
FILL FILL_0_OAI21X1_1018 ( );
FILL FILL_1_OAI21X1_1018 ( );
FILL FILL_0_BUFX4_183 ( );
FILL FILL_1_BUFX4_183 ( );
FILL FILL_2_BUFX4_183 ( );
FILL FILL_0_BUFX4_49 ( );
FILL FILL_1_BUFX4_49 ( );
FILL FILL_0_DFFPOSX1_463 ( );
FILL FILL_1_DFFPOSX1_463 ( );
FILL FILL_2_DFFPOSX1_463 ( );
FILL FILL_3_DFFPOSX1_463 ( );
FILL FILL_4_DFFPOSX1_463 ( );
FILL FILL_5_DFFPOSX1_463 ( );
FILL FILL_0_BUFX4_282 ( );
FILL FILL_1_BUFX4_282 ( );
FILL FILL_0_BUFX2_998 ( );
FILL FILL_1_BUFX2_998 ( );
FILL FILL_0_BUFX2_646 ( );
FILL FILL_0_DFFPOSX1_327 ( );
FILL FILL_1_DFFPOSX1_327 ( );
FILL FILL_2_DFFPOSX1_327 ( );
FILL FILL_3_DFFPOSX1_327 ( );
FILL FILL_4_DFFPOSX1_327 ( );
FILL FILL_5_DFFPOSX1_327 ( );
FILL FILL_0_OAI21X1_271 ( );
FILL FILL_1_OAI21X1_271 ( );
FILL FILL_0_OAI21X1_270 ( );
FILL FILL_1_OAI21X1_270 ( );
FILL FILL_0_BUFX4_2 ( );
FILL FILL_1_BUFX4_2 ( );
FILL FILL_0_DFFPOSX1_555 ( );
FILL FILL_1_DFFPOSX1_555 ( );
FILL FILL_2_DFFPOSX1_555 ( );
FILL FILL_3_DFFPOSX1_555 ( );
FILL FILL_4_DFFPOSX1_555 ( );
FILL FILL_5_DFFPOSX1_555 ( );
FILL FILL_6_DFFPOSX1_555 ( );
FILL FILL_0_OAI21X1_681 ( );
FILL FILL_1_OAI21X1_681 ( );
FILL FILL_0_OAI21X1_680 ( );
FILL FILL_1_OAI21X1_680 ( );
FILL FILL_2_OAI21X1_680 ( );
FILL FILL_0_BUFX2_431 ( );
FILL FILL_1_BUFX2_431 ( );
FILL FILL_0_BUFX4_290 ( );
FILL FILL_1_BUFX4_290 ( );
FILL FILL_0_BUFX4_252 ( );
FILL FILL_1_BUFX4_252 ( );
FILL FILL_0_BUFX4_9 ( );
FILL FILL_1_BUFX4_9 ( );
FILL FILL_0_OAI21X1_607 ( );
FILL FILL_1_OAI21X1_607 ( );
FILL FILL_0_BUFX4_204 ( );
FILL FILL_1_BUFX4_204 ( );
FILL FILL_0_OAI21X1_608 ( );
FILL FILL_1_OAI21X1_608 ( );
FILL FILL_0_OAI21X1_631 ( );
FILL FILL_1_OAI21X1_631 ( );
FILL FILL_2_OAI21X1_631 ( );
FILL FILL_0_OAI21X1_633 ( );
FILL FILL_1_OAI21X1_633 ( );
FILL FILL_2_OAI21X1_633 ( );
FILL FILL_0_OAI21X1_632 ( );
FILL FILL_1_OAI21X1_632 ( );
FILL FILL_0_DFFPOSX1_399 ( );
FILL FILL_1_DFFPOSX1_399 ( );
FILL FILL_2_DFFPOSX1_399 ( );
FILL FILL_3_DFFPOSX1_399 ( );
FILL FILL_4_DFFPOSX1_399 ( );
FILL FILL_5_DFFPOSX1_399 ( );
FILL FILL_6_DFFPOSX1_399 ( );
FILL FILL_0_NOR2X1_43 ( );
FILL FILL_1_NOR2X1_43 ( );
FILL FILL_0_AOI21X1_19 ( );
FILL FILL_1_AOI21X1_19 ( );
FILL FILL_0_NAND2X1_483 ( );
FILL FILL_1_NAND2X1_483 ( );
FILL FILL_0_INVX1_19 ( );
FILL FILL_0_OAI21X1_810 ( );
FILL FILL_1_OAI21X1_810 ( );
FILL FILL_2_OAI21X1_810 ( );
FILL FILL_0_NAND2X1_243 ( );
FILL FILL_1_NAND2X1_243 ( );
FILL FILL_0_INVX2_45 ( );
FILL FILL_0_DFFPOSX1_395 ( );
FILL FILL_1_DFFPOSX1_395 ( );
FILL FILL_2_DFFPOSX1_395 ( );
FILL FILL_3_DFFPOSX1_395 ( );
FILL FILL_4_DFFPOSX1_395 ( );
FILL FILL_5_DFFPOSX1_395 ( );
FILL FILL_6_DFFPOSX1_395 ( );
FILL FILL_0_NAND2X1_111 ( );
FILL FILL_0_BUFX4_213 ( );
FILL FILL_1_BUFX4_213 ( );
FILL FILL_0_NAND2X1_214 ( );
FILL FILL_1_NAND2X1_214 ( );
FILL FILL_0_OAI21X1_457 ( );
FILL FILL_1_OAI21X1_457 ( );
FILL FILL_0_NAND2X1_253 ( );
FILL FILL_0_INVX2_47 ( );
FILL FILL_0_NAND2X1_254 ( );
FILL FILL_0_OAI21X1_488 ( );
FILL FILL_1_OAI21X1_488 ( );
FILL FILL_2_OAI21X1_488 ( );
FILL FILL_0_INVX2_37 ( );
FILL FILL_0_NAND3X1_35 ( );
FILL FILL_1_NAND3X1_35 ( );
FILL FILL_0_NAND3X1_36 ( );
FILL FILL_1_NAND3X1_36 ( );
FILL FILL_0_NOR3X1_10 ( );
FILL FILL_1_NOR3X1_10 ( );
FILL FILL_2_NOR3X1_10 ( );
FILL FILL_3_NOR3X1_10 ( );
FILL FILL_0_INVX1_44 ( );
FILL FILL_0_AOI21X1_5 ( );
FILL FILL_1_AOI21X1_5 ( );
FILL FILL_0_OAI21X1_493 ( );
FILL FILL_1_OAI21X1_493 ( );
FILL FILL_0_NOR2X1_120 ( );
FILL FILL_1_NOR2X1_120 ( );
FILL FILL_0_NAND3X1_37 ( );
FILL FILL_1_NAND3X1_37 ( );
FILL FILL_0_NAND2X1_335 ( );
FILL FILL_1_NAND2X1_335 ( );
FILL FILL_0_BUFX2_615 ( );
FILL FILL_0_NAND2X1_337 ( );
FILL FILL_0_OAI21X1_762 ( );
FILL FILL_1_OAI21X1_762 ( );
FILL FILL_0_OAI21X1_763 ( );
FILL FILL_1_OAI21X1_763 ( );
FILL FILL_0_OAI21X1_759 ( );
FILL FILL_1_OAI21X1_759 ( );
FILL FILL_0_DFFPOSX1_87 ( );
FILL FILL_1_DFFPOSX1_87 ( );
FILL FILL_2_DFFPOSX1_87 ( );
FILL FILL_3_DFFPOSX1_87 ( );
FILL FILL_4_DFFPOSX1_87 ( );
FILL FILL_5_DFFPOSX1_87 ( );
FILL FILL_6_DFFPOSX1_87 ( );
FILL FILL_0_OAI21X1_1749 ( );
FILL FILL_1_OAI21X1_1749 ( );
FILL FILL_2_OAI21X1_1749 ( );
FILL FILL_0_OAI21X1_1748 ( );
FILL FILL_1_OAI21X1_1748 ( );
FILL FILL_0_OAI21X1_717 ( );
FILL FILL_1_OAI21X1_717 ( );
FILL FILL_0_NAND2X1_91 ( );
FILL FILL_1_NAND2X1_91 ( );
FILL FILL_0_DFFPOSX1_375 ( );
FILL FILL_1_DFFPOSX1_375 ( );
FILL FILL_2_DFFPOSX1_375 ( );
FILL FILL_3_DFFPOSX1_375 ( );
FILL FILL_4_DFFPOSX1_375 ( );
FILL FILL_5_DFFPOSX1_375 ( );
FILL FILL_6_DFFPOSX1_375 ( );
FILL FILL_0_OAI21X1_347 ( );
FILL FILL_1_OAI21X1_347 ( );
FILL FILL_0_CLKBUF1_1 ( );
FILL FILL_1_CLKBUF1_1 ( );
FILL FILL_2_CLKBUF1_1 ( );
FILL FILL_3_CLKBUF1_1 ( );
FILL FILL_4_CLKBUF1_1 ( );
FILL FILL_0_OAI21X1_384 ( );
FILL FILL_1_OAI21X1_384 ( );
FILL FILL_0_NAND2X1_128 ( );
FILL FILL_1_NAND2X1_128 ( );
FILL FILL_0_BUFX2_620 ( );
FILL FILL_0_BUFX4_91 ( );
FILL FILL_1_BUFX4_91 ( );
FILL FILL_0_OAI21X1_738 ( );
FILL FILL_1_OAI21X1_738 ( );
FILL FILL_2_OAI21X1_738 ( );
FILL FILL_0_BUFX2_542 ( );
FILL FILL_0_NAND2X1_98 ( );
FILL FILL_1_NAND2X1_98 ( );
FILL FILL_0_OAI21X1_737 ( );
FILL FILL_1_OAI21X1_737 ( );
FILL FILL_0_BUFX4_283 ( );
FILL FILL_1_BUFX4_283 ( );
FILL FILL_0_BUFX4_147 ( );
FILL FILL_1_BUFX4_147 ( );
FILL FILL_0_BUFX4_209 ( );
FILL FILL_1_BUFX4_209 ( );
FILL FILL_2_BUFX4_209 ( );
FILL FILL_0_DFFPOSX1_93 ( );
FILL FILL_1_DFFPOSX1_93 ( );
FILL FILL_2_DFFPOSX1_93 ( );
FILL FILL_3_DFFPOSX1_93 ( );
FILL FILL_4_DFFPOSX1_93 ( );
FILL FILL_5_DFFPOSX1_93 ( );
FILL FILL_0_OAI21X1_437 ( );
FILL FILL_1_OAI21X1_437 ( );
FILL FILL_0_DFFPOSX1_836 ( );
FILL FILL_1_DFFPOSX1_836 ( );
FILL FILL_2_DFFPOSX1_836 ( );
FILL FILL_3_DFFPOSX1_836 ( );
FILL FILL_4_DFFPOSX1_836 ( );
FILL FILL_5_DFFPOSX1_836 ( );
FILL FILL_0_NAND2X1_524 ( );
FILL FILL_1_NAND2X1_524 ( );
FILL FILL_0_OAI21X1_1148 ( );
FILL FILL_1_OAI21X1_1148 ( );
FILL FILL_0_NAND2X1_97 ( );
FILL FILL_1_NAND2X1_97 ( );
FILL FILL_0_INVX1_203 ( );
FILL FILL_0_NAND2X1_600 ( );
FILL FILL_0_NOR2X1_190 ( );
FILL FILL_0_NAND3X1_54 ( );
FILL FILL_1_NAND3X1_54 ( );
FILL FILL_2_NAND3X1_54 ( );
FILL FILL_0_INVX1_204 ( );
FILL FILL_0_BUFX4_317 ( );
FILL FILL_1_BUFX4_317 ( );
FILL FILL_2_BUFX4_317 ( );
FILL FILL_0_OR2X2_19 ( );
FILL FILL_1_OR2X2_19 ( );
FILL FILL_0_NOR2X1_191 ( );
FILL FILL_1_NOR2X1_191 ( );
FILL FILL_0_NOR2X1_193 ( );
FILL FILL_1_NOR2X1_193 ( );
FILL FILL_0_NAND2X1_606 ( );
FILL FILL_0_OAI21X1_1289 ( );
FILL FILL_1_OAI21X1_1289 ( );
FILL FILL_2_OAI21X1_1289 ( );
FILL FILL_0_OAI21X1_1288 ( );
FILL FILL_1_OAI21X1_1288 ( );
FILL FILL_0_OAI21X1_1290 ( );
FILL FILL_1_OAI21X1_1290 ( );
FILL FILL_0_BUFX2_151 ( );
FILL FILL_1_BUFX2_151 ( );
FILL FILL_0_INVX1_205 ( );
FILL FILL_0_NOR2X1_192 ( );
FILL FILL_1_NOR2X1_192 ( );
FILL FILL_0_XNOR2X1_80 ( );
FILL FILL_1_XNOR2X1_80 ( );
FILL FILL_2_XNOR2X1_80 ( );
FILL FILL_0_DFFPOSX1_321 ( );
FILL FILL_1_DFFPOSX1_321 ( );
FILL FILL_2_DFFPOSX1_321 ( );
FILL FILL_3_DFFPOSX1_321 ( );
FILL FILL_4_DFFPOSX1_321 ( );
FILL FILL_5_DFFPOSX1_321 ( );
FILL FILL_6_DFFPOSX1_321 ( );
FILL FILL_0_OAI21X1_1284 ( );
FILL FILL_1_OAI21X1_1284 ( );
FILL FILL_0_OAI21X1_1283 ( );
FILL FILL_1_OAI21X1_1283 ( );
FILL FILL_2_OAI21X1_1283 ( );
FILL FILL_0_OAI21X1_1780 ( );
FILL FILL_1_OAI21X1_1780 ( );
FILL FILL_0_NAND2X1_721 ( );
FILL FILL_1_NAND2X1_721 ( );
FILL FILL_0_BUFX2_167 ( );
FILL FILL_1_BUFX2_167 ( );
FILL FILL_0_DFFPOSX1_916 ( );
FILL FILL_1_DFFPOSX1_916 ( );
FILL FILL_2_DFFPOSX1_916 ( );
FILL FILL_3_DFFPOSX1_916 ( );
FILL FILL_4_DFFPOSX1_916 ( );
FILL FILL_5_DFFPOSX1_916 ( );
FILL FILL_0_BUFX2_833 ( );
FILL FILL_0_NOR2X1_162 ( );
FILL FILL_1_NOR2X1_162 ( );
FILL FILL_0_NAND3X1_45 ( );
FILL FILL_1_NAND3X1_45 ( );
FILL FILL_0_NAND2X1_617 ( );
FILL FILL_1_NAND2X1_617 ( );
FILL FILL_0_NOR2X1_204 ( );
FILL FILL_0_OAI21X1_1516 ( );
FILL FILL_1_OAI21X1_1516 ( );
FILL FILL_0_OAI21X1_1518 ( );
FILL FILL_1_OAI21X1_1518 ( );
FILL FILL_0_INVX2_81 ( );
FILL FILL_0_OAI21X1_1517 ( );
FILL FILL_1_OAI21X1_1517 ( );
FILL FILL_0_DFFPOSX1_918 ( );
FILL FILL_1_DFFPOSX1_918 ( );
FILL FILL_2_DFFPOSX1_918 ( );
FILL FILL_3_DFFPOSX1_918 ( );
FILL FILL_4_DFFPOSX1_918 ( );
FILL FILL_5_DFFPOSX1_918 ( );
FILL FILL_0_NAND3X1_46 ( );
FILL FILL_1_NAND3X1_46 ( );
FILL FILL_0_OAI21X1_1335 ( );
FILL FILL_1_OAI21X1_1335 ( );
FILL FILL_0_INVX2_111 ( );
FILL FILL_0_AOI21X1_39 ( );
FILL FILL_1_AOI21X1_39 ( );
FILL FILL_0_BUFX4_121 ( );
FILL FILL_1_BUFX4_121 ( );
FILL FILL_0_NAND2X1_557 ( );
FILL FILL_1_NAND2X1_557 ( );
FILL FILL_0_OAI21X1_1174 ( );
FILL FILL_1_OAI21X1_1174 ( );
FILL FILL_0_DFFPOSX1_854 ( );
FILL FILL_1_DFFPOSX1_854 ( );
FILL FILL_2_DFFPOSX1_854 ( );
FILL FILL_3_DFFPOSX1_854 ( );
FILL FILL_4_DFFPOSX1_854 ( );
FILL FILL_5_DFFPOSX1_854 ( );
FILL FILL_6_DFFPOSX1_854 ( );
FILL FILL_0_NAND2X1_558 ( );
FILL FILL_1_NAND2X1_558 ( );
FILL FILL_0_BUFX2_106 ( );
FILL FILL_1_BUFX2_106 ( );
FILL FILL_0_BUFX4_270 ( );
FILL FILL_1_BUFX4_270 ( );
FILL FILL_0_BUFX4_38 ( );
FILL FILL_1_BUFX4_38 ( );
FILL FILL_0_BUFX4_47 ( );
FILL FILL_1_BUFX4_47 ( );
FILL FILL_0_BUFX4_51 ( );
FILL FILL_1_BUFX4_51 ( );
FILL FILL_0_OAI21X1_1528 ( );
FILL FILL_1_OAI21X1_1528 ( );
FILL FILL_2_OAI21X1_1528 ( );
FILL FILL_0_BUFX2_45 ( );
FILL FILL_1_BUFX2_45 ( );
FILL FILL_0_DFFPOSX1_932 ( );
FILL FILL_1_DFFPOSX1_932 ( );
FILL FILL_2_DFFPOSX1_932 ( );
FILL FILL_3_DFFPOSX1_932 ( );
FILL FILL_4_DFFPOSX1_932 ( );
FILL FILL_5_DFFPOSX1_932 ( );
FILL FILL_6_DFFPOSX1_932 ( );
FILL FILL_0_OAI21X1_1381 ( );
FILL FILL_1_OAI21X1_1381 ( );
FILL FILL_0_BUFX4_162 ( );
FILL FILL_1_BUFX4_162 ( );
FILL FILL_0_OAI21X1_1333 ( );
FILL FILL_1_OAI21X1_1333 ( );
FILL FILL_0_OAI21X1_1375 ( );
FILL FILL_1_OAI21X1_1375 ( );
FILL FILL_0_OAI21X1_1374 ( );
FILL FILL_1_OAI21X1_1374 ( );
FILL FILL_0_OAI21X1_244 ( );
FILL FILL_1_OAI21X1_244 ( );
FILL FILL_0_OAI21X1_245 ( );
FILL FILL_1_OAI21X1_245 ( );
FILL FILL_0_DFFPOSX1_314 ( );
FILL FILL_1_DFFPOSX1_314 ( );
FILL FILL_2_DFFPOSX1_314 ( );
FILL FILL_3_DFFPOSX1_314 ( );
FILL FILL_4_DFFPOSX1_314 ( );
FILL FILL_5_DFFPOSX1_314 ( );
FILL FILL_0_DFFPOSX1_299 ( );
FILL FILL_1_DFFPOSX1_299 ( );
FILL FILL_2_DFFPOSX1_299 ( );
FILL FILL_3_DFFPOSX1_299 ( );
FILL FILL_4_DFFPOSX1_299 ( );
FILL FILL_5_DFFPOSX1_299 ( );
FILL FILL_6_DFFPOSX1_299 ( );
FILL FILL_0_OAI21X1_214 ( );
FILL FILL_1_OAI21X1_214 ( );
FILL FILL_2_OAI21X1_214 ( );
FILL FILL_0_OAI21X1_215 ( );
FILL FILL_1_OAI21X1_215 ( );
FILL FILL_0_OAI21X1_1781 ( );
FILL FILL_1_OAI21X1_1781 ( );
FILL FILL_0_NAND2X1_722 ( );
FILL FILL_1_NAND2X1_722 ( );
FILL FILL_0_DFFPOSX1_107 ( );
FILL FILL_1_DFFPOSX1_107 ( );
FILL FILL_2_DFFPOSX1_107 ( );
FILL FILL_3_DFFPOSX1_107 ( );
FILL FILL_4_DFFPOSX1_107 ( );
FILL FILL_5_DFFPOSX1_107 ( );
FILL FILL_6_DFFPOSX1_107 ( );
FILL FILL_0_BUFX2_838 ( );
FILL FILL_1_BUFX2_838 ( );
FILL FILL_0_BUFX2_966 ( );
FILL FILL_0_DFFPOSX1_642 ( );
FILL FILL_1_DFFPOSX1_642 ( );
FILL FILL_2_DFFPOSX1_642 ( );
FILL FILL_3_DFFPOSX1_642 ( );
FILL FILL_4_DFFPOSX1_642 ( );
FILL FILL_5_DFFPOSX1_642 ( );
FILL FILL_6_DFFPOSX1_642 ( );
FILL FILL_0_INVX1_56 ( );
FILL FILL_0_INVX1_157 ( );
FILL FILL_0_BUFX2_336 ( );
FILL FILL_1_BUFX2_336 ( );
FILL FILL_0_INVX2_197 ( );
FILL FILL_1_INVX2_197 ( );
FILL FILL_0_BUFX2_810 ( );
FILL FILL_0_NAND2X1_345 ( );
FILL FILL_1_NAND2X1_345 ( );
FILL FILL_0_BUFX2_326 ( );
FILL FILL_0_BUFX2_711 ( );
FILL FILL_0_INVX1_131 ( );
FILL FILL_0_NAND2X1_364 ( );
FILL FILL_1_NAND2X1_364 ( );
FILL FILL_0_INVX1_156 ( );
FILL FILL_0_BUFX2_321 ( );
FILL FILL_0_INVX1_71 ( );
FILL FILL_0_INVX1_82 ( );
FILL FILL_0_BUFX4_265 ( );
FILL FILL_1_BUFX4_265 ( );
FILL FILL_0_DFFPOSX1_22 ( );
FILL FILL_1_DFFPOSX1_22 ( );
FILL FILL_2_DFFPOSX1_22 ( );
FILL FILL_3_DFFPOSX1_22 ( );
FILL FILL_4_DFFPOSX1_22 ( );
FILL FILL_5_DFFPOSX1_22 ( );
FILL FILL_6_DFFPOSX1_22 ( );
FILL FILL_0_OAI21X1_1632 ( );
FILL FILL_1_OAI21X1_1632 ( );
FILL FILL_2_OAI21X1_1632 ( );
FILL FILL_0_BUFX2_755 ( );
FILL FILL_0_DFFPOSX1_1022 ( );
FILL FILL_1_DFFPOSX1_1022 ( );
FILL FILL_2_DFFPOSX1_1022 ( );
FILL FILL_3_DFFPOSX1_1022 ( );
FILL FILL_4_DFFPOSX1_1022 ( );
FILL FILL_5_DFFPOSX1_1022 ( );
FILL FILL_0_OAI21X1_1599 ( );
FILL FILL_1_OAI21X1_1599 ( );
FILL FILL_0_OAI21X1_1747 ( );
FILL FILL_1_OAI21X1_1747 ( );
FILL FILL_0_OAI21X1_1746 ( );
FILL FILL_1_OAI21X1_1746 ( );
FILL FILL_0_DFFPOSX1_86 ( );
FILL FILL_1_DFFPOSX1_86 ( );
FILL FILL_2_DFFPOSX1_86 ( );
FILL FILL_3_DFFPOSX1_86 ( );
FILL FILL_4_DFFPOSX1_86 ( );
FILL FILL_5_DFFPOSX1_86 ( );
FILL FILL_0_INVX1_164 ( );
FILL FILL_0_OAI21X1_1019 ( );
FILL FILL_1_OAI21X1_1019 ( );
FILL FILL_0_DFFPOSX1_735 ( );
FILL FILL_1_DFFPOSX1_735 ( );
FILL FILL_2_DFFPOSX1_735 ( );
FILL FILL_3_DFFPOSX1_735 ( );
FILL FILL_4_DFFPOSX1_735 ( );
FILL FILL_5_DFFPOSX1_735 ( );
FILL FILL_6_DFFPOSX1_735 ( );
FILL FILL_0_CLKBUF1_73 ( );
FILL FILL_1_CLKBUF1_73 ( );
FILL FILL_2_CLKBUF1_73 ( );
FILL FILL_3_CLKBUF1_73 ( );
FILL FILL_4_CLKBUF1_73 ( );
FILL FILL_0_BUFX4_98 ( );
FILL FILL_1_BUFX4_98 ( );
FILL FILL_2_BUFX4_98 ( );
FILL FILL_0_OAI21X1_475 ( );
FILL FILL_1_OAI21X1_475 ( );
FILL FILL_0_BUFX2_585 ( );
FILL FILL_1_BUFX2_585 ( );
FILL FILL_0_OAI21X1_659 ( );
FILL FILL_1_OAI21X1_659 ( );
FILL FILL_0_DFFPOSX1_548 ( );
FILL FILL_1_DFFPOSX1_548 ( );
FILL FILL_2_DFFPOSX1_548 ( );
FILL FILL_3_DFFPOSX1_548 ( );
FILL FILL_4_DFFPOSX1_548 ( );
FILL FILL_5_DFFPOSX1_548 ( );
FILL FILL_0_OAI21X1_658 ( );
FILL FILL_1_OAI21X1_658 ( );
FILL FILL_0_CLKBUF1_91 ( );
FILL FILL_1_CLKBUF1_91 ( );
FILL FILL_2_CLKBUF1_91 ( );
FILL FILL_3_CLKBUF1_91 ( );
FILL FILL_4_CLKBUF1_91 ( );
FILL FILL_0_BUFX4_145 ( );
FILL FILL_1_BUFX4_145 ( );
FILL FILL_0_BUFX2_569 ( );
FILL FILL_1_BUFX2_569 ( );
FILL FILL_0_DFFPOSX1_535 ( );
FILL FILL_1_DFFPOSX1_535 ( );
FILL FILL_2_DFFPOSX1_535 ( );
FILL FILL_3_DFFPOSX1_535 ( );
FILL FILL_4_DFFPOSX1_535 ( );
FILL FILL_5_DFFPOSX1_535 ( );
FILL FILL_0_OAI21X1_630 ( );
FILL FILL_1_OAI21X1_630 ( );
FILL FILL_0_BUFX4_93 ( );
FILL FILL_1_BUFX4_93 ( );
FILL FILL_0_BUFX4_112 ( );
FILL FILL_1_BUFX4_112 ( );
FILL FILL_0_DFFPOSX1_526 ( );
FILL FILL_1_DFFPOSX1_526 ( );
FILL FILL_2_DFFPOSX1_526 ( );
FILL FILL_3_DFFPOSX1_526 ( );
FILL FILL_4_DFFPOSX1_526 ( );
FILL FILL_5_DFFPOSX1_526 ( );
FILL FILL_0_DFFPOSX1_536 ( );
FILL FILL_1_DFFPOSX1_536 ( );
FILL FILL_2_DFFPOSX1_536 ( );
FILL FILL_3_DFFPOSX1_536 ( );
FILL FILL_4_DFFPOSX1_536 ( );
FILL FILL_5_DFFPOSX1_536 ( );
FILL FILL_6_DFFPOSX1_536 ( );
FILL FILL_0_NAND2X1_234 ( );
FILL FILL_1_NAND2X1_234 ( );
FILL FILL_0_NAND2X1_236 ( );
FILL FILL_0_NAND2X1_235 ( );
FILL FILL_1_NAND2X1_235 ( );
FILL FILL_0_OAI21X1_473 ( );
FILL FILL_1_OAI21X1_473 ( );
FILL FILL_0_XNOR2X1_38 ( );
FILL FILL_1_XNOR2X1_38 ( );
FILL FILL_2_XNOR2X1_38 ( );
FILL FILL_3_XNOR2X1_38 ( );
FILL FILL_0_OAI21X1_472 ( );
FILL FILL_1_OAI21X1_472 ( );
FILL FILL_0_INVX2_34 ( );
FILL FILL_0_OAI21X1_811 ( );
FILL FILL_1_OAI21X1_811 ( );
FILL FILL_0_NOR2X1_51 ( );
FILL FILL_0_OAI21X1_806 ( );
FILL FILL_1_OAI21X1_806 ( );
FILL FILL_0_OAI21X1_807 ( );
FILL FILL_1_OAI21X1_807 ( );
FILL FILL_0_OR2X2_13 ( );
FILL FILL_1_OR2X2_13 ( );
FILL FILL_0_BUFX4_62 ( );
FILL FILL_1_BUFX4_62 ( );
FILL FILL_0_BUFX4_18 ( );
FILL FILL_1_BUFX4_18 ( );
FILL FILL_0_DFFPOSX1_459 ( );
FILL FILL_1_DFFPOSX1_459 ( );
FILL FILL_2_DFFPOSX1_459 ( );
FILL FILL_3_DFFPOSX1_459 ( );
FILL FILL_4_DFFPOSX1_459 ( );
FILL FILL_5_DFFPOSX1_459 ( );
FILL FILL_0_NOR2X1_52 ( );
FILL FILL_1_NOR2X1_52 ( );
FILL FILL_0_NAND2X1_252 ( );
FILL FILL_1_NAND2X1_252 ( );
FILL FILL_0_NOR2X1_53 ( );
FILL FILL_0_NAND2X1_250 ( );
FILL FILL_1_NAND2X1_250 ( );
FILL FILL_0_OAI21X1_486 ( );
FILL FILL_1_OAI21X1_486 ( );
FILL FILL_0_OAI21X1_487 ( );
FILL FILL_1_OAI21X1_487 ( );
FILL FILL_2_OAI21X1_487 ( );
FILL FILL_0_OAI21X1_822 ( );
FILL FILL_1_OAI21X1_822 ( );
FILL FILL_0_NAND2X1_260 ( );
FILL FILL_1_NAND2X1_260 ( );
FILL FILL_0_INVX1_23 ( );
FILL FILL_0_NAND2X1_262 ( );
FILL FILL_0_OAI21X1_499 ( );
FILL FILL_1_OAI21X1_499 ( );
FILL FILL_0_INVX2_39 ( );
FILL FILL_0_OAI21X1_842 ( );
FILL FILL_1_OAI21X1_842 ( );
FILL FILL_0_NOR3X1_11 ( );
FILL FILL_1_NOR3X1_11 ( );
FILL FILL_2_NOR3X1_11 ( );
FILL FILL_3_NOR3X1_11 ( );
FILL FILL_0_NAND2X1_336 ( );
FILL FILL_1_NAND2X1_336 ( );
FILL FILL_0_BUFX2_598 ( );
FILL FILL_1_BUFX2_598 ( );
FILL FILL_0_BUFX2_756 ( );
FILL FILL_1_BUFX2_756 ( );
FILL FILL_0_DFFPOSX1_583 ( );
FILL FILL_1_DFFPOSX1_583 ( );
FILL FILL_2_DFFPOSX1_583 ( );
FILL FILL_3_DFFPOSX1_583 ( );
FILL FILL_4_DFFPOSX1_583 ( );
FILL FILL_5_DFFPOSX1_583 ( );
FILL FILL_6_DFFPOSX1_583 ( );
FILL FILL_0_BUFX4_221 ( );
FILL FILL_1_BUFX4_221 ( );
FILL FILL_0_BUFX4_25 ( );
FILL FILL_1_BUFX4_25 ( );
FILL FILL_0_XNOR2X1_15 ( );
FILL FILL_1_XNOR2X1_15 ( );
FILL FILL_2_XNOR2X1_15 ( );
FILL FILL_0_CLKBUF1_19 ( );
FILL FILL_1_CLKBUF1_19 ( );
FILL FILL_2_CLKBUF1_19 ( );
FILL FILL_3_CLKBUF1_19 ( );
FILL FILL_4_CLKBUF1_19 ( );
FILL FILL_0_DFFPOSX1_439 ( );
FILL FILL_1_DFFPOSX1_439 ( );
FILL FILL_2_DFFPOSX1_439 ( );
FILL FILL_3_DFFPOSX1_439 ( );
FILL FILL_4_DFFPOSX1_439 ( );
FILL FILL_5_DFFPOSX1_439 ( );
FILL FILL_0_OAI21X1_454 ( );
FILL FILL_1_OAI21X1_454 ( );
FILL FILL_0_NAND2X1_210 ( );
FILL FILL_1_NAND2X1_210 ( );
FILL FILL_0_BUFX4_224 ( );
FILL FILL_1_BUFX4_224 ( );
FILL FILL_0_DFFPOSX1_109 ( );
FILL FILL_1_DFFPOSX1_109 ( );
FILL FILL_2_DFFPOSX1_109 ( );
FILL FILL_3_DFFPOSX1_109 ( );
FILL FILL_4_DFFPOSX1_109 ( );
FILL FILL_5_DFFPOSX1_109 ( );
FILL FILL_6_DFFPOSX1_109 ( );
FILL FILL_0_DFFPOSX1_575 ( );
FILL FILL_1_DFFPOSX1_575 ( );
FILL FILL_2_DFFPOSX1_575 ( );
FILL FILL_3_DFFPOSX1_575 ( );
FILL FILL_4_DFFPOSX1_575 ( );
FILL FILL_5_DFFPOSX1_575 ( );
FILL FILL_6_DFFPOSX1_575 ( );
FILL FILL_0_CLKBUF1_50 ( );
FILL FILL_1_CLKBUF1_50 ( );
FILL FILL_2_CLKBUF1_50 ( );
FILL FILL_3_CLKBUF1_50 ( );
FILL FILL_4_CLKBUF1_50 ( );
FILL FILL_0_OAI21X1_445 ( );
FILL FILL_1_OAI21X1_445 ( );
FILL FILL_0_DFFPOSX1_450 ( );
FILL FILL_1_DFFPOSX1_450 ( );
FILL FILL_2_DFFPOSX1_450 ( );
FILL FILL_3_DFFPOSX1_450 ( );
FILL FILL_4_DFFPOSX1_450 ( );
FILL FILL_5_DFFPOSX1_450 ( );
FILL FILL_0_OAI21X1_1697 ( );
FILL FILL_1_OAI21X1_1697 ( );
FILL FILL_0_DFFPOSX1_445 ( );
FILL FILL_1_DFFPOSX1_445 ( );
FILL FILL_2_DFFPOSX1_445 ( );
FILL FILL_3_DFFPOSX1_445 ( );
FILL FILL_4_DFFPOSX1_445 ( );
FILL FILL_5_DFFPOSX1_445 ( );
FILL FILL_6_DFFPOSX1_445 ( );
FILL FILL_0_BUFX4_334 ( );
FILL FILL_1_BUFX4_334 ( );
FILL FILL_0_OAI21X1_1639 ( );
FILL FILL_1_OAI21X1_1639 ( );
FILL FILL_0_NAND2X1_707 ( );
FILL FILL_0_BUFX4_311 ( );
FILL FILL_1_BUFX4_311 ( );
FILL FILL_2_BUFX4_311 ( );
FILL FILL_0_INVX4_51 ( );
FILL FILL_0_BUFX4_255 ( );
FILL FILL_1_BUFX4_255 ( );
FILL FILL_0_CLKBUF1_35 ( );
FILL FILL_1_CLKBUF1_35 ( );
FILL FILL_2_CLKBUF1_35 ( );
FILL FILL_3_CLKBUF1_35 ( );
FILL FILL_4_CLKBUF1_35 ( );
FILL FILL_0_XNOR2X1_79 ( );
FILL FILL_1_XNOR2X1_79 ( );
FILL FILL_2_XNOR2X1_79 ( );
FILL FILL_0_INVX1_206 ( );
FILL FILL_0_NAND2X1_605 ( );
FILL FILL_1_NAND2X1_605 ( );
FILL FILL_0_XNOR2X1_65 ( );
FILL FILL_1_XNOR2X1_65 ( );
FILL FILL_2_XNOR2X1_65 ( );
FILL FILL_3_XNOR2X1_65 ( );
FILL FILL_0_AOI21X1_47 ( );
FILL FILL_1_AOI21X1_47 ( );
FILL FILL_0_INVX1_207 ( );
FILL FILL_0_OAI21X1_1286 ( );
FILL FILL_1_OAI21X1_1286 ( );
FILL FILL_0_NAND2X1_604 ( );
FILL FILL_0_DFFPOSX1_253 ( );
FILL FILL_1_DFFPOSX1_253 ( );
FILL FILL_2_DFFPOSX1_253 ( );
FILL FILL_3_DFFPOSX1_253 ( );
FILL FILL_4_DFFPOSX1_253 ( );
FILL FILL_5_DFFPOSX1_253 ( );
FILL FILL_0_AND2X2_28 ( );
FILL FILL_1_AND2X2_28 ( );
FILL FILL_0_BUFX4_117 ( );
FILL FILL_1_BUFX4_117 ( );
FILL FILL_0_NAND3X1_42 ( );
FILL FILL_1_NAND3X1_42 ( );
FILL FILL_0_DFFPOSX1_899 ( );
FILL FILL_1_DFFPOSX1_899 ( );
FILL FILL_2_DFFPOSX1_899 ( );
FILL FILL_3_DFFPOSX1_899 ( );
FILL FILL_4_DFFPOSX1_899 ( );
FILL FILL_5_DFFPOSX1_899 ( );
FILL FILL_0_BUFX4_14 ( );
FILL FILL_1_BUFX4_14 ( );
FILL FILL_2_BUFX4_14 ( );
FILL FILL_0_BUFX4_92 ( );
FILL FILL_1_BUFX4_92 ( );
FILL FILL_2_BUFX4_92 ( );
FILL FILL_0_INVX1_192 ( );
FILL FILL_0_NAND3X1_56 ( );
FILL FILL_1_NAND3X1_56 ( );
FILL FILL_0_AND2X2_29 ( );
FILL FILL_1_AND2X2_29 ( );
FILL FILL_0_NAND3X1_55 ( );
FILL FILL_1_NAND3X1_55 ( );
FILL FILL_0_OAI21X1_1298 ( );
FILL FILL_1_OAI21X1_1298 ( );
FILL FILL_0_NOR2X1_196 ( );
FILL FILL_0_OAI21X1_1300 ( );
FILL FILL_1_OAI21X1_1300 ( );
FILL FILL_0_OAI21X1_1301 ( );
FILL FILL_1_OAI21X1_1301 ( );
FILL FILL_2_OAI21X1_1301 ( );
FILL FILL_0_DFFPOSX1_980 ( );
FILL FILL_1_DFFPOSX1_980 ( );
FILL FILL_2_DFFPOSX1_980 ( );
FILL FILL_3_DFFPOSX1_980 ( );
FILL FILL_4_DFFPOSX1_980 ( );
FILL FILL_5_DFFPOSX1_980 ( );
FILL FILL_6_DFFPOSX1_980 ( );
FILL FILL_0_XNOR2X1_72 ( );
FILL FILL_1_XNOR2X1_72 ( );
FILL FILL_2_XNOR2X1_72 ( );
FILL FILL_3_XNOR2X1_72 ( );
FILL FILL_0_BUFX4_310 ( );
FILL FILL_1_BUFX4_310 ( );
FILL FILL_0_BUFX2_168 ( );
FILL FILL_0_OAI21X1_1519 ( );
FILL FILL_1_OAI21X1_1519 ( );
FILL FILL_2_OAI21X1_1519 ( );
FILL FILL_0_DFFPOSX1_852 ( );
FILL FILL_1_DFFPOSX1_852 ( );
FILL FILL_2_DFFPOSX1_852 ( );
FILL FILL_3_DFFPOSX1_852 ( );
FILL FILL_4_DFFPOSX1_852 ( );
FILL FILL_5_DFFPOSX1_852 ( );
FILL FILL_6_DFFPOSX1_852 ( );
FILL FILL_0_CLKBUF1_36 ( );
FILL FILL_1_CLKBUF1_36 ( );
FILL FILL_2_CLKBUF1_36 ( );
FILL FILL_3_CLKBUF1_36 ( );
FILL FILL_0_BUFX4_87 ( );
FILL FILL_1_BUFX4_87 ( );
FILL FILL_0_NOR2X1_226 ( );
FILL FILL_1_NOR2X1_226 ( );
FILL FILL_0_OAI21X1_1522 ( );
FILL FILL_1_OAI21X1_1522 ( );
FILL FILL_0_NAND2X1_640 ( );
FILL FILL_0_INVX2_102 ( );
FILL FILL_1_INVX2_102 ( );
FILL FILL_0_INVX1_178 ( );
FILL FILL_0_NAND2X1_641 ( );
FILL FILL_1_NAND2X1_641 ( );
FILL FILL_0_BUFX4_45 ( );
FILL FILL_1_BUFX4_45 ( );
FILL FILL_0_OAI21X1_1529 ( );
FILL FILL_1_OAI21X1_1529 ( );
FILL FILL_0_OAI21X1_1530 ( );
FILL FILL_1_OAI21X1_1530 ( );
FILL FILL_0_DFFPOSX1_984 ( );
FILL FILL_1_DFFPOSX1_984 ( );
FILL FILL_2_DFFPOSX1_984 ( );
FILL FILL_3_DFFPOSX1_984 ( );
FILL FILL_4_DFFPOSX1_984 ( );
FILL FILL_5_DFFPOSX1_984 ( );
FILL FILL_6_DFFPOSX1_984 ( );
FILL FILL_0_DFFPOSX1_934 ( );
FILL FILL_1_DFFPOSX1_934 ( );
FILL FILL_2_DFFPOSX1_934 ( );
FILL FILL_3_DFFPOSX1_934 ( );
FILL FILL_4_DFFPOSX1_934 ( );
FILL FILL_5_DFFPOSX1_934 ( );
FILL FILL_6_DFFPOSX1_934 ( );
FILL FILL_0_OAI21X1_1379 ( );
FILL FILL_1_OAI21X1_1379 ( );
FILL FILL_0_CLKBUF1_97 ( );
FILL FILL_1_CLKBUF1_97 ( );
FILL FILL_2_CLKBUF1_97 ( );
FILL FILL_3_CLKBUF1_97 ( );
FILL FILL_4_CLKBUF1_97 ( );
FILL FILL_0_BUFX2_170 ( );
FILL FILL_0_BUFX2_236 ( );
FILL FILL_1_BUFX2_236 ( );
FILL FILL_0_OAI21X1_1082 ( );
FILL FILL_1_OAI21X1_1082 ( );
FILL FILL_0_NAND2X1_448 ( );
FILL FILL_1_NAND2X1_448 ( );
FILL FILL_0_OAI21X1_1099 ( );
FILL FILL_1_OAI21X1_1099 ( );
FILL FILL_0_NAND2X1_465 ( );
FILL FILL_1_NAND2X1_465 ( );
FILL FILL_0_DFFPOSX1_807 ( );
FILL FILL_1_DFFPOSX1_807 ( );
FILL FILL_2_DFFPOSX1_807 ( );
FILL FILL_3_DFFPOSX1_807 ( );
FILL FILL_4_DFFPOSX1_807 ( );
FILL FILL_5_DFFPOSX1_807 ( );
FILL FILL_0_BUFX2_61 ( );
FILL FILL_0_BUFX2_186 ( );
FILL FILL_0_BUFX2_188 ( );
FILL FILL_1_BUFX2_188 ( );
FILL FILL_0_CLKBUF1_26 ( );
FILL FILL_1_CLKBUF1_26 ( );
FILL FILL_2_CLKBUF1_26 ( );
FILL FILL_3_CLKBUF1_26 ( );
FILL FILL_4_CLKBUF1_26 ( );
FILL FILL_0_DFFPOSX1_215 ( );
FILL FILL_1_DFFPOSX1_215 ( );
FILL FILL_2_DFFPOSX1_215 ( );
FILL FILL_3_DFFPOSX1_215 ( );
FILL FILL_4_DFFPOSX1_215 ( );
FILL FILL_5_DFFPOSX1_215 ( );
FILL FILL_6_DFFPOSX1_215 ( );
FILL FILL_0_OAI21X1_59 ( );
FILL FILL_1_OAI21X1_59 ( );
FILL FILL_0_OAI21X1_1825 ( );
FILL FILL_1_OAI21X1_1825 ( );
FILL FILL_0_NAND2X1_766 ( );
FILL FILL_0_DFFPOSX1_151 ( );
FILL FILL_1_DFFPOSX1_151 ( );
FILL FILL_2_DFFPOSX1_151 ( );
FILL FILL_3_DFFPOSX1_151 ( );
FILL FILL_4_DFFPOSX1_151 ( );
FILL FILL_5_DFFPOSX1_151 ( );
FILL FILL_0_BUFX2_984 ( );
FILL FILL_0_NAND2X1_376 ( );
FILL FILL_0_DFFPOSX1_727 ( );
FILL FILL_1_DFFPOSX1_727 ( );
FILL FILL_2_DFFPOSX1_727 ( );
FILL FILL_3_DFFPOSX1_727 ( );
FILL FILL_4_DFFPOSX1_727 ( );
FILL FILL_5_DFFPOSX1_727 ( );
FILL FILL_0_BUFX2_298 ( );
FILL FILL_0_INVX2_195 ( );
FILL FILL_0_OAI21X1_881 ( );
FILL FILL_1_OAI21X1_881 ( );
FILL FILL_2_OAI21X1_881 ( );
FILL FILL_0_BUFX2_723 ( );
FILL FILL_1_BUFX2_723 ( );
FILL FILL_0_BUFX2_691 ( );
FILL FILL_1_BUFX2_691 ( );
FILL FILL_0_INVX2_135 ( );
FILL FILL_0_BUFX2_659 ( );
FILL FILL_0_BUFX2_501 ( );
FILL FILL_0_NAND2X1_700 ( );
FILL FILL_0_DFFPOSX1_54 ( );
FILL FILL_1_DFFPOSX1_54 ( );
FILL FILL_2_DFFPOSX1_54 ( );
FILL FILL_3_DFFPOSX1_54 ( );
FILL FILL_4_DFFPOSX1_54 ( );
FILL FILL_5_DFFPOSX1_54 ( );
FILL FILL_0_OAI21X1_1682 ( );
FILL FILL_1_OAI21X1_1682 ( );
FILL FILL_0_OAI21X1_1683 ( );
FILL FILL_1_OAI21X1_1683 ( );
FILL FILL_0_NAND2X1_668 ( );
FILL FILL_0_OAI21X1_1210 ( );
FILL FILL_1_OAI21X1_1210 ( );
FILL FILL_2_OAI21X1_1210 ( );
FILL FILL_0_OAI21X1_1211 ( );
FILL FILL_1_OAI21X1_1211 ( );
FILL FILL_0_DFFPOSX1_873 ( );
FILL FILL_1_DFFPOSX1_873 ( );
FILL FILL_2_DFFPOSX1_873 ( );
FILL FILL_3_DFFPOSX1_873 ( );
FILL FILL_4_DFFPOSX1_873 ( );
FILL FILL_5_DFFPOSX1_873 ( );
FILL FILL_0_BUFX2_373 ( );
FILL FILL_0_CLKBUF1_78 ( );
FILL FILL_1_CLKBUF1_78 ( );
FILL FILL_2_CLKBUF1_78 ( );
FILL FILL_3_CLKBUF1_78 ( );
FILL FILL_4_CLKBUF1_78 ( );
FILL FILL_0_BUFX4_125 ( );
FILL FILL_1_BUFX4_125 ( );
FILL FILL_0_BUFX4_83 ( );
FILL FILL_1_BUFX4_83 ( );
FILL FILL_0_DFFPOSX1_469 ( );
FILL FILL_1_DFFPOSX1_469 ( );
FILL FILL_2_DFFPOSX1_469 ( );
FILL FILL_3_DFFPOSX1_469 ( );
FILL FILL_4_DFFPOSX1_469 ( );
FILL FILL_5_DFFPOSX1_469 ( );
FILL FILL_0_NAND2X1_237 ( );
FILL FILL_1_NAND2X1_237 ( );
FILL FILL_0_BUFX2_592 ( );
FILL FILL_0_OAI21X1_1702 ( );
FILL FILL_1_OAI21X1_1702 ( );
FILL FILL_0_BUFX4_85 ( );
FILL FILL_1_BUFX4_85 ( );
FILL FILL_2_BUFX4_85 ( );
FILL FILL_0_DFFPOSX1_563 ( );
FILL FILL_1_DFFPOSX1_563 ( );
FILL FILL_2_DFFPOSX1_563 ( );
FILL FILL_3_DFFPOSX1_563 ( );
FILL FILL_4_DFFPOSX1_563 ( );
FILL FILL_5_DFFPOSX1_563 ( );
FILL FILL_0_OAI21X1_702 ( );
FILL FILL_1_OAI21X1_702 ( );
FILL FILL_0_OAI21X1_703 ( );
FILL FILL_1_OAI21X1_703 ( );
FILL FILL_0_OAI21X1_1411 ( );
FILL FILL_1_OAI21X1_1411 ( );
FILL FILL_0_BUFX4_24 ( );
FILL FILL_1_BUFX4_24 ( );
FILL FILL_0_BUFX2_631 ( );
FILL FILL_0_BUFX4_323 ( );
FILL FILL_1_BUFX4_323 ( );
FILL FILL_0_OAI21X1_629 ( );
FILL FILL_1_OAI21X1_629 ( );
FILL FILL_0_OAI21X1_605 ( );
FILL FILL_1_OAI21X1_605 ( );
FILL FILL_0_OAI21X1_606 ( );
FILL FILL_1_OAI21X1_606 ( );
FILL FILL_0_DFFPOSX1_598 ( );
FILL FILL_1_DFFPOSX1_598 ( );
FILL FILL_2_DFFPOSX1_598 ( );
FILL FILL_3_DFFPOSX1_598 ( );
FILL FILL_4_DFFPOSX1_598 ( );
FILL FILL_5_DFFPOSX1_598 ( );
FILL FILL_6_DFFPOSX1_598 ( );
FILL FILL_0_OAI21X1_804 ( );
FILL FILL_1_OAI21X1_804 ( );
FILL FILL_2_OAI21X1_804 ( );
FILL FILL_0_OAI21X1_805 ( );
FILL FILL_1_OAI21X1_805 ( );
FILL FILL_0_BUFX2_500 ( );
FILL FILL_1_BUFX2_500 ( );
FILL FILL_0_DFFPOSX1_468 ( );
FILL FILL_1_DFFPOSX1_468 ( );
FILL FILL_2_DFFPOSX1_468 ( );
FILL FILL_3_DFFPOSX1_468 ( );
FILL FILL_4_DFFPOSX1_468 ( );
FILL FILL_5_DFFPOSX1_468 ( );
FILL FILL_6_DFFPOSX1_468 ( );
FILL FILL_0_OAI21X1_802 ( );
FILL FILL_1_OAI21X1_802 ( );
FILL FILL_0_OAI21X1_803 ( );
FILL FILL_1_OAI21X1_803 ( );
FILL FILL_0_NOR2X1_46 ( );
FILL FILL_1_NOR2X1_46 ( );
FILL FILL_0_NOR2X1_94 ( );
FILL FILL_0_INVX2_51 ( );
FILL FILL_0_BUFX2_426 ( );
FILL FILL_1_BUFX2_426 ( );
FILL FILL_0_BUFX4_63 ( );
FILL FILL_1_BUFX4_63 ( );
FILL FILL_0_NAND2X1_299 ( );
FILL FILL_0_NAND2X1_242 ( );
FILL FILL_0_BUFX4_289 ( );
FILL FILL_1_BUFX4_289 ( );
FILL FILL_0_NOR2X1_97 ( );
FILL FILL_1_NOR2X1_97 ( );
FILL FILL_0_OAI21X1_642 ( );
FILL FILL_1_OAI21X1_642 ( );
FILL FILL_0_NAND2X1_649 ( );
FILL FILL_1_NAND2X1_649 ( );
FILL FILL_0_OAI21X1_1576 ( );
FILL FILL_1_OAI21X1_1576 ( );
FILL FILL_0_XNOR2X1_23 ( );
FILL FILL_1_XNOR2X1_23 ( );
FILL FILL_2_XNOR2X1_23 ( );
FILL FILL_3_XNOR2X1_23 ( );
FILL FILL_0_NAND2X1_213 ( );
FILL FILL_1_NAND2X1_213 ( );
FILL FILL_0_OAI21X1_456 ( );
FILL FILL_1_OAI21X1_456 ( );
FILL FILL_0_XNOR2X1_55 ( );
FILL FILL_1_XNOR2X1_55 ( );
FILL FILL_2_XNOR2X1_55 ( );
FILL FILL_3_XNOR2X1_55 ( );
FILL FILL_0_INVX1_22 ( );
FILL FILL_0_OAI21X1_491 ( );
FILL FILL_1_OAI21X1_491 ( );
FILL FILL_0_NOR2X1_55 ( );
FILL FILL_1_NOR2X1_55 ( );
FILL FILL_0_NAND2X1_333 ( );
FILL FILL_1_NAND2X1_333 ( );
FILL FILL_0_BUFX2_618 ( );
FILL FILL_0_NAND3X1_13 ( );
FILL FILL_1_NAND3X1_13 ( );
FILL FILL_0_NAND3X1_12 ( );
FILL FILL_1_NAND3X1_12 ( );
FILL FILL_0_OAI21X1_497 ( );
FILL FILL_1_OAI21X1_497 ( );
FILL FILL_0_OAI21X1_495 ( );
FILL FILL_1_OAI21X1_495 ( );
FILL FILL_2_OAI21X1_495 ( );
FILL FILL_0_OAI21X1_496 ( );
FILL FILL_1_OAI21X1_496 ( );
FILL FILL_0_NAND2X1_261 ( );
FILL FILL_1_NAND2X1_261 ( );
FILL FILL_0_DFFPOSX1_481 ( );
FILL FILL_1_DFFPOSX1_481 ( );
FILL FILL_2_DFFPOSX1_481 ( );
FILL FILL_3_DFFPOSX1_481 ( );
FILL FILL_4_DFFPOSX1_481 ( );
FILL FILL_5_DFFPOSX1_481 ( );
FILL FILL_6_DFFPOSX1_481 ( );
FILL FILL_0_DFFPOSX1_607 ( );
FILL FILL_1_DFFPOSX1_607 ( );
FILL FILL_2_DFFPOSX1_607 ( );
FILL FILL_3_DFFPOSX1_607 ( );
FILL FILL_4_DFFPOSX1_607 ( );
FILL FILL_5_DFFPOSX1_607 ( );
FILL FILL_6_DFFPOSX1_607 ( );
FILL FILL_0_OAI21X1_826 ( );
FILL FILL_1_OAI21X1_826 ( );
FILL FILL_0_DFFPOSX1_605 ( );
FILL FILL_1_DFFPOSX1_605 ( );
FILL FILL_2_DFFPOSX1_605 ( );
FILL FILL_3_DFFPOSX1_605 ( );
FILL FILL_4_DFFPOSX1_605 ( );
FILL FILL_5_DFFPOSX1_605 ( );
FILL FILL_6_DFFPOSX1_605 ( );
FILL FILL_0_BUFX2_532 ( );
FILL FILL_0_BUFX4_77 ( );
FILL FILL_1_BUFX4_77 ( );
FILL FILL_0_NAND2X1_176 ( );
FILL FILL_0_OAI21X1_715 ( );
FILL FILL_1_OAI21X1_715 ( );
FILL FILL_0_OAI21X1_429 ( );
FILL FILL_1_OAI21X1_429 ( );
FILL FILL_0_DFFPOSX1_456 ( );
FILL FILL_1_DFFPOSX1_456 ( );
FILL FILL_2_DFFPOSX1_456 ( );
FILL FILL_3_DFFPOSX1_456 ( );
FILL FILL_4_DFFPOSX1_456 ( );
FILL FILL_5_DFFPOSX1_456 ( );
FILL FILL_0_BUFX2_840 ( );
FILL FILL_1_BUFX2_840 ( );
FILL FILL_0_OAI21X1_1783 ( );
FILL FILL_1_OAI21X1_1783 ( );
FILL FILL_0_NAND2X1_724 ( );
FILL FILL_1_NAND2X1_724 ( );
FILL FILL_0_OAI21X1_824 ( );
FILL FILL_1_OAI21X1_824 ( );
FILL FILL_0_DFFPOSX1_604 ( );
FILL FILL_1_DFFPOSX1_604 ( );
FILL FILL_2_DFFPOSX1_604 ( );
FILL FILL_3_DFFPOSX1_604 ( );
FILL FILL_4_DFFPOSX1_604 ( );
FILL FILL_5_DFFPOSX1_604 ( );
FILL FILL_0_OAI21X1_745 ( );
FILL FILL_1_OAI21X1_745 ( );
FILL FILL_2_OAI21X1_745 ( );
FILL FILL_0_BUFX2_411 ( );
FILL FILL_1_BUFX2_411 ( );
FILL FILL_0_NAND2X1_200 ( );
FILL FILL_1_NAND2X1_200 ( );
FILL FILL_0_DFFPOSX1_61 ( );
FILL FILL_1_DFFPOSX1_61 ( );
FILL FILL_2_DFFPOSX1_61 ( );
FILL FILL_3_DFFPOSX1_61 ( );
FILL FILL_4_DFFPOSX1_61 ( );
FILL FILL_5_DFFPOSX1_61 ( );
FILL FILL_6_DFFPOSX1_61 ( );
FILL FILL_0_OAI21X1_1696 ( );
FILL FILL_1_OAI21X1_1696 ( );
FILL FILL_0_NAND2X1_189 ( );
FILL FILL_1_NAND2X1_189 ( );
FILL FILL_0_DFFPOSX1_29 ( );
FILL FILL_1_DFFPOSX1_29 ( );
FILL FILL_2_DFFPOSX1_29 ( );
FILL FILL_3_DFFPOSX1_29 ( );
FILL FILL_4_DFFPOSX1_29 ( );
FILL FILL_5_DFFPOSX1_29 ( );
FILL FILL_6_DFFPOSX1_29 ( );
FILL FILL_0_OAI21X1_314 ( );
FILL FILL_1_OAI21X1_314 ( );
FILL FILL_0_NAND2X1_420 ( );
FILL FILL_1_NAND2X1_420 ( );
FILL FILL_0_OAI21X1_1054 ( );
FILL FILL_1_OAI21X1_1054 ( );
FILL FILL_0_BUFX4_95 ( );
FILL FILL_1_BUFX4_95 ( );
FILL FILL_0_BUFX4_109 ( );
FILL FILL_1_BUFX4_109 ( );
FILL FILL_0_BUFX4_104 ( );
FILL FILL_1_BUFX4_104 ( );
FILL FILL_0_CLKBUF1_55 ( );
FILL FILL_1_CLKBUF1_55 ( );
FILL FILL_2_CLKBUF1_55 ( );
FILL FILL_3_CLKBUF1_55 ( );
FILL FILL_4_CLKBUF1_55 ( );
FILL FILL_0_NAND2X1_603 ( );
FILL FILL_0_OAI21X1_1458 ( );
FILL FILL_1_OAI21X1_1458 ( );
FILL FILL_0_NOR2X1_224 ( );
FILL FILL_1_NOR2X1_224 ( );
FILL FILL_0_NOR2X1_144 ( );
FILL FILL_0_NAND2X1_523 ( );
FILL FILL_1_NAND2X1_523 ( );
FILL FILL_0_NOR2X1_194 ( );
FILL FILL_1_NOR2X1_194 ( );
FILL FILL_0_NOR2X1_195 ( );
FILL FILL_1_NOR2X1_195 ( );
FILL FILL_0_OAI21X1_1287 ( );
FILL FILL_1_OAI21X1_1287 ( );
FILL FILL_0_NAND3X1_40 ( );
FILL FILL_1_NAND3X1_40 ( );
FILL FILL_0_OAI21X1_122 ( );
FILL FILL_1_OAI21X1_122 ( );
FILL FILL_0_BUFX2_907 ( );
FILL FILL_1_BUFX2_907 ( );
FILL FILL_0_INVX2_109 ( );
FILL FILL_1_INVX2_109 ( );
FILL FILL_0_NAND3X1_64 ( );
FILL FILL_1_NAND3X1_64 ( );
FILL FILL_0_NOR2X1_151 ( );
FILL FILL_1_NOR2X1_151 ( );
FILL FILL_0_INVX1_189 ( );
FILL FILL_0_NAND2X1_520 ( );
FILL FILL_1_NAND2X1_520 ( );
FILL FILL_0_BUFX2_935 ( );
FILL FILL_0_CLKBUF1_49 ( );
FILL FILL_1_CLKBUF1_49 ( );
FILL FILL_2_CLKBUF1_49 ( );
FILL FILL_3_CLKBUF1_49 ( );
FILL FILL_0_BUFX2_149 ( );
FILL FILL_1_BUFX2_149 ( );
FILL FILL_0_DFFPOSX1_905 ( );
FILL FILL_1_DFFPOSX1_905 ( );
FILL FILL_2_DFFPOSX1_905 ( );
FILL FILL_3_DFFPOSX1_905 ( );
FILL FILL_4_DFFPOSX1_905 ( );
FILL FILL_5_DFFPOSX1_905 ( );
FILL FILL_0_OAI21X1_1297 ( );
FILL FILL_1_OAI21X1_1297 ( );
FILL FILL_0_OAI21X1_1299 ( );
FILL FILL_1_OAI21X1_1299 ( );
FILL FILL_2_OAI21X1_1299 ( );
FILL FILL_0_AND2X2_30 ( );
FILL FILL_1_AND2X2_30 ( );
FILL FILL_0_OAI21X1_1461 ( );
FILL FILL_1_OAI21X1_1461 ( );
FILL FILL_0_CLKBUF1_68 ( );
FILL FILL_1_CLKBUF1_68 ( );
FILL FILL_2_CLKBUF1_68 ( );
FILL FILL_3_CLKBUF1_68 ( );
FILL FILL_4_CLKBUF1_68 ( );
FILL FILL_0_NAND2X1_607 ( );
FILL FILL_1_NAND2X1_607 ( );
FILL FILL_0_OAI21X1_1515 ( );
FILL FILL_1_OAI21X1_1515 ( );
FILL FILL_0_INVX1_177 ( );
FILL FILL_1_INVX1_177 ( );
FILL FILL_0_OAI21X1_1171 ( );
FILL FILL_1_OAI21X1_1171 ( );
FILL FILL_0_NAND2X1_554 ( );
FILL FILL_0_XNOR2X1_73 ( );
FILL FILL_1_XNOR2X1_73 ( );
FILL FILL_2_XNOR2X1_73 ( );
FILL FILL_3_XNOR2X1_73 ( );
FILL FILL_0_NOR2X1_161 ( );
FILL FILL_1_NOR2X1_161 ( );
FILL FILL_0_OAI21X1_1172 ( );
FILL FILL_1_OAI21X1_1172 ( );
FILL FILL_2_OAI21X1_1172 ( );
FILL FILL_0_NAND2X1_636 ( );
FILL FILL_0_OAI21X1_1482 ( );
FILL FILL_1_OAI21X1_1482 ( );
FILL FILL_0_OAI21X1_1480 ( );
FILL FILL_1_OAI21X1_1480 ( );
FILL FILL_0_DFFPOSX1_969 ( );
FILL FILL_1_DFFPOSX1_969 ( );
FILL FILL_2_DFFPOSX1_969 ( );
FILL FILL_3_DFFPOSX1_969 ( );
FILL FILL_4_DFFPOSX1_969 ( );
FILL FILL_5_DFFPOSX1_969 ( );
FILL FILL_6_DFFPOSX1_969 ( );
FILL FILL_0_BUFX2_220 ( );
FILL FILL_0_DFFPOSX1_982 ( );
FILL FILL_1_DFFPOSX1_982 ( );
FILL FILL_2_DFFPOSX1_982 ( );
FILL FILL_3_DFFPOSX1_982 ( );
FILL FILL_4_DFFPOSX1_982 ( );
FILL FILL_5_DFFPOSX1_982 ( );
FILL FILL_6_DFFPOSX1_982 ( );
FILL FILL_0_OAI21X1_1524 ( );
FILL FILL_1_OAI21X1_1524 ( );
FILL FILL_0_OAI21X1_1523 ( );
FILL FILL_1_OAI21X1_1523 ( );
FILL FILL_0_INVX1_225 ( );
FILL FILL_0_AOI21X1_62 ( );
FILL FILL_1_AOI21X1_62 ( );
FILL FILL_0_NOR2X1_227 ( );
FILL FILL_1_NOR2X1_227 ( );
FILL FILL_0_OAI21X1_1526 ( );
FILL FILL_1_OAI21X1_1526 ( );
FILL FILL_0_OAI21X1_1527 ( );
FILL FILL_1_OAI21X1_1527 ( );
FILL FILL_0_OAI21X1_1525 ( );
FILL FILL_1_OAI21X1_1525 ( );
FILL FILL_0_DFFPOSX1_983 ( );
FILL FILL_1_DFFPOSX1_983 ( );
FILL FILL_2_DFFPOSX1_983 ( );
FILL FILL_3_DFFPOSX1_983 ( );
FILL FILL_4_DFFPOSX1_983 ( );
FILL FILL_5_DFFPOSX1_983 ( );
FILL FILL_0_OAI21X1_1521 ( );
FILL FILL_1_OAI21X1_1521 ( );
FILL FILL_0_DFFPOSX1_981 ( );
FILL FILL_1_DFFPOSX1_981 ( );
FILL FILL_2_DFFPOSX1_981 ( );
FILL FILL_3_DFFPOSX1_981 ( );
FILL FILL_4_DFFPOSX1_981 ( );
FILL FILL_5_DFFPOSX1_981 ( );
FILL FILL_0_DFFPOSX1_790 ( );
FILL FILL_1_DFFPOSX1_790 ( );
FILL FILL_2_DFFPOSX1_790 ( );
FILL FILL_3_DFFPOSX1_790 ( );
FILL FILL_4_DFFPOSX1_790 ( );
FILL FILL_5_DFFPOSX1_790 ( );
FILL FILL_0_OAI21X1_1572 ( );
FILL FILL_1_OAI21X1_1572 ( );
FILL FILL_0_OAI21X1_1098 ( );
FILL FILL_1_OAI21X1_1098 ( );
FILL FILL_2_OAI21X1_1098 ( );
FILL FILL_0_OAI21X1_26 ( );
FILL FILL_1_OAI21X1_26 ( );
FILL FILL_0_DFFPOSX1_182 ( );
FILL FILL_1_DFFPOSX1_182 ( );
FILL FILL_2_DFFPOSX1_182 ( );
FILL FILL_3_DFFPOSX1_182 ( );
FILL FILL_4_DFFPOSX1_182 ( );
FILL FILL_5_DFFPOSX1_182 ( );
FILL FILL_6_DFFPOSX1_182 ( );
FILL FILL_0_OAI21X1_279 ( );
FILL FILL_1_OAI21X1_279 ( );
FILL FILL_2_OAI21X1_279 ( );
FILL FILL_0_DFFPOSX1_331 ( );
FILL FILL_1_DFFPOSX1_331 ( );
FILL FILL_2_DFFPOSX1_331 ( );
FILL FILL_3_DFFPOSX1_331 ( );
FILL FILL_4_DFFPOSX1_331 ( );
FILL FILL_5_DFFPOSX1_331 ( );
FILL FILL_0_NAND2X1_26 ( );
FILL FILL_1_NAND2X1_26 ( );
FILL FILL_0_NAND2X1_59 ( );
FILL FILL_0_DFFPOSX1_170 ( );
FILL FILL_1_DFFPOSX1_170 ( );
FILL FILL_2_DFFPOSX1_170 ( );
FILL FILL_3_DFFPOSX1_170 ( );
FILL FILL_4_DFFPOSX1_170 ( );
FILL FILL_5_DFFPOSX1_170 ( );
FILL FILL_0_OAI21X1_14 ( );
FILL FILL_1_OAI21X1_14 ( );
FILL FILL_0_BUFX2_851 ( );
FILL FILL_1_BUFX2_851 ( );
FILL FILL_0_DFFPOSX1_171 ( );
FILL FILL_1_DFFPOSX1_171 ( );
FILL FILL_2_DFFPOSX1_171 ( );
FILL FILL_3_DFFPOSX1_171 ( );
FILL FILL_4_DFFPOSX1_171 ( );
FILL FILL_5_DFFPOSX1_171 ( );
FILL FILL_0_OAI21X1_15 ( );
FILL FILL_1_OAI21X1_15 ( );
FILL FILL_2_OAI21X1_15 ( );
FILL FILL_0_NAND2X1_15 ( );
FILL FILL_0_BUFX2_902 ( );
FILL FILL_1_BUFX2_902 ( );
FILL FILL_0_BUFX2_824 ( );
FILL FILL_1_BUFX2_824 ( );
FILL FILL_0_INVX2_55 ( );
FILL FILL_0_BUFX2_930 ( );
FILL FILL_0_BUFX2_866 ( );
FILL FILL_1_BUFX2_866 ( );
FILL FILL_0_BUFX4_263 ( );
FILL FILL_1_BUFX4_263 ( );
FILL FILL_0_NAND2X1_39 ( );
FILL FILL_1_NAND2X1_39 ( );
FILL FILL_0_OAI21X1_1101 ( );
FILL FILL_1_OAI21X1_1101 ( );
FILL FILL_2_OAI21X1_1101 ( );
FILL FILL_0_NAND2X1_467 ( );
FILL FILL_0_DFFPOSX1_809 ( );
FILL FILL_1_DFFPOSX1_809 ( );
FILL FILL_2_DFFPOSX1_809 ( );
FILL FILL_3_DFFPOSX1_809 ( );
FILL FILL_4_DFFPOSX1_809 ( );
FILL FILL_5_DFFPOSX1_809 ( );
FILL FILL_6_DFFPOSX1_809 ( );
FILL FILL_0_BUFX2_130 ( );
FILL FILL_1_BUFX2_130 ( );
FILL FILL_0_BUFX4_230 ( );
FILL FILL_1_BUFX4_230 ( );
FILL FILL_0_OAI21X1_134 ( );
FILL FILL_1_OAI21X1_134 ( );
FILL FILL_0_OAI21X1_135 ( );
FILL FILL_1_OAI21X1_135 ( );
FILL FILL_0_DFFPOSX1_259 ( );
FILL FILL_1_DFFPOSX1_259 ( );
FILL FILL_2_DFFPOSX1_259 ( );
FILL FILL_3_DFFPOSX1_259 ( );
FILL FILL_4_DFFPOSX1_259 ( );
FILL FILL_5_DFFPOSX1_259 ( );
FILL FILL_0_DFFPOSX1_729 ( );
FILL FILL_1_DFFPOSX1_729 ( );
FILL FILL_2_DFFPOSX1_729 ( );
FILL FILL_3_DFFPOSX1_729 ( );
FILL FILL_4_DFFPOSX1_729 ( );
FILL FILL_5_DFFPOSX1_729 ( );
FILL FILL_0_DFFPOSX1_313 ( );
FILL FILL_1_DFFPOSX1_313 ( );
FILL FILL_2_DFFPOSX1_313 ( );
FILL FILL_3_DFFPOSX1_313 ( );
FILL FILL_4_DFFPOSX1_313 ( );
FILL FILL_5_DFFPOSX1_313 ( );
FILL FILL_0_OAI21X1_243 ( );
FILL FILL_1_OAI21X1_243 ( );
FILL FILL_0_OAI21X1_242 ( );
FILL FILL_1_OAI21X1_242 ( );
FILL FILL_0_OAI21X1_1703 ( );
FILL FILL_1_OAI21X1_1703 ( );
FILL FILL_0_DFFPOSX1_64 ( );
FILL FILL_1_DFFPOSX1_64 ( );
FILL FILL_2_DFFPOSX1_64 ( );
FILL FILL_3_DFFPOSX1_64 ( );
FILL FILL_4_DFFPOSX1_64 ( );
FILL FILL_5_DFFPOSX1_64 ( );
FILL FILL_0_BUFX4_179 ( );
FILL FILL_1_BUFX4_179 ( );
FILL FILL_0_CLKBUF1_22 ( );
FILL FILL_1_CLKBUF1_22 ( );
FILL FILL_2_CLKBUF1_22 ( );
FILL FILL_3_CLKBUF1_22 ( );
FILL FILL_4_CLKBUF1_22 ( );
FILL FILL_0_DFFPOSX1_945 ( );
FILL FILL_1_DFFPOSX1_945 ( );
FILL FILL_2_DFFPOSX1_945 ( );
FILL FILL_3_DFFPOSX1_945 ( );
FILL FILL_4_DFFPOSX1_945 ( );
FILL FILL_5_DFFPOSX1_945 ( );
FILL FILL_6_DFFPOSX1_945 ( );
FILL FILL_0_OAI21X1_1412 ( );
FILL FILL_1_OAI21X1_1412 ( );
FILL FILL_0_DFFPOSX1_525 ( );
FILL FILL_1_DFFPOSX1_525 ( );
FILL FILL_2_DFFPOSX1_525 ( );
FILL FILL_3_DFFPOSX1_525 ( );
FILL FILL_4_DFFPOSX1_525 ( );
FILL FILL_5_DFFPOSX1_525 ( );
FILL FILL_6_DFFPOSX1_525 ( );
FILL FILL_0_NAND2X1_121 ( );
FILL FILL_1_NAND2X1_121 ( );
FILL FILL_0_OAI21X1_377 ( );
FILL FILL_1_OAI21X1_377 ( );
FILL FILL_0_NOR2X1_92 ( );
FILL FILL_1_NOR2X1_92 ( );
FILL FILL_0_DFFPOSX1_470 ( );
FILL FILL_1_DFFPOSX1_470 ( );
FILL FILL_2_DFFPOSX1_470 ( );
FILL FILL_3_DFFPOSX1_470 ( );
FILL FILL_4_DFFPOSX1_470 ( );
FILL FILL_5_DFFPOSX1_470 ( );
FILL FILL_0_NAND2X1_239 ( );
FILL FILL_1_NAND2X1_239 ( );
FILL FILL_0_OAI21X1_477 ( );
FILL FILL_1_OAI21X1_477 ( );
FILL FILL_0_NOR2X1_45 ( );
FILL FILL_1_NOR2X1_45 ( );
FILL FILL_0_OAI21X1_476 ( );
FILL FILL_1_OAI21X1_476 ( );
FILL FILL_0_NAND2X1_238 ( );
FILL FILL_1_NAND2X1_238 ( );
FILL FILL_0_NOR2X1_44 ( );
FILL FILL_0_OAI21X1_627 ( );
FILL FILL_1_OAI21X1_627 ( );
FILL FILL_2_OAI21X1_627 ( );
FILL FILL_0_BUFX4_107 ( );
FILL FILL_1_BUFX4_107 ( );
FILL FILL_0_CLKBUF1_72 ( );
FILL FILL_1_CLKBUF1_72 ( );
FILL FILL_2_CLKBUF1_72 ( );
FILL FILL_3_CLKBUF1_72 ( );
FILL FILL_4_CLKBUF1_72 ( );
FILL FILL_0_DFFPOSX1_599 ( );
FILL FILL_1_DFFPOSX1_599 ( );
FILL FILL_2_DFFPOSX1_599 ( );
FILL FILL_3_DFFPOSX1_599 ( );
FILL FILL_4_DFFPOSX1_599 ( );
FILL FILL_5_DFFPOSX1_599 ( );
FILL FILL_0_OAI21X1_809 ( );
FILL FILL_1_OAI21X1_809 ( );
FILL FILL_0_OAI21X1_808 ( );
FILL FILL_1_OAI21X1_808 ( );
FILL FILL_0_DFFPOSX1_1001 ( );
FILL FILL_1_DFFPOSX1_1001 ( );
FILL FILL_2_DFFPOSX1_1001 ( );
FILL FILL_3_DFFPOSX1_1001 ( );
FILL FILL_4_DFFPOSX1_1001 ( );
FILL FILL_5_DFFPOSX1_1001 ( );
FILL FILL_6_DFFPOSX1_1001 ( );
FILL FILL_0_DFFPOSX1_458 ( );
FILL FILL_1_DFFPOSX1_458 ( );
FILL FILL_2_DFFPOSX1_458 ( );
FILL FILL_3_DFFPOSX1_458 ( );
FILL FILL_4_DFFPOSX1_458 ( );
FILL FILL_5_DFFPOSX1_458 ( );
FILL FILL_6_DFFPOSX1_458 ( );
FILL FILL_0_NAND2X1_257 ( );
FILL FILL_0_OAI21X1_827 ( );
FILL FILL_1_OAI21X1_827 ( );
FILL FILL_0_OAI21X1_828 ( );
FILL FILL_1_OAI21X1_828 ( );
FILL FILL_0_NOR2X1_116 ( );
FILL FILL_0_INVX1_43 ( );
FILL FILL_0_NOR2X1_117 ( );
FILL FILL_1_NOR2X1_117 ( );
FILL FILL_0_DFFPOSX1_610 ( );
FILL FILL_1_DFFPOSX1_610 ( );
FILL FILL_2_DFFPOSX1_610 ( );
FILL FILL_3_DFFPOSX1_610 ( );
FILL FILL_4_DFFPOSX1_610 ( );
FILL FILL_5_DFFPOSX1_610 ( );
FILL FILL_0_OAI21X1_840 ( );
FILL FILL_1_OAI21X1_840 ( );
FILL FILL_0_INVX2_38 ( );
FILL FILL_0_NOR2X1_99 ( );
FILL FILL_0_OAI21X1_839 ( );
FILL FILL_1_OAI21X1_839 ( );
FILL FILL_0_NOR2X1_56 ( );
FILL FILL_1_NOR2X1_56 ( );
FILL FILL_0_AOI21X1_6 ( );
FILL FILL_1_AOI21X1_6 ( );
FILL FILL_0_NOR2X1_118 ( );
FILL FILL_0_OAI21X1_498 ( );
FILL FILL_1_OAI21X1_498 ( );
FILL FILL_0_NAND2X1_263 ( );
FILL FILL_0_OAI21X1_758 ( );
FILL FILL_1_OAI21X1_758 ( );
FILL FILL_2_OAI21X1_758 ( );
FILL FILL_0_NAND2X1_334 ( );
FILL FILL_1_NAND2X1_334 ( );
FILL FILL_0_OAI21X1_832 ( );
FILL FILL_1_OAI21X1_832 ( );
FILL FILL_0_OAI21X1_831 ( );
FILL FILL_1_OAI21X1_831 ( );
FILL FILL_0_OAI21X1_825 ( );
FILL FILL_1_OAI21X1_825 ( );
FILL FILL_0_BUFX4_43 ( );
FILL FILL_1_BUFX4_43 ( );
FILL FILL_0_NAND2X1_108 ( );
FILL FILL_0_OAI21X1_364 ( );
FILL FILL_1_OAI21X1_364 ( );
FILL FILL_0_DFFPOSX1_567 ( );
FILL FILL_1_DFFPOSX1_567 ( );
FILL FILL_2_DFFPOSX1_567 ( );
FILL FILL_3_DFFPOSX1_567 ( );
FILL FILL_4_DFFPOSX1_567 ( );
FILL FILL_5_DFFPOSX1_567 ( );
FILL FILL_0_BUFX4_48 ( );
FILL FILL_1_BUFX4_48 ( );
FILL FILL_0_BUFX4_305 ( );
FILL FILL_1_BUFX4_305 ( );
FILL FILL_0_OAI21X1_17 ( );
FILL FILL_1_OAI21X1_17 ( );
FILL FILL_0_DFFPOSX1_173 ( );
FILL FILL_1_DFFPOSX1_173 ( );
FILL FILL_2_DFFPOSX1_173 ( );
FILL FILL_3_DFFPOSX1_173 ( );
FILL FILL_4_DFFPOSX1_173 ( );
FILL FILL_5_DFFPOSX1_173 ( );
FILL FILL_0_OAI21X1_823 ( );
FILL FILL_1_OAI21X1_823 ( );
FILL FILL_0_DFFPOSX1_578 ( );
FILL FILL_1_DFFPOSX1_578 ( );
FILL FILL_2_DFFPOSX1_578 ( );
FILL FILL_3_DFFPOSX1_578 ( );
FILL FILL_4_DFFPOSX1_578 ( );
FILL FILL_5_DFFPOSX1_578 ( );
FILL FILL_0_OAI21X1_232 ( );
FILL FILL_1_OAI21X1_232 ( );
FILL FILL_0_DFFPOSX1_308 ( );
FILL FILL_1_DFFPOSX1_308 ( );
FILL FILL_2_DFFPOSX1_308 ( );
FILL FILL_3_DFFPOSX1_308 ( );
FILL FILL_4_DFFPOSX1_308 ( );
FILL FILL_5_DFFPOSX1_308 ( );
FILL FILL_6_DFFPOSX1_308 ( );
FILL FILL_0_OAI21X1_233 ( );
FILL FILL_1_OAI21X1_233 ( );
FILL FILL_2_OAI21X1_233 ( );
FILL FILL_0_OAI21X1_571 ( );
FILL FILL_1_OAI21X1_571 ( );
FILL FILL_0_OAI21X1_568 ( );
FILL FILL_1_OAI21X1_568 ( );
FILL FILL_0_BUFX2_475 ( );
FILL FILL_0_OAI21X1_105 ( );
FILL FILL_1_OAI21X1_105 ( );
FILL FILL_0_DFFPOSX1_244 ( );
FILL FILL_1_DFFPOSX1_244 ( );
FILL FILL_2_DFFPOSX1_244 ( );
FILL FILL_3_DFFPOSX1_244 ( );
FILL FILL_4_DFFPOSX1_244 ( );
FILL FILL_5_DFFPOSX1_244 ( );
FILL FILL_0_NOR2X1_220 ( );
FILL FILL_1_NOR2X1_220 ( );
FILL FILL_0_OAI21X1_1436 ( );
FILL FILL_1_OAI21X1_1436 ( );
FILL FILL_0_NAND2X1_628 ( );
FILL FILL_0_OAI21X1_315 ( );
FILL FILL_1_OAI21X1_315 ( );
FILL FILL_0_DFFPOSX1_762 ( );
FILL FILL_1_DFFPOSX1_762 ( );
FILL FILL_2_DFFPOSX1_762 ( );
FILL FILL_3_DFFPOSX1_762 ( );
FILL FILL_4_DFFPOSX1_762 ( );
FILL FILL_5_DFFPOSX1_762 ( );
FILL FILL_0_BUFX4_253 ( );
FILL FILL_1_BUFX4_253 ( );
FILL FILL_0_NAND2X1_633 ( );
FILL FILL_1_NAND2X1_633 ( );
FILL FILL_0_NAND2X1_526 ( );
FILL FILL_1_NAND2X1_526 ( );
FILL FILL_0_DFFPOSX1_898 ( );
FILL FILL_1_DFFPOSX1_898 ( );
FILL FILL_2_DFFPOSX1_898 ( );
FILL FILL_3_DFFPOSX1_898 ( );
FILL FILL_4_DFFPOSX1_898 ( );
FILL FILL_5_DFFPOSX1_898 ( );
FILL FILL_0_INVX2_71 ( );
FILL FILL_0_NAND2X1_632 ( );
FILL FILL_0_BUFX4_26 ( );
FILL FILL_1_BUFX4_26 ( );
FILL FILL_0_OAI21X1_123 ( );
FILL FILL_1_OAI21X1_123 ( );
FILL FILL_2_OAI21X1_123 ( );
FILL FILL_0_DFFPOSX1_900 ( );
FILL FILL_1_DFFPOSX1_900 ( );
FILL FILL_2_DFFPOSX1_900 ( );
FILL FILL_3_DFFPOSX1_900 ( );
FILL FILL_4_DFFPOSX1_900 ( );
FILL FILL_5_DFFPOSX1_900 ( );
FILL FILL_6_DFFPOSX1_900 ( );
FILL FILL_0_INVX2_72 ( );
FILL FILL_0_XNOR2X1_98 ( );
FILL FILL_1_XNOR2X1_98 ( );
FILL FILL_2_XNOR2X1_98 ( );
FILL FILL_3_XNOR2X1_98 ( );
FILL FILL_0_DFFPOSX1_317 ( );
FILL FILL_1_DFFPOSX1_317 ( );
FILL FILL_2_DFFPOSX1_317 ( );
FILL FILL_3_DFFPOSX1_317 ( );
FILL FILL_4_DFFPOSX1_317 ( );
FILL FILL_5_DFFPOSX1_317 ( );
FILL FILL_6_DFFPOSX1_317 ( );
FILL FILL_0_OAI21X1_1467 ( );
FILL FILL_1_OAI21X1_1467 ( );
FILL FILL_0_OAI21X1_1468 ( );
FILL FILL_1_OAI21X1_1468 ( );
FILL FILL_0_INVX2_98 ( );
FILL FILL_0_NAND2X1_527 ( );
FILL FILL_1_NAND2X1_527 ( );
FILL FILL_0_OAI21X1_1471 ( );
FILL FILL_1_OAI21X1_1471 ( );
FILL FILL_0_OAI21X1_1462 ( );
FILL FILL_1_OAI21X1_1462 ( );
FILL FILL_0_DFFPOSX1_963 ( );
FILL FILL_1_DFFPOSX1_963 ( );
FILL FILL_2_DFFPOSX1_963 ( );
FILL FILL_3_DFFPOSX1_963 ( );
FILL FILL_4_DFFPOSX1_963 ( );
FILL FILL_5_DFFPOSX1_963 ( );
FILL FILL_0_NAND2X1_634 ( );
FILL FILL_1_NAND2X1_634 ( );
FILL FILL_0_DFFPOSX1_787 ( );
FILL FILL_1_DFFPOSX1_787 ( );
FILL FILL_2_DFFPOSX1_787 ( );
FILL FILL_3_DFFPOSX1_787 ( );
FILL FILL_4_DFFPOSX1_787 ( );
FILL FILL_5_DFFPOSX1_787 ( );
FILL FILL_6_DFFPOSX1_787 ( );
FILL FILL_0_OAI21X1_1079 ( );
FILL FILL_1_OAI21X1_1079 ( );
FILL FILL_0_NAND2X1_445 ( );
FILL FILL_0_INVX2_99 ( );
FILL FILL_0_NOR2X1_233 ( );
FILL FILL_1_NOR2X1_233 ( );
FILL FILL_0_OAI21X1_1481 ( );
FILL FILL_1_OAI21X1_1481 ( );
FILL FILL_2_OAI21X1_1481 ( );
FILL FILL_0_AOI21X1_49 ( );
FILL FILL_1_AOI21X1_49 ( );
FILL FILL_0_OAI21X1_1296 ( );
FILL FILL_1_OAI21X1_1296 ( );
FILL FILL_0_NAND2X1_552 ( );
FILL FILL_0_INVX4_39 ( );
FILL FILL_1_INVX4_39 ( );
FILL FILL_0_DFFPOSX1_904 ( );
FILL FILL_1_DFFPOSX1_904 ( );
FILL FILL_2_DFFPOSX1_904 ( );
FILL FILL_3_DFFPOSX1_904 ( );
FILL FILL_4_DFFPOSX1_904 ( );
FILL FILL_5_DFFPOSX1_904 ( );
FILL FILL_6_DFFPOSX1_904 ( );
FILL FILL_0_OAI21X1_1173 ( );
FILL FILL_1_OAI21X1_1173 ( );
FILL FILL_0_DFFPOSX1_853 ( );
FILL FILL_1_DFFPOSX1_853 ( );
FILL FILL_2_DFFPOSX1_853 ( );
FILL FILL_3_DFFPOSX1_853 ( );
FILL FILL_4_DFFPOSX1_853 ( );
FILL FILL_5_DFFPOSX1_853 ( );
FILL FILL_0_OAI21X1_1081 ( );
FILL FILL_1_OAI21X1_1081 ( );
FILL FILL_0_DFFPOSX1_789 ( );
FILL FILL_1_DFFPOSX1_789 ( );
FILL FILL_2_DFFPOSX1_789 ( );
FILL FILL_3_DFFPOSX1_789 ( );
FILL FILL_4_DFFPOSX1_789 ( );
FILL FILL_5_DFFPOSX1_789 ( );
FILL FILL_6_DFFPOSX1_789 ( );
FILL FILL_0_NAND2X1_561 ( );
FILL FILL_1_NAND2X1_561 ( );
FILL FILL_0_AOI21X1_40 ( );
FILL FILL_1_AOI21X1_40 ( );
FILL FILL_0_INVX2_82 ( );
FILL FILL_0_NOR2X1_164 ( );
FILL FILL_0_OAI21X1_1340 ( );
FILL FILL_1_OAI21X1_1340 ( );
FILL FILL_0_OAI21X1_1337 ( );
FILL FILL_1_OAI21X1_1337 ( );
FILL FILL_0_OAI21X1_1520 ( );
FILL FILL_1_OAI21X1_1520 ( );
FILL FILL_0_INVX1_212 ( );
FILL FILL_0_AOI21X1_53 ( );
FILL FILL_1_AOI21X1_53 ( );
FILL FILL_0_NOR2X1_205 ( );
FILL FILL_0_CLKBUF1_30 ( );
FILL FILL_1_CLKBUF1_30 ( );
FILL FILL_2_CLKBUF1_30 ( );
FILL FILL_3_CLKBUF1_30 ( );
FILL FILL_0_OAI21X1_1571 ( );
FILL FILL_1_OAI21X1_1571 ( );
FILL FILL_0_DFFPOSX1_998 ( );
FILL FILL_1_DFFPOSX1_998 ( );
FILL FILL_2_DFFPOSX1_998 ( );
FILL FILL_3_DFFPOSX1_998 ( );
FILL FILL_4_DFFPOSX1_998 ( );
FILL FILL_5_DFFPOSX1_998 ( );
FILL FILL_0_DFFPOSX1_806 ( );
FILL FILL_1_DFFPOSX1_806 ( );
FILL FILL_2_DFFPOSX1_806 ( );
FILL FILL_3_DFFPOSX1_806 ( );
FILL FILL_4_DFFPOSX1_806 ( );
FILL FILL_5_DFFPOSX1_806 ( );
FILL FILL_6_DFFPOSX1_806 ( );
FILL FILL_0_OAI21X1_278 ( );
FILL FILL_1_OAI21X1_278 ( );
FILL FILL_0_DFFPOSX1_615 ( );
FILL FILL_1_DFFPOSX1_615 ( );
FILL FILL_2_DFFPOSX1_615 ( );
FILL FILL_3_DFFPOSX1_615 ( );
FILL FILL_4_DFFPOSX1_615 ( );
FILL FILL_5_DFFPOSX1_615 ( );
FILL FILL_0_INVX1_179 ( );
FILL FILL_0_OAI21X1_1084 ( );
FILL FILL_1_OAI21X1_1084 ( );
FILL FILL_0_NAND2X1_450 ( );
FILL FILL_1_NAND2X1_450 ( );
FILL FILL_0_DFFPOSX1_792 ( );
FILL FILL_1_DFFPOSX1_792 ( );
FILL FILL_2_DFFPOSX1_792 ( );
FILL FILL_3_DFFPOSX1_792 ( );
FILL FILL_4_DFFPOSX1_792 ( );
FILL FILL_5_DFFPOSX1_792 ( );
FILL FILL_0_NAND2X1_14 ( );
FILL FILL_1_NAND2X1_14 ( );
FILL FILL_0_OAI21X1_1813 ( );
FILL FILL_1_OAI21X1_1813 ( );
FILL FILL_0_DFFPOSX1_139 ( );
FILL FILL_1_DFFPOSX1_139 ( );
FILL FILL_2_DFFPOSX1_139 ( );
FILL FILL_3_DFFPOSX1_139 ( );
FILL FILL_4_DFFPOSX1_139 ( );
FILL FILL_5_DFFPOSX1_139 ( );
FILL FILL_6_DFFPOSX1_139 ( );
FILL FILL_0_BUFX2_252 ( );
FILL FILL_1_BUFX2_252 ( );
FILL FILL_0_BUFX2_1030 ( );
FILL FILL_1_BUFX2_1030 ( );
FILL FILL_0_BUFX2_888 ( );
FILL FILL_0_INVX2_153 ( );
FILL FILL_0_BUFX2_266 ( );
FILL FILL_1_BUFX2_266 ( );
FILL FILL_0_OAI21X1_849 ( );
FILL FILL_1_OAI21X1_849 ( );
FILL FILL_0_INVX1_50 ( );
FILL FILL_0_DFFPOSX1_621 ( );
FILL FILL_1_DFFPOSX1_621 ( );
FILL FILL_2_DFFPOSX1_621 ( );
FILL FILL_3_DFFPOSX1_621 ( );
FILL FILL_4_DFFPOSX1_621 ( );
FILL FILL_5_DFFPOSX1_621 ( );
FILL FILL_0_BUFX2_66 ( );
FILL FILL_0_OAI21X1_39 ( );
FILL FILL_1_OAI21X1_39 ( );
FILL FILL_0_DFFPOSX1_195 ( );
FILL FILL_1_DFFPOSX1_195 ( );
FILL FILL_2_DFFPOSX1_195 ( );
FILL FILL_3_DFFPOSX1_195 ( );
FILL FILL_4_DFFPOSX1_195 ( );
FILL FILL_5_DFFPOSX1_195 ( );
FILL FILL_6_DFFPOSX1_195 ( );
FILL FILL_0_BUFX2_899 ( );
FILL FILL_1_BUFX2_899 ( );
FILL FILL_0_NAND2X1_69 ( );
FILL FILL_1_NAND2X1_69 ( );
FILL FILL_0_OAI21X1_69 ( );
FILL FILL_1_OAI21X1_69 ( );
FILL FILL_0_DFFPOSX1_225 ( );
FILL FILL_1_DFFPOSX1_225 ( );
FILL FILL_2_DFFPOSX1_225 ( );
FILL FILL_3_DFFPOSX1_225 ( );
FILL FILL_4_DFFPOSX1_225 ( );
FILL FILL_5_DFFPOSX1_225 ( );
FILL FILL_0_CLKBUF1_61 ( );
FILL FILL_1_CLKBUF1_61 ( );
FILL FILL_2_CLKBUF1_61 ( );
FILL FILL_3_CLKBUF1_61 ( );
FILL FILL_4_CLKBUF1_61 ( );
FILL FILL_0_BUFX2_983 ( );
FILL FILL_1_BUFX2_983 ( );
FILL FILL_0_DFFPOSX1_79 ( );
FILL FILL_1_DFFPOSX1_79 ( );
FILL FILL_2_DFFPOSX1_79 ( );
FILL FILL_3_DFFPOSX1_79 ( );
FILL FILL_4_DFFPOSX1_79 ( );
FILL FILL_5_DFFPOSX1_79 ( );
FILL FILL_0_CLKBUF1_64 ( );
FILL FILL_1_CLKBUF1_64 ( );
FILL FILL_2_CLKBUF1_64 ( );
FILL FILL_3_CLKBUF1_64 ( );
FILL FILL_4_CLKBUF1_64 ( );
FILL FILL_0_BUFX2_734 ( );
FILL FILL_1_BUFX2_734 ( );
FILL FILL_0_OAI21X1_323 ( );
FILL FILL_1_OAI21X1_323 ( );
FILL FILL_0_DFFPOSX1_353 ( );
FILL FILL_1_DFFPOSX1_353 ( );
FILL FILL_2_DFFPOSX1_353 ( );
FILL FILL_3_DFFPOSX1_353 ( );
FILL FILL_4_DFFPOSX1_353 ( );
FILL FILL_5_DFFPOSX1_353 ( );
FILL FILL_0_BUFX2_557 ( );
FILL FILL_1_BUFX2_557 ( );
FILL FILL_0_BUFX2_256 ( );
FILL FILL_0_OAI21X1_635 ( );
FILL FILL_1_OAI21X1_635 ( );
FILL FILL_0_DFFPOSX1_537 ( );
FILL FILL_1_DFFPOSX1_537 ( );
FILL FILL_2_DFFPOSX1_537 ( );
FILL FILL_3_DFFPOSX1_537 ( );
FILL FILL_4_DFFPOSX1_537 ( );
FILL FILL_5_DFFPOSX1_537 ( );
FILL FILL_0_BUFX2_439 ( );
FILL FILL_1_BUFX2_439 ( );
FILL FILL_0_DFFPOSX1_406 ( );
FILL FILL_1_DFFPOSX1_406 ( );
FILL FILL_2_DFFPOSX1_406 ( );
FILL FILL_3_DFFPOSX1_406 ( );
FILL FILL_4_DFFPOSX1_406 ( );
FILL FILL_5_DFFPOSX1_406 ( );
FILL FILL_6_DFFPOSX1_406 ( );
FILL FILL_0_NAND2X1_122 ( );
FILL FILL_0_OAI21X1_378 ( );
FILL FILL_1_OAI21X1_378 ( );
FILL FILL_2_OAI21X1_378 ( );
FILL FILL_0_NOR2X1_93 ( );
FILL FILL_0_DFFPOSX1_405 ( );
FILL FILL_1_DFFPOSX1_405 ( );
FILL FILL_2_DFFPOSX1_405 ( );
FILL FILL_3_DFFPOSX1_405 ( );
FILL FILL_4_DFFPOSX1_405 ( );
FILL FILL_5_DFFPOSX1_405 ( );
FILL FILL_0_OAI21X1_525 ( );
FILL FILL_1_OAI21X1_525 ( );
FILL FILL_0_OAI21X1_526 ( );
FILL FILL_1_OAI21X1_526 ( );
FILL FILL_0_INVX2_33 ( );
FILL FILL_0_BUFX2_628 ( );
FILL FILL_0_OAI21X1_798 ( );
FILL FILL_1_OAI21X1_798 ( );
FILL FILL_0_OAI21X1_799 ( );
FILL FILL_1_OAI21X1_799 ( );
FILL FILL_0_DFFPOSX1_596 ( );
FILL FILL_1_DFFPOSX1_596 ( );
FILL FILL_2_DFFPOSX1_596 ( );
FILL FILL_3_DFFPOSX1_596 ( );
FILL FILL_4_DFFPOSX1_596 ( );
FILL FILL_5_DFFPOSX1_596 ( );
FILL FILL_6_DFFPOSX1_596 ( );
FILL FILL_0_DFFPOSX1_595 ( );
FILL FILL_1_DFFPOSX1_595 ( );
FILL FILL_2_DFFPOSX1_595 ( );
FILL FILL_3_DFFPOSX1_595 ( );
FILL FILL_4_DFFPOSX1_595 ( );
FILL FILL_5_DFFPOSX1_595 ( );
FILL FILL_0_OAI21X1_796 ( );
FILL FILL_1_OAI21X1_796 ( );
FILL FILL_0_OAI21X1_813 ( );
FILL FILL_1_OAI21X1_813 ( );
FILL FILL_0_OAI21X1_812 ( );
FILL FILL_1_OAI21X1_812 ( );
FILL FILL_0_BUFX4_161 ( );
FILL FILL_1_BUFX4_161 ( );
FILL FILL_0_CLKBUF1_5 ( );
FILL FILL_1_CLKBUF1_5 ( );
FILL FILL_2_CLKBUF1_5 ( );
FILL FILL_3_CLKBUF1_5 ( );
FILL FILL_4_CLKBUF1_5 ( );
FILL FILL_0_BUFX4_156 ( );
FILL FILL_1_BUFX4_156 ( );
FILL FILL_0_OAI21X1_240 ( );
FILL FILL_1_OAI21X1_240 ( );
FILL FILL_2_OAI21X1_240 ( );
FILL FILL_0_OAI21X1_241 ( );
FILL FILL_1_OAI21X1_241 ( );
FILL FILL_0_DFFPOSX1_479 ( );
FILL FILL_1_DFFPOSX1_479 ( );
FILL FILL_2_DFFPOSX1_479 ( );
FILL FILL_3_DFFPOSX1_479 ( );
FILL FILL_4_DFFPOSX1_479 ( );
FILL FILL_5_DFFPOSX1_479 ( );
FILL FILL_6_DFFPOSX1_479 ( );
FILL FILL_0_OAI21X1_492 ( );
FILL FILL_1_OAI21X1_492 ( );
FILL FILL_0_AOI21X1_4 ( );
FILL FILL_1_AOI21X1_4 ( );
FILL FILL_0_NAND2X1_258 ( );
FILL FILL_1_NAND2X1_258 ( );
FILL FILL_0_OAI21X1_838 ( );
FILL FILL_1_OAI21X1_838 ( );
FILL FILL_0_DFFPOSX1_609 ( );
FILL FILL_1_DFFPOSX1_609 ( );
FILL FILL_2_DFFPOSX1_609 ( );
FILL FILL_3_DFFPOSX1_609 ( );
FILL FILL_4_DFFPOSX1_609 ( );
FILL FILL_5_DFFPOSX1_609 ( );
FILL FILL_6_DFFPOSX1_609 ( );
FILL FILL_0_OAI21X1_837 ( );
FILL FILL_1_OAI21X1_837 ( );
FILL FILL_0_OAI21X1_836 ( );
FILL FILL_1_OAI21X1_836 ( );
FILL FILL_0_NOR2X1_119 ( );
FILL FILL_1_NOR2X1_119 ( );
FILL FILL_0_AOI21X1_35 ( );
FILL FILL_1_AOI21X1_35 ( );
FILL FILL_2_AOI21X1_35 ( );
FILL FILL_0_BUFX2_515 ( );
FILL FILL_1_BUFX2_515 ( );
FILL FILL_0_OAI21X1_388 ( );
FILL FILL_1_OAI21X1_388 ( );
FILL FILL_2_OAI21X1_388 ( );
FILL FILL_0_BUFX2_614 ( );
FILL FILL_1_BUFX2_614 ( );
FILL FILL_0_DFFPOSX1_482 ( );
FILL FILL_1_DFFPOSX1_482 ( );
FILL FILL_2_DFFPOSX1_482 ( );
FILL FILL_3_DFFPOSX1_482 ( );
FILL FILL_4_DFFPOSX1_482 ( );
FILL FILL_5_DFFPOSX1_482 ( );
FILL FILL_0_NAND2X1_110 ( );
FILL FILL_1_NAND2X1_110 ( );
FILL FILL_0_OAI21X1_366 ( );
FILL FILL_1_OAI21X1_366 ( );
FILL FILL_0_OAI21X1_346 ( );
FILL FILL_1_OAI21X1_346 ( );
FILL FILL_0_DFFPOSX1_392 ( );
FILL FILL_1_DFFPOSX1_392 ( );
FILL FILL_2_DFFPOSX1_392 ( );
FILL FILL_3_DFFPOSX1_392 ( );
FILL FILL_4_DFFPOSX1_392 ( );
FILL FILL_5_DFFPOSX1_392 ( );
FILL FILL_0_OAI21X1_714 ( );
FILL FILL_1_OAI21X1_714 ( );
FILL FILL_2_OAI21X1_714 ( );
FILL FILL_0_BUFX4_281 ( );
FILL FILL_1_BUFX4_281 ( );
FILL FILL_0_BUFX4_64 ( );
FILL FILL_1_BUFX4_64 ( );
FILL FILL_0_NAND2X1_17 ( );
FILL FILL_1_NAND2X1_17 ( );
FILL FILL_0_BUFX2_487 ( );
FILL FILL_1_BUFX2_487 ( );
FILL FILL_0_DFFPOSX1_951 ( );
FILL FILL_1_DFFPOSX1_951 ( );
FILL FILL_2_DFFPOSX1_951 ( );
FILL FILL_3_DFFPOSX1_951 ( );
FILL FILL_4_DFFPOSX1_951 ( );
FILL FILL_5_DFFPOSX1_951 ( );
FILL FILL_0_OAI21X1_765 ( );
FILL FILL_1_OAI21X1_765 ( );
FILL FILL_0_OAI21X1_764 ( );
FILL FILL_1_OAI21X1_764 ( );
FILL FILL_0_OAI21X1_744 ( );
FILL FILL_1_OAI21X1_744 ( );
FILL FILL_0_CLKBUF1_23 ( );
FILL FILL_1_CLKBUF1_23 ( );
FILL FILL_2_CLKBUF1_23 ( );
FILL FILL_3_CLKBUF1_23 ( );
FILL FILL_0_BUFX4_127 ( );
FILL FILL_1_BUFX4_127 ( );
FILL FILL_0_OAI21X1_1245 ( );
FILL FILL_1_OAI21X1_1245 ( );
FILL FILL_0_DFFPOSX1_885 ( );
FILL FILL_1_DFFPOSX1_885 ( );
FILL FILL_2_DFFPOSX1_885 ( );
FILL FILL_3_DFFPOSX1_885 ( );
FILL FILL_4_DFFPOSX1_885 ( );
FILL FILL_5_DFFPOSX1_885 ( );
FILL FILL_0_OAI21X1_1244 ( );
FILL FILL_1_OAI21X1_1244 ( );
FILL FILL_2_OAI21X1_1244 ( );
FILL FILL_0_OAI21X1_104 ( );
FILL FILL_1_OAI21X1_104 ( );
FILL FILL_0_DFFPOSX1_510 ( );
FILL FILL_1_DFFPOSX1_510 ( );
FILL FILL_2_DFFPOSX1_510 ( );
FILL FILL_3_DFFPOSX1_510 ( );
FILL FILL_4_DFFPOSX1_510 ( );
FILL FILL_5_DFFPOSX1_510 ( );
FILL FILL_6_DFFPOSX1_510 ( );
FILL FILL_0_AND2X2_26 ( );
FILL FILL_1_AND2X2_26 ( );
FILL FILL_2_AND2X2_26 ( );
FILL FILL_0_NAND2X1_598 ( );
FILL FILL_1_NAND2X1_598 ( );
FILL FILL_0_DFFPOSX1_349 ( );
FILL FILL_1_DFFPOSX1_349 ( );
FILL FILL_2_DFFPOSX1_349 ( );
FILL FILL_3_DFFPOSX1_349 ( );
FILL FILL_4_DFFPOSX1_349 ( );
FILL FILL_5_DFFPOSX1_349 ( );
FILL FILL_6_DFFPOSX1_349 ( );
FILL FILL_0_BUFX4_291 ( );
FILL FILL_1_BUFX4_291 ( );
FILL FILL_2_BUFX4_291 ( );
FILL FILL_0_BUFX2_699 ( );
FILL FILL_1_BUFX2_699 ( );
FILL FILL_0_OAI21X1_195 ( );
FILL FILL_1_OAI21X1_195 ( );
FILL FILL_0_BUFX2_11 ( );
FILL FILL_1_BUFX2_11 ( );
FILL FILL_0_OAI21X1_1282 ( );
FILL FILL_1_OAI21X1_1282 ( );
FILL FILL_2_OAI21X1_1282 ( );
FILL FILL_0_OAI21X1_1281 ( );
FILL FILL_1_OAI21X1_1281 ( );
FILL FILL_0_OAI21X1_1457 ( );
FILL FILL_1_OAI21X1_1457 ( );
FILL FILL_0_DFFPOSX1_961 ( );
FILL FILL_1_DFFPOSX1_961 ( );
FILL FILL_2_DFFPOSX1_961 ( );
FILL FILL_3_DFFPOSX1_961 ( );
FILL FILL_4_DFFPOSX1_961 ( );
FILL FILL_5_DFFPOSX1_961 ( );
FILL FILL_0_CLKBUF1_3 ( );
FILL FILL_1_CLKBUF1_3 ( );
FILL FILL_2_CLKBUF1_3 ( );
FILL FILL_3_CLKBUF1_3 ( );
FILL FILL_4_CLKBUF1_3 ( );
FILL FILL_0_OAI21X1_1285 ( );
FILL FILL_1_OAI21X1_1285 ( );
FILL FILL_0_DFFPOSX1_772 ( );
FILL FILL_1_DFFPOSX1_772 ( );
FILL FILL_2_DFFPOSX1_772 ( );
FILL FILL_3_DFFPOSX1_772 ( );
FILL FILL_4_DFFPOSX1_772 ( );
FILL FILL_5_DFFPOSX1_772 ( );
FILL FILL_6_DFFPOSX1_772 ( );
FILL FILL_0_OAI21X1_1064 ( );
FILL FILL_1_OAI21X1_1064 ( );
FILL FILL_0_OAI21X1_1463 ( );
FILL FILL_1_OAI21X1_1463 ( );
FILL FILL_0_INVX1_176 ( );
FILL FILL_0_OAI21X1_1063 ( );
FILL FILL_1_OAI21X1_1063 ( );
FILL FILL_0_NAND2X1_429 ( );
FILL FILL_1_NAND2X1_429 ( );
FILL FILL_0_OAI21X1_1464 ( );
FILL FILL_1_OAI21X1_1464 ( );
FILL FILL_0_OAI21X1_250 ( );
FILL FILL_1_OAI21X1_250 ( );
FILL FILL_0_OAI21X1_251 ( );
FILL FILL_1_OAI21X1_251 ( );
FILL FILL_0_NOR2X1_145 ( );
FILL FILL_0_XNOR2X1_66 ( );
FILL FILL_1_XNOR2X1_66 ( );
FILL FILL_2_XNOR2X1_66 ( );
FILL FILL_3_XNOR2X1_66 ( );
FILL FILL_0_OAI21X1_75 ( );
FILL FILL_1_OAI21X1_75 ( );
FILL FILL_0_DFFPOSX1_902 ( );
FILL FILL_1_DFFPOSX1_902 ( );
FILL FILL_2_DFFPOSX1_902 ( );
FILL FILL_3_DFFPOSX1_902 ( );
FILL FILL_4_DFFPOSX1_902 ( );
FILL FILL_5_DFFPOSX1_902 ( );
FILL FILL_6_DFFPOSX1_902 ( );
FILL FILL_0_BUFX4_292 ( );
FILL FILL_1_BUFX4_292 ( );
FILL FILL_0_OAI21X1_1473 ( );
FILL FILL_1_OAI21X1_1473 ( );
FILL FILL_0_NOR2X1_150 ( );
FILL FILL_1_NOR2X1_150 ( );
FILL FILL_0_DFFPOSX1_966 ( );
FILL FILL_1_DFFPOSX1_966 ( );
FILL FILL_2_DFFPOSX1_966 ( );
FILL FILL_3_DFFPOSX1_966 ( );
FILL FILL_4_DFFPOSX1_966 ( );
FILL FILL_5_DFFPOSX1_966 ( );
FILL FILL_0_CLKBUF1_27 ( );
FILL FILL_1_CLKBUF1_27 ( );
FILL FILL_2_CLKBUF1_27 ( );
FILL FILL_3_CLKBUF1_27 ( );
FILL FILL_4_CLKBUF1_27 ( );
FILL FILL_0_NAND3X1_41 ( );
FILL FILL_1_NAND3X1_41 ( );
FILL FILL_0_BUFX4_23 ( );
FILL FILL_1_BUFX4_23 ( );
FILL FILL_0_OAI21X1_1477 ( );
FILL FILL_1_OAI21X1_1477 ( );
FILL FILL_0_OAI21X1_1476 ( );
FILL FILL_1_OAI21X1_1476 ( );
FILL FILL_0_INVX2_75 ( );
FILL FILL_0_BUFX2_156 ( );
FILL FILL_1_BUFX2_156 ( );
FILL FILL_0_NAND2X1_555 ( );
FILL FILL_0_OAI21X1_1069 ( );
FILL FILL_1_OAI21X1_1069 ( );
FILL FILL_0_NAND2X1_435 ( );
FILL FILL_1_NAND2X1_435 ( );
FILL FILL_0_DFFPOSX1_777 ( );
FILL FILL_1_DFFPOSX1_777 ( );
FILL FILL_2_DFFPOSX1_777 ( );
FILL FILL_3_DFFPOSX1_777 ( );
FILL FILL_4_DFFPOSX1_777 ( );
FILL FILL_5_DFFPOSX1_777 ( );
FILL FILL_0_OAI21X1_1303 ( );
FILL FILL_1_OAI21X1_1303 ( );
FILL FILL_0_OAI21X1_1178 ( );
FILL FILL_1_OAI21X1_1178 ( );
FILL FILL_0_OAI21X1_1177 ( );
FILL FILL_1_OAI21X1_1177 ( );
FILL FILL_0_OAI21X1_1295 ( );
FILL FILL_1_OAI21X1_1295 ( );
FILL FILL_0_NAND2X1_447 ( );
FILL FILL_1_NAND2X1_447 ( );
FILL FILL_0_BUFX4_381 ( );
FILL FILL_1_BUFX4_381 ( );
FILL FILL_0_OAI21X1_1176 ( );
FILL FILL_1_OAI21X1_1176 ( );
FILL FILL_0_OAI21X1_1175 ( );
FILL FILL_1_OAI21X1_1175 ( );
FILL FILL_0_OAI21X1_1341 ( );
FILL FILL_1_OAI21X1_1341 ( );
FILL FILL_0_OAI21X1_1339 ( );
FILL FILL_1_OAI21X1_1339 ( );
FILL FILL_0_DFFPOSX1_906 ( );
FILL FILL_1_DFFPOSX1_906 ( );
FILL FILL_2_DFFPOSX1_906 ( );
FILL FILL_3_DFFPOSX1_906 ( );
FILL FILL_4_DFFPOSX1_906 ( );
FILL FILL_5_DFFPOSX1_906 ( );
FILL FILL_6_DFFPOSX1_906 ( );
FILL FILL_0_OAI21X1_1338 ( );
FILL FILL_1_OAI21X1_1338 ( );
FILL FILL_2_OAI21X1_1338 ( );
FILL FILL_0_OAI21X1_1336 ( );
FILL FILL_1_OAI21X1_1336 ( );
FILL FILL_0_BUFX2_234 ( );
FILL FILL_1_BUFX2_234 ( );
FILL FILL_0_BUFX2_41 ( );
FILL FILL_1_BUFX2_41 ( );
FILL FILL_0_NAND2X1_464 ( );
FILL FILL_0_OAI21X1_1083 ( );
FILL FILL_1_OAI21X1_1083 ( );
FILL FILL_0_DFFPOSX1_791 ( );
FILL FILL_1_DFFPOSX1_791 ( );
FILL FILL_2_DFFPOSX1_791 ( );
FILL FILL_3_DFFPOSX1_791 ( );
FILL FILL_4_DFFPOSX1_791 ( );
FILL FILL_5_DFFPOSX1_791 ( );
FILL FILL_6_DFFPOSX1_791 ( );
FILL FILL_0_NAND2X1_449 ( );
FILL FILL_1_NAND2X1_449 ( );
FILL FILL_0_BUFX2_235 ( );
FILL FILL_0_BUFX2_60 ( );
FILL FILL_1_BUFX2_60 ( );
FILL FILL_0_DFFPOSX1_24 ( );
FILL FILL_1_DFFPOSX1_24 ( );
FILL FILL_2_DFFPOSX1_24 ( );
FILL FILL_3_DFFPOSX1_24 ( );
FILL FILL_4_DFFPOSX1_24 ( );
FILL FILL_5_DFFPOSX1_24 ( );
FILL FILL_6_DFFPOSX1_24 ( );
FILL FILL_0_OAI21X1_1634 ( );
FILL FILL_1_OAI21X1_1634 ( );
FILL FILL_0_NAND2X1_702 ( );
FILL FILL_1_NAND2X1_702 ( );
FILL FILL_0_NAND2X1_754 ( );
FILL FILL_1_NAND2X1_754 ( );
FILL FILL_0_BUFX4_219 ( );
FILL FILL_1_BUFX4_219 ( );
FILL FILL_0_BUFX2_44 ( );
FILL FILL_1_BUFX2_44 ( );
FILL FILL_0_BUFX2_1002 ( );
FILL FILL_0_BUFX2_42 ( );
FILL FILL_1_BUFX2_42 ( );
FILL FILL_0_BUFX2_694 ( );
FILL FILL_1_BUFX2_694 ( );
FILL FILL_0_BUFX2_897 ( );
FILL FILL_1_BUFX2_897 ( );
FILL FILL_0_BUFX2_260 ( );
FILL FILL_1_BUFX2_260 ( );
FILL FILL_0_BUFX2_288 ( );
FILL FILL_1_BUFX2_288 ( );
FILL FILL_0_INVX1_158 ( );
FILL FILL_0_INVX1_79 ( );
FILL FILL_0_BUFX2_802 ( );
FILL FILL_0_OAI21X1_878 ( );
FILL FILL_1_OAI21X1_878 ( );
FILL FILL_0_DFFPOSX1_650 ( );
FILL FILL_1_DFFPOSX1_650 ( );
FILL FILL_2_DFFPOSX1_650 ( );
FILL FILL_3_DFFPOSX1_650 ( );
FILL FILL_4_DFFPOSX1_650 ( );
FILL FILL_5_DFFPOSX1_650 ( );
FILL FILL_6_DFFPOSX1_650 ( );
FILL FILL_0_BUFX2_366 ( );
FILL FILL_1_BUFX2_366 ( );
FILL FILL_0_NAND2X1_746 ( );
FILL FILL_0_OAI21X1_1805 ( );
FILL FILL_1_OAI21X1_1805 ( );
FILL FILL_0_DFFPOSX1_131 ( );
FILL FILL_1_DFFPOSX1_131 ( );
FILL FILL_2_DFFPOSX1_131 ( );
FILL FILL_3_DFFPOSX1_131 ( );
FILL FILL_4_DFFPOSX1_131 ( );
FILL FILL_5_DFFPOSX1_131 ( );
FILL FILL_0_BUFX4_366 ( );
FILL FILL_1_BUFX4_366 ( );
FILL FILL_0_OAI21X1_1007 ( );
FILL FILL_1_OAI21X1_1007 ( );
FILL FILL_0_OAI21X1_1006 ( );
FILL FILL_1_OAI21X1_1006 ( );
FILL FILL_2_OAI21X1_1006 ( );
FILL FILL_0_OAI21X1_1732 ( );
FILL FILL_1_OAI21X1_1732 ( );
FILL FILL_0_OAI21X1_1733 ( );
FILL FILL_1_OAI21X1_1733 ( );
FILL FILL_0_NAND2X1_29 ( );
FILL FILL_0_OAI21X1_29 ( );
FILL FILL_1_OAI21X1_29 ( );
FILL FILL_0_BUFX4_151 ( );
FILL FILL_1_BUFX4_151 ( );
FILL FILL_0_DFFPOSX1_96 ( );
FILL FILL_1_DFFPOSX1_96 ( );
FILL FILL_2_DFFPOSX1_96 ( );
FILL FILL_3_DFFPOSX1_96 ( );
FILL FILL_4_DFFPOSX1_96 ( );
FILL FILL_5_DFFPOSX1_96 ( );
FILL FILL_6_DFFPOSX1_96 ( );
FILL FILL_0_OAI21X1_322 ( );
FILL FILL_1_OAI21X1_322 ( );
FILL FILL_0_DFFPOSX1_938 ( );
FILL FILL_1_DFFPOSX1_938 ( );
FILL FILL_2_DFFPOSX1_938 ( );
FILL FILL_3_DFFPOSX1_938 ( );
FILL FILL_4_DFFPOSX1_938 ( );
FILL FILL_5_DFFPOSX1_938 ( );
FILL FILL_0_BUFX4_296 ( );
FILL FILL_1_BUFX4_296 ( );
FILL FILL_0_BUFX2_568 ( );
FILL FILL_0_DFFPOSX1_471 ( );
FILL FILL_1_DFFPOSX1_471 ( );
FILL FILL_2_DFFPOSX1_471 ( );
FILL FILL_3_DFFPOSX1_471 ( );
FILL FILL_4_DFFPOSX1_471 ( );
FILL FILL_5_DFFPOSX1_471 ( );
FILL FILL_6_DFFPOSX1_471 ( );
FILL FILL_0_OAI21X1_478 ( );
FILL FILL_1_OAI21X1_478 ( );
FILL FILL_0_BUFX2_437 ( );
FILL FILL_1_BUFX2_437 ( );
FILL FILL_0_DFFPOSX1_407 ( );
FILL FILL_1_DFFPOSX1_407 ( );
FILL FILL_2_DFFPOSX1_407 ( );
FILL FILL_3_DFFPOSX1_407 ( );
FILL FILL_4_DFFPOSX1_407 ( );
FILL FILL_5_DFFPOSX1_407 ( );
FILL FILL_0_NAND2X1_123 ( );
FILL FILL_0_OAI21X1_379 ( );
FILL FILL_1_OAI21X1_379 ( );
FILL FILL_0_XNOR2X1_21 ( );
FILL FILL_1_XNOR2X1_21 ( );
FILL FILL_2_XNOR2X1_21 ( );
FILL FILL_3_XNOR2X1_21 ( );
FILL FILL_0_BUFX2_503 ( );
FILL FILL_0_BUFX4_200 ( );
FILL FILL_1_BUFX4_200 ( );
FILL FILL_0_BUFX4_115 ( );
FILL FILL_1_BUFX4_115 ( );
FILL FILL_0_BUFX2_627 ( );
FILL FILL_1_BUFX2_627 ( );
FILL FILL_0_NAND2X1_241 ( );
FILL FILL_0_DFFPOSX1_591 ( );
FILL FILL_1_DFFPOSX1_591 ( );
FILL FILL_2_DFFPOSX1_591 ( );
FILL FILL_3_DFFPOSX1_591 ( );
FILL FILL_4_DFFPOSX1_591 ( );
FILL FILL_5_DFFPOSX1_591 ( );
FILL FILL_0_OAI21X1_781 ( );
FILL FILL_1_OAI21X1_781 ( );
FILL FILL_0_OAI21X1_782 ( );
FILL FILL_1_OAI21X1_782 ( );
FILL FILL_0_DFFPOSX1_600 ( );
FILL FILL_1_DFFPOSX1_600 ( );
FILL FILL_2_DFFPOSX1_600 ( );
FILL FILL_3_DFFPOSX1_600 ( );
FILL FILL_4_DFFPOSX1_600 ( );
FILL FILL_5_DFFPOSX1_600 ( );
FILL FILL_0_OAI21X1_795 ( );
FILL FILL_1_OAI21X1_795 ( );
FILL FILL_0_DFFPOSX1_886 ( );
FILL FILL_1_DFFPOSX1_886 ( );
FILL FILL_2_DFFPOSX1_886 ( );
FILL FILL_3_DFFPOSX1_886 ( );
FILL FILL_4_DFFPOSX1_886 ( );
FILL FILL_5_DFFPOSX1_886 ( );
FILL FILL_0_OAI21X1_829 ( );
FILL FILL_1_OAI21X1_829 ( );
FILL FILL_2_OAI21X1_829 ( );
FILL FILL_0_DFFPOSX1_606 ( );
FILL FILL_1_DFFPOSX1_606 ( );
FILL FILL_2_DFFPOSX1_606 ( );
FILL FILL_3_DFFPOSX1_606 ( );
FILL FILL_4_DFFPOSX1_606 ( );
FILL FILL_5_DFFPOSX1_606 ( );
FILL FILL_0_OAI21X1_830 ( );
FILL FILL_1_OAI21X1_830 ( );
FILL FILL_0_DFFPOSX1_312 ( );
FILL FILL_1_DFFPOSX1_312 ( );
FILL FILL_2_DFFPOSX1_312 ( );
FILL FILL_3_DFFPOSX1_312 ( );
FILL FILL_4_DFFPOSX1_312 ( );
FILL FILL_5_DFFPOSX1_312 ( );
FILL FILL_6_DFFPOSX1_312 ( );
FILL FILL_0_DFFPOSX1_301 ( );
FILL FILL_1_DFFPOSX1_301 ( );
FILL FILL_2_DFFPOSX1_301 ( );
FILL FILL_3_DFFPOSX1_301 ( );
FILL FILL_4_DFFPOSX1_301 ( );
FILL FILL_5_DFFPOSX1_301 ( );
FILL FILL_0_OAI21X1_219 ( );
FILL FILL_1_OAI21X1_219 ( );
FILL FILL_0_OAI21X1_218 ( );
FILL FILL_1_OAI21X1_218 ( );
FILL FILL_0_AOI21X1_27 ( );
FILL FILL_1_AOI21X1_27 ( );
FILL FILL_2_AOI21X1_27 ( );
FILL FILL_0_AOI21X1_28 ( );
FILL FILL_1_AOI21X1_28 ( );
FILL FILL_0_NOR2X1_101 ( );
FILL FILL_0_OR2X2_14 ( );
FILL FILL_1_OR2X2_14 ( );
FILL FILL_0_NOR2X1_57 ( );
FILL FILL_1_NOR2X1_57 ( );
FILL FILL_0_NAND3X1_26 ( );
FILL FILL_1_NAND3X1_26 ( );
FILL FILL_0_INVX4_28 ( );
FILL FILL_1_INVX4_28 ( );
FILL FILL_0_DFFPOSX1_416 ( );
FILL FILL_1_DFFPOSX1_416 ( );
FILL FILL_2_DFFPOSX1_416 ( );
FILL FILL_3_DFFPOSX1_416 ( );
FILL FILL_4_DFFPOSX1_416 ( );
FILL FILL_5_DFFPOSX1_416 ( );
FILL FILL_6_DFFPOSX1_416 ( );
FILL FILL_0_NAND2X1_132 ( );
FILL FILL_0_BUFX4_171 ( );
FILL FILL_1_BUFX4_171 ( );
FILL FILL_0_BUFX2_423 ( );
FILL FILL_0_DFFPOSX1_394 ( );
FILL FILL_1_DFFPOSX1_394 ( );
FILL FILL_2_DFFPOSX1_394 ( );
FILL FILL_3_DFFPOSX1_394 ( );
FILL FILL_4_DFFPOSX1_394 ( );
FILL FILL_5_DFFPOSX1_394 ( );
FILL FILL_0_DFFPOSX1_374 ( );
FILL FILL_1_DFFPOSX1_374 ( );
FILL FILL_2_DFFPOSX1_374 ( );
FILL FILL_3_DFFPOSX1_374 ( );
FILL FILL_4_DFFPOSX1_374 ( );
FILL FILL_5_DFFPOSX1_374 ( );
FILL FILL_0_BUFX2_595 ( );
FILL FILL_1_BUFX2_595 ( );
FILL FILL_0_BUFX2_596 ( );
FILL FILL_1_BUFX2_596 ( );
FILL FILL_0_BUFX2_200 ( );
FILL FILL_1_BUFX2_200 ( );
FILL FILL_0_OAI21X1_1428 ( );
FILL FILL_1_OAI21X1_1428 ( );
FILL FILL_0_OAI21X1_1429 ( );
FILL FILL_1_OAI21X1_1429 ( );
FILL FILL_0_DFFPOSX1_760 ( );
FILL FILL_1_DFFPOSX1_760 ( );
FILL FILL_2_DFFPOSX1_760 ( );
FILL FILL_3_DFFPOSX1_760 ( );
FILL FILL_4_DFFPOSX1_760 ( );
FILL FILL_5_DFFPOSX1_760 ( );
FILL FILL_0_DFFPOSX1_585 ( );
FILL FILL_1_DFFPOSX1_585 ( );
FILL FILL_2_DFFPOSX1_585 ( );
FILL FILL_3_DFFPOSX1_585 ( );
FILL FILL_4_DFFPOSX1_585 ( );
FILL FILL_5_DFFPOSX1_585 ( );
FILL FILL_6_DFFPOSX1_585 ( );
FILL FILL_0_BUFX2_637 ( );
FILL FILL_1_BUFX2_637 ( );
FILL FILL_0_BUFX2_609 ( );
FILL FILL_1_BUFX2_609 ( );
FILL FILL_0_DFFPOSX1_247 ( );
FILL FILL_1_DFFPOSX1_247 ( );
FILL FILL_2_DFFPOSX1_247 ( );
FILL FILL_3_DFFPOSX1_247 ( );
FILL FILL_4_DFFPOSX1_247 ( );
FILL FILL_5_DFFPOSX1_247 ( );
FILL FILL_6_DFFPOSX1_247 ( );
FILL FILL_0_BUFX4_223 ( );
FILL FILL_1_BUFX4_223 ( );
FILL FILL_0_DFFPOSX1_116 ( );
FILL FILL_1_DFFPOSX1_116 ( );
FILL FILL_2_DFFPOSX1_116 ( );
FILL FILL_3_DFFPOSX1_116 ( );
FILL FILL_4_DFFPOSX1_116 ( );
FILL FILL_5_DFFPOSX1_116 ( );
FILL FILL_0_OAI21X1_1790 ( );
FILL FILL_1_OAI21X1_1790 ( );
FILL FILL_0_BUFX2_731 ( );
FILL FILL_1_BUFX2_731 ( );
FILL FILL_0_CLKBUF1_47 ( );
FILL FILL_1_CLKBUF1_47 ( );
FILL FILL_2_CLKBUF1_47 ( );
FILL FILL_3_CLKBUF1_47 ( );
FILL FILL_4_CLKBUF1_47 ( );
FILL FILL_0_BUFX2_913 ( );
FILL FILL_1_BUFX2_913 ( );
FILL FILL_0_OAI21X1_1438 ( );
FILL FILL_1_OAI21X1_1438 ( );
FILL FILL_0_INVX1_201 ( );
FILL FILL_0_BUFX2_1022 ( );
FILL FILL_1_BUFX2_1022 ( );
FILL FILL_0_DFFPOSX1_289 ( );
FILL FILL_1_DFFPOSX1_289 ( );
FILL FILL_2_DFFPOSX1_289 ( );
FILL FILL_3_DFFPOSX1_289 ( );
FILL FILL_4_DFFPOSX1_289 ( );
FILL FILL_5_DFFPOSX1_289 ( );
FILL FILL_6_DFFPOSX1_289 ( );
FILL FILL_0_DFFPOSX1_962 ( );
FILL FILL_1_DFFPOSX1_962 ( );
FILL FILL_2_DFFPOSX1_962 ( );
FILL FILL_3_DFFPOSX1_962 ( );
FILL FILL_4_DFFPOSX1_962 ( );
FILL FILL_5_DFFPOSX1_962 ( );
FILL FILL_6_DFFPOSX1_962 ( );
FILL FILL_0_OAI21X1_194 ( );
FILL FILL_1_OAI21X1_194 ( );
FILL FILL_2_OAI21X1_194 ( );
FILL FILL_0_DFFPOSX1_834 ( );
FILL FILL_1_DFFPOSX1_834 ( );
FILL FILL_2_DFFPOSX1_834 ( );
FILL FILL_3_DFFPOSX1_834 ( );
FILL FILL_4_DFFPOSX1_834 ( );
FILL FILL_5_DFFPOSX1_834 ( );
FILL FILL_0_NOR2X1_143 ( );
FILL FILL_0_INVX1_190 ( );
FILL FILL_1_INVX1_190 ( );
FILL FILL_0_OAI21X1_1456 ( );
FILL FILL_1_OAI21X1_1456 ( );
FILL FILL_0_DFFPOSX1_81 ( );
FILL FILL_1_DFFPOSX1_81 ( );
FILL FILL_2_DFFPOSX1_81 ( );
FILL FILL_3_DFFPOSX1_81 ( );
FILL FILL_4_DFFPOSX1_81 ( );
FILL FILL_5_DFFPOSX1_81 ( );
FILL FILL_6_DFFPOSX1_81 ( );
FILL FILL_0_BUFX4_138 ( );
FILL FILL_1_BUFX4_138 ( );
FILL FILL_0_BUFX4_118 ( );
FILL FILL_1_BUFX4_118 ( );
FILL FILL_2_BUFX4_118 ( );
FILL FILL_0_NAND2X1_430 ( );
FILL FILL_1_NAND2X1_430 ( );
FILL FILL_0_INVX4_38 ( );
FILL FILL_1_INVX4_38 ( );
FILL FILL_0_DFFPOSX1_771 ( );
FILL FILL_1_DFFPOSX1_771 ( );
FILL FILL_2_DFFPOSX1_771 ( );
FILL FILL_3_DFFPOSX1_771 ( );
FILL FILL_4_DFFPOSX1_771 ( );
FILL FILL_5_DFFPOSX1_771 ( );
FILL FILL_0_AOI21X1_48 ( );
FILL FILL_1_AOI21X1_48 ( );
FILL FILL_0_OR2X2_20 ( );
FILL FILL_1_OR2X2_20 ( );
FILL FILL_0_OAI21X1_1292 ( );
FILL FILL_1_OAI21X1_1292 ( );
FILL FILL_2_OAI21X1_1292 ( );
FILL FILL_0_OAI21X1_1291 ( );
FILL FILL_1_OAI21X1_1291 ( );
FILL FILL_0_BUFX4_318 ( );
FILL FILL_1_BUFX4_318 ( );
FILL FILL_0_NAND2X1_529 ( );
FILL FILL_0_DFFPOSX1_229 ( );
FILL FILL_1_DFFPOSX1_229 ( );
FILL FILL_2_DFFPOSX1_229 ( );
FILL FILL_3_DFFPOSX1_229 ( );
FILL FILL_4_DFFPOSX1_229 ( );
FILL FILL_5_DFFPOSX1_229 ( );
FILL FILL_0_NAND2X1_528 ( );
FILL FILL_1_NAND2X1_528 ( );
FILL FILL_0_AOI21X1_37 ( );
FILL FILL_1_AOI21X1_37 ( );
FILL FILL_0_OAI21X1_1151 ( );
FILL FILL_1_OAI21X1_1151 ( );
FILL FILL_0_BUFX2_39 ( );
FILL FILL_1_BUFX2_39 ( );
FILL FILL_0_OAI21X1_1472 ( );
FILL FILL_1_OAI21X1_1472 ( );
FILL FILL_0_XNOR2X1_81 ( );
FILL FILL_1_XNOR2X1_81 ( );
FILL FILL_2_XNOR2X1_81 ( );
FILL FILL_0_OAI21X1_1152 ( );
FILL FILL_1_OAI21X1_1152 ( );
FILL FILL_0_INVX1_191 ( );
FILL FILL_0_DFFPOSX1_839 ( );
FILL FILL_1_DFFPOSX1_839 ( );
FILL FILL_2_DFFPOSX1_839 ( );
FILL FILL_3_DFFPOSX1_839 ( );
FILL FILL_4_DFFPOSX1_839 ( );
FILL FILL_5_DFFPOSX1_839 ( );
FILL FILL_6_DFFPOSX1_839 ( );
FILL FILL_0_CLKBUF1_89 ( );
FILL FILL_1_CLKBUF1_89 ( );
FILL FILL_2_CLKBUF1_89 ( );
FILL FILL_3_CLKBUF1_89 ( );
FILL FILL_4_CLKBUF1_89 ( );
FILL FILL_0_BUFX2_104 ( );
FILL FILL_1_BUFX2_104 ( );
FILL FILL_0_XNOR2X1_99 ( );
FILL FILL_1_XNOR2X1_99 ( );
FILL FILL_2_XNOR2X1_99 ( );
FILL FILL_3_XNOR2X1_99 ( );
FILL FILL_0_OAI21X1_1080 ( );
FILL FILL_1_OAI21X1_1080 ( );
FILL FILL_0_NAND2X1_446 ( );
FILL FILL_0_DFFPOSX1_788 ( );
FILL FILL_1_DFFPOSX1_788 ( );
FILL FILL_2_DFFPOSX1_788 ( );
FILL FILL_3_DFFPOSX1_788 ( );
FILL FILL_4_DFFPOSX1_788 ( );
FILL FILL_5_DFFPOSX1_788 ( );
FILL FILL_0_NAND2X1_560 ( );
FILL FILL_1_NAND2X1_560 ( );
FILL FILL_0_OAI21X1_1302 ( );
FILL FILL_1_OAI21X1_1302 ( );
FILL FILL_0_DFFPOSX1_920 ( );
FILL FILL_1_DFFPOSX1_920 ( );
FILL FILL_2_DFFPOSX1_920 ( );
FILL FILL_3_DFFPOSX1_920 ( );
FILL FILL_4_DFFPOSX1_920 ( );
FILL FILL_5_DFFPOSX1_920 ( );
FILL FILL_0_BUFX4_339 ( );
FILL FILL_1_BUFX4_339 ( );
FILL FILL_0_BUFX2_107 ( );
FILL FILL_1_BUFX2_107 ( );
FILL FILL_0_NAND2X1_559 ( );
FILL FILL_0_DFFPOSX1_716 ( );
FILL FILL_1_DFFPOSX1_716 ( );
FILL FILL_2_DFFPOSX1_716 ( );
FILL FILL_3_DFFPOSX1_716 ( );
FILL FILL_4_DFFPOSX1_716 ( );
FILL FILL_5_DFFPOSX1_716 ( );
FILL FILL_0_BUFX2_233 ( );
FILL FILL_0_BUFX2_172 ( );
FILL FILL_1_BUFX2_172 ( );
FILL FILL_0_DFFPOSX1_613 ( );
FILL FILL_1_DFFPOSX1_613 ( );
FILL FILL_2_DFFPOSX1_613 ( );
FILL FILL_3_DFFPOSX1_613 ( );
FILL FILL_4_DFFPOSX1_613 ( );
FILL FILL_5_DFFPOSX1_613 ( );
FILL FILL_0_DFFPOSX1_919 ( );
FILL FILL_1_DFFPOSX1_919 ( );
FILL FILL_2_DFFPOSX1_919 ( );
FILL FILL_3_DFFPOSX1_919 ( );
FILL FILL_4_DFFPOSX1_919 ( );
FILL FILL_5_DFFPOSX1_919 ( );
FILL FILL_6_DFFPOSX1_919 ( );
FILL FILL_0_CLKBUF1_67 ( );
FILL FILL_1_CLKBUF1_67 ( );
FILL FILL_2_CLKBUF1_67 ( );
FILL FILL_3_CLKBUF1_67 ( );
FILL FILL_4_CLKBUF1_67 ( );
FILL FILL_0_BUFX4_375 ( );
FILL FILL_1_BUFX4_375 ( );
FILL FILL_0_DFFPOSX1_122 ( );
FILL FILL_1_DFFPOSX1_122 ( );
FILL FILL_2_DFFPOSX1_122 ( );
FILL FILL_3_DFFPOSX1_122 ( );
FILL FILL_4_DFFPOSX1_122 ( );
FILL FILL_5_DFFPOSX1_122 ( );
FILL FILL_6_DFFPOSX1_122 ( );
FILL FILL_0_OAI21X1_1796 ( );
FILL FILL_1_OAI21X1_1796 ( );
FILL FILL_0_NAND2X1_737 ( );
FILL FILL_1_NAND2X1_737 ( );
FILL FILL_0_BUFX4_195 ( );
FILL FILL_1_BUFX4_195 ( );
FILL FILL_0_OAI21X1_57 ( );
FILL FILL_1_OAI21X1_57 ( );
FILL FILL_0_NAND2X1_57 ( );
FILL FILL_1_NAND2X1_57 ( );
FILL FILL_0_DFFPOSX1_213 ( );
FILL FILL_1_DFFPOSX1_213 ( );
FILL FILL_2_DFFPOSX1_213 ( );
FILL FILL_3_DFFPOSX1_213 ( );
FILL FILL_4_DFFPOSX1_213 ( );
FILL FILL_5_DFFPOSX1_213 ( );
FILL FILL_6_DFFPOSX1_213 ( );
FILL FILL_0_DFFPOSX1_627 ( );
FILL FILL_1_DFFPOSX1_627 ( );
FILL FILL_2_DFFPOSX1_627 ( );
FILL FILL_3_DFFPOSX1_627 ( );
FILL FILL_4_DFFPOSX1_627 ( );
FILL FILL_5_DFFPOSX1_627 ( );
FILL FILL_6_DFFPOSX1_627 ( );
FILL FILL_0_OAI21X1_855 ( );
FILL FILL_1_OAI21X1_855 ( );
FILL FILL_2_OAI21X1_855 ( );
FILL FILL_0_BUFX2_684 ( );
FILL FILL_1_BUFX2_684 ( );
FILL FILL_0_BUFX2_305 ( );
FILL FILL_1_BUFX2_305 ( );
FILL FILL_0_BUFX2_652 ( );
FILL FILL_1_BUFX2_652 ( );
FILL FILL_0_NAND2X1_372 ( );
FILL FILL_1_NAND2X1_372 ( );
FILL FILL_0_DFFPOSX1_15 ( );
FILL FILL_1_DFFPOSX1_15 ( );
FILL FILL_2_DFFPOSX1_15 ( );
FILL FILL_3_DFFPOSX1_15 ( );
FILL FILL_4_DFFPOSX1_15 ( );
FILL FILL_5_DFFPOSX1_15 ( );
FILL FILL_0_NAND2X1_693 ( );
FILL FILL_0_OAI21X1_1625 ( );
FILL FILL_1_OAI21X1_1625 ( );
FILL FILL_2_OAI21X1_1625 ( );
FILL FILL_0_NAND2X1_661 ( );
FILL FILL_1_NAND2X1_661 ( );
FILL FILL_0_OAI21X1_1592 ( );
FILL FILL_1_OAI21X1_1592 ( );
FILL FILL_0_DFFPOSX1_1015 ( );
FILL FILL_1_DFFPOSX1_1015 ( );
FILL FILL_2_DFFPOSX1_1015 ( );
FILL FILL_3_DFFPOSX1_1015 ( );
FILL FILL_4_DFFPOSX1_1015 ( );
FILL FILL_5_DFFPOSX1_1015 ( );
FILL FILL_0_BUFX2_748 ( );
FILL FILL_0_OAI21X1_262 ( );
FILL FILL_1_OAI21X1_262 ( );
FILL FILL_0_BUFX2_205 ( );
FILL FILL_1_BUFX2_205 ( );
FILL FILL_0_BUFX2_504 ( );
FILL FILL_1_BUFX2_504 ( );
FILL FILL_0_DFFPOSX1_185 ( );
FILL FILL_1_DFFPOSX1_185 ( );
FILL FILL_2_DFFPOSX1_185 ( );
FILL FILL_3_DFFPOSX1_185 ( );
FILL FILL_4_DFFPOSX1_185 ( );
FILL FILL_5_DFFPOSX1_185 ( );
FILL FILL_6_DFFPOSX1_185 ( );
FILL FILL_0_BUFX2_1027 ( );
FILL FILL_1_BUFX2_1027 ( );
FILL FILL_0_BUFX4_42 ( );
FILL FILL_1_BUFX4_42 ( );
FILL FILL_0_OAI21X1_1766 ( );
FILL FILL_1_OAI21X1_1766 ( );
FILL FILL_0_OAI21X1_1767 ( );
FILL FILL_1_OAI21X1_1767 ( );
FILL FILL_0_OAI21X1_1407 ( );
FILL FILL_1_OAI21X1_1407 ( );
FILL FILL_0_OAI21X1_1388 ( );
FILL FILL_1_OAI21X1_1388 ( );
FILL FILL_0_OAI21X1_1389 ( );
FILL FILL_1_OAI21X1_1389 ( );
FILL FILL_0_INVX8_7 ( );
FILL FILL_1_INVX8_7 ( );
FILL FILL_0_CLKBUF1_31 ( );
FILL FILL_1_CLKBUF1_31 ( );
FILL FILL_2_CLKBUF1_31 ( );
FILL FILL_3_CLKBUF1_31 ( );
FILL FILL_4_CLKBUF1_31 ( );
FILL FILL_0_OAI21X1_634 ( );
FILL FILL_1_OAI21X1_634 ( );
FILL FILL_0_NAND2X1_240 ( );
FILL FILL_1_NAND2X1_240 ( );
FILL FILL_0_BUFX4_347 ( );
FILL FILL_1_BUFX4_347 ( );
FILL FILL_0_NAND2X1_714 ( );
FILL FILL_1_NAND2X1_714 ( );
FILL FILL_0_BUFX2_633 ( );
FILL FILL_0_DFFPOSX1_534 ( );
FILL FILL_1_DFFPOSX1_534 ( );
FILL FILL_2_DFFPOSX1_534 ( );
FILL FILL_3_DFFPOSX1_534 ( );
FILL FILL_4_DFFPOSX1_534 ( );
FILL FILL_5_DFFPOSX1_534 ( );
FILL FILL_0_OAI21X1_628 ( );
FILL FILL_1_OAI21X1_628 ( );
FILL FILL_0_CLKBUF1_100 ( );
FILL FILL_1_CLKBUF1_100 ( );
FILL FILL_2_CLKBUF1_100 ( );
FILL FILL_3_CLKBUF1_100 ( );
FILL FILL_4_CLKBUF1_100 ( );
FILL FILL_0_CLKBUF1_12 ( );
FILL FILL_1_CLKBUF1_12 ( );
FILL FILL_2_CLKBUF1_12 ( );
FILL FILL_3_CLKBUF1_12 ( );
FILL FILL_4_CLKBUF1_12 ( );
FILL FILL_0_DFFPOSX1_493 ( );
FILL FILL_1_DFFPOSX1_493 ( );
FILL FILL_2_DFFPOSX1_493 ( );
FILL FILL_3_DFFPOSX1_493 ( );
FILL FILL_4_DFFPOSX1_493 ( );
FILL FILL_5_DFFPOSX1_493 ( );
FILL FILL_0_DFFPOSX1_943 ( );
FILL FILL_1_DFFPOSX1_943 ( );
FILL FILL_2_DFFPOSX1_943 ( );
FILL FILL_3_DFFPOSX1_943 ( );
FILL FILL_4_DFFPOSX1_943 ( );
FILL FILL_5_DFFPOSX1_943 ( );
FILL FILL_6_DFFPOSX1_943 ( );
FILL FILL_0_BUFX4_57 ( );
FILL FILL_1_BUFX4_57 ( );
FILL FILL_0_OAI21X1_238 ( );
FILL FILL_1_OAI21X1_238 ( );
FILL FILL_0_OAI21X1_239 ( );
FILL FILL_1_OAI21X1_239 ( );
FILL FILL_0_BUFX2_512 ( );
FILL FILL_1_BUFX2_512 ( );
FILL FILL_0_BUFX4_82 ( );
FILL FILL_1_BUFX4_82 ( );
FILL FILL_0_BUFX4_328 ( );
FILL FILL_1_BUFX4_328 ( );
FILL FILL_0_OAI21X1_1248 ( );
FILL FILL_1_OAI21X1_1248 ( );
FILL FILL_0_DFFPOSX1_1000 ( );
FILL FILL_1_DFFPOSX1_1000 ( );
FILL FILL_2_DFFPOSX1_1000 ( );
FILL FILL_3_DFFPOSX1_1000 ( );
FILL FILL_4_DFFPOSX1_1000 ( );
FILL FILL_5_DFFPOSX1_1000 ( );
FILL FILL_0_OAI21X1_1575 ( );
FILL FILL_1_OAI21X1_1575 ( );
FILL FILL_0_OAI21X1_835 ( );
FILL FILL_1_OAI21X1_835 ( );
FILL FILL_0_DFFPOSX1_413 ( );
FILL FILL_1_DFFPOSX1_413 ( );
FILL FILL_2_DFFPOSX1_413 ( );
FILL FILL_3_DFFPOSX1_413 ( );
FILL FILL_4_DFFPOSX1_413 ( );
FILL FILL_5_DFFPOSX1_413 ( );
FILL FILL_0_OAI21X1_1419 ( );
FILL FILL_1_OAI21X1_1419 ( );
FILL FILL_0_NAND2X1_129 ( );
FILL FILL_0_OAI21X1_385 ( );
FILL FILL_1_OAI21X1_385 ( );
FILL FILL_2_OAI21X1_385 ( );
FILL FILL_0_NOR2X1_54 ( );
FILL FILL_1_NOR2X1_54 ( );
FILL FILL_0_BUFX2_450 ( );
FILL FILL_1_BUFX2_450 ( );
FILL FILL_0_DFFPOSX1_547 ( );
FILL FILL_1_DFFPOSX1_547 ( );
FILL FILL_2_DFFPOSX1_547 ( );
FILL FILL_3_DFFPOSX1_547 ( );
FILL FILL_4_DFFPOSX1_547 ( );
FILL FILL_5_DFFPOSX1_547 ( );
FILL FILL_0_BUFX2_425 ( );
FILL FILL_0_INVX4_27 ( );
FILL FILL_0_OAI21X1_390 ( );
FILL FILL_1_OAI21X1_390 ( );
FILL FILL_0_INVX1_5 ( );
FILL FILL_0_BUFX2_640 ( );
FILL FILL_1_BUFX2_640 ( );
FILL FILL_0_OAI21X1_1417 ( );
FILL FILL_1_OAI21X1_1417 ( );
FILL FILL_0_BUFX2_613 ( );
FILL FILL_1_BUFX2_613 ( );
FILL FILL_0_BUFX2_638 ( );
FILL FILL_0_BUFX2_404 ( );
FILL FILL_0_OAI21X1_1416 ( );
FILL FILL_1_OAI21X1_1416 ( );
FILL FILL_0_OAI21X1_1426 ( );
FILL FILL_1_OAI21X1_1426 ( );
FILL FILL_0_DFFPOSX1_823 ( );
FILL FILL_1_DFFPOSX1_823 ( );
FILL FILL_2_DFFPOSX1_823 ( );
FILL FILL_3_DFFPOSX1_823 ( );
FILL FILL_4_DFFPOSX1_823 ( );
FILL FILL_5_DFFPOSX1_823 ( );
FILL FILL_0_XNOR2X1_92 ( );
FILL FILL_1_XNOR2X1_92 ( );
FILL FILL_2_XNOR2X1_92 ( );
FILL FILL_3_XNOR2X1_92 ( );
FILL FILL_0_NAND2X1_90 ( );
FILL FILL_1_NAND2X1_90 ( );
FILL FILL_0_BUFX4_351 ( );
FILL FILL_1_BUFX4_351 ( );
FILL FILL_0_BUFX4_356 ( );
FILL FILL_1_BUFX4_356 ( );
FILL FILL_2_BUFX4_356 ( );
FILL FILL_0_CLKBUF1_59 ( );
FILL FILL_1_CLKBUF1_59 ( );
FILL FILL_2_CLKBUF1_59 ( );
FILL FILL_3_CLKBUF1_59 ( );
FILL FILL_4_CLKBUF1_59 ( );
FILL FILL_0_NAND2X1_418 ( );
FILL FILL_1_NAND2X1_418 ( );
FILL FILL_0_OAI21X1_1052 ( );
FILL FILL_1_OAI21X1_1052 ( );
FILL FILL_0_OAI21X1_1435 ( );
FILL FILL_1_OAI21X1_1435 ( );
FILL FILL_0_BUFX4_108 ( );
FILL FILL_1_BUFX4_108 ( );
FILL FILL_0_OAI21X1_1434 ( );
FILL FILL_1_OAI21X1_1434 ( );
FILL FILL_0_CLKBUF1_102 ( );
FILL FILL_1_CLKBUF1_102 ( );
FILL FILL_2_CLKBUF1_102 ( );
FILL FILL_3_CLKBUF1_102 ( );
FILL FILL_4_CLKBUF1_102 ( );
FILL FILL_0_BUFX2_977 ( );
FILL FILL_1_BUFX2_977 ( );
FILL FILL_0_OAI21X1_111 ( );
FILL FILL_1_OAI21X1_111 ( );
FILL FILL_0_BUFX2_134 ( );
FILL FILL_0_OAI21X1_110 ( );
FILL FILL_1_OAI21X1_110 ( );
FILL FILL_2_OAI21X1_110 ( );
FILL FILL_0_OAI21X1_584 ( );
FILL FILL_1_OAI21X1_584 ( );
FILL FILL_0_DFFPOSX1_515 ( );
FILL FILL_1_DFFPOSX1_515 ( );
FILL FILL_2_DFFPOSX1_515 ( );
FILL FILL_3_DFFPOSX1_515 ( );
FILL FILL_4_DFFPOSX1_515 ( );
FILL FILL_5_DFFPOSX1_515 ( );
FILL FILL_0_OAI21X1_583 ( );
FILL FILL_1_OAI21X1_583 ( );
FILL FILL_2_OAI21X1_583 ( );
FILL FILL_0_NOR2X1_134 ( );
FILL FILL_1_NOR2X1_134 ( );
FILL FILL_0_NAND2X1_731 ( );
FILL FILL_1_NAND2X1_731 ( );
FILL FILL_0_CLKBUF1_43 ( );
FILL FILL_1_CLKBUF1_43 ( );
FILL FILL_2_CLKBUF1_43 ( );
FILL FILL_3_CLKBUF1_43 ( );
FILL FILL_0_BUFX2_540 ( );
FILL FILL_0_DFFPOSX1_954 ( );
FILL FILL_1_DFFPOSX1_954 ( );
FILL FILL_2_DFFPOSX1_954 ( );
FILL FILL_3_DFFPOSX1_954 ( );
FILL FILL_4_DFFPOSX1_954 ( );
FILL FILL_5_DFFPOSX1_954 ( );
FILL FILL_6_DFFPOSX1_954 ( );
FILL FILL_0_DFFPOSX1_833 ( );
FILL FILL_1_DFFPOSX1_833 ( );
FILL FILL_2_DFFPOSX1_833 ( );
FILL FILL_3_DFFPOSX1_833 ( );
FILL FILL_4_DFFPOSX1_833 ( );
FILL FILL_5_DFFPOSX1_833 ( );
FILL FILL_0_NAND2X1_516 ( );
FILL FILL_1_NAND2X1_516 ( );
FILL FILL_0_OAI21X1_1144 ( );
FILL FILL_1_OAI21X1_1144 ( );
FILL FILL_0_BUFX4_159 ( );
FILL FILL_1_BUFX4_159 ( );
FILL FILL_0_OAI21X1_1460 ( );
FILL FILL_1_OAI21X1_1460 ( );
FILL FILL_0_BUFX4_40 ( );
FILL FILL_1_BUFX4_40 ( );
FILL FILL_2_BUFX4_40 ( );
FILL FILL_0_BUFX4_67 ( );
FILL FILL_1_BUFX4_67 ( );
FILL FILL_0_BUFX2_768 ( );
FILL FILL_0_NAND2X1_521 ( );
FILL FILL_0_OAI21X1_1146 ( );
FILL FILL_1_OAI21X1_1146 ( );
FILL FILL_0_OAI21X1_1145 ( );
FILL FILL_1_OAI21X1_1145 ( );
FILL FILL_0_OAI21X1_1737 ( );
FILL FILL_1_OAI21X1_1737 ( );
FILL FILL_0_OAI21X1_1736 ( );
FILL FILL_1_OAI21X1_1736 ( );
FILL FILL_2_OAI21X1_1736 ( );
FILL FILL_0_DFFPOSX1_964 ( );
FILL FILL_1_DFFPOSX1_964 ( );
FILL FILL_2_DFFPOSX1_964 ( );
FILL FILL_3_DFFPOSX1_964 ( );
FILL FILL_4_DFFPOSX1_964 ( );
FILL FILL_5_DFFPOSX1_964 ( );
FILL FILL_0_BUFX4_273 ( );
FILL FILL_1_BUFX4_273 ( );
FILL FILL_0_BUFX4_35 ( );
FILL FILL_1_BUFX4_35 ( );
FILL FILL_0_BUFX4_257 ( );
FILL FILL_1_BUFX4_257 ( );
FILL FILL_0_OAI21X1_286 ( );
FILL FILL_1_OAI21X1_286 ( );
FILL FILL_0_OAI21X1_1466 ( );
FILL FILL_1_OAI21X1_1466 ( );
FILL FILL_0_BUFX2_21 ( );
FILL FILL_1_BUFX2_21 ( );
FILL FILL_0_BUFX2_991 ( );
FILL FILL_1_BUFX2_991 ( );
FILL FILL_0_INVX2_73 ( );
FILL FILL_0_CLKBUF1_57 ( );
FILL FILL_1_CLKBUF1_57 ( );
FILL FILL_2_CLKBUF1_57 ( );
FILL FILL_3_CLKBUF1_57 ( );
FILL FILL_4_CLKBUF1_57 ( );
FILL FILL_0_BUFX2_153 ( );
FILL FILL_1_BUFX2_153 ( );
FILL FILL_0_NOR2X1_146 ( );
FILL FILL_1_NOR2X1_146 ( );
FILL FILL_0_OAI21X1_1150 ( );
FILL FILL_1_OAI21X1_1150 ( );
FILL FILL_0_OAI21X1_1149 ( );
FILL FILL_1_OAI21X1_1149 ( );
FILL FILL_0_OAI21X1_74 ( );
FILL FILL_1_OAI21X1_74 ( );
FILL FILL_0_NAND2X1_530 ( );
FILL FILL_1_NAND2X1_530 ( );
FILL FILL_0_OAI21X1_1153 ( );
FILL FILL_1_OAI21X1_1153 ( );
FILL FILL_0_NOR2X1_147 ( );
FILL FILL_1_NOR2X1_147 ( );
FILL FILL_0_OAI21X1_1170 ( );
FILL FILL_1_OAI21X1_1170 ( );
FILL FILL_0_NAND2X1_551 ( );
FILL FILL_1_NAND2X1_551 ( );
FILL FILL_0_INVX2_74 ( );
FILL FILL_0_OAI21X1_1068 ( );
FILL FILL_1_OAI21X1_1068 ( );
FILL FILL_0_NAND2X1_434 ( );
FILL FILL_0_DFFPOSX1_776 ( );
FILL FILL_1_DFFPOSX1_776 ( );
FILL FILL_2_DFFPOSX1_776 ( );
FILL FILL_3_DFFPOSX1_776 ( );
FILL FILL_4_DFFPOSX1_776 ( );
FILL FILL_5_DFFPOSX1_776 ( );
FILL FILL_6_DFFPOSX1_776 ( );
FILL FILL_0_CLKBUF1_21 ( );
FILL FILL_1_CLKBUF1_21 ( );
FILL FILL_2_CLKBUF1_21 ( );
FILL FILL_3_CLKBUF1_21 ( );
FILL FILL_4_CLKBUF1_21 ( );
FILL FILL_0_OAI21X1_1478 ( );
FILL FILL_1_OAI21X1_1478 ( );
FILL FILL_2_OAI21X1_1478 ( );
FILL FILL_0_OAI21X1_1479 ( );
FILL FILL_1_OAI21X1_1479 ( );
FILL FILL_0_DFFPOSX1_856 ( );
FILL FILL_1_DFFPOSX1_856 ( );
FILL FILL_2_DFFPOSX1_856 ( );
FILL FILL_3_DFFPOSX1_856 ( );
FILL FILL_4_DFFPOSX1_856 ( );
FILL FILL_5_DFFPOSX1_856 ( );
FILL FILL_6_DFFPOSX1_856 ( );
FILL FILL_0_OAI21X1_1475 ( );
FILL FILL_1_OAI21X1_1475 ( );
FILL FILL_0_OAI21X1_1474 ( );
FILL FILL_1_OAI21X1_1474 ( );
FILL FILL_0_DFFPOSX1_855 ( );
FILL FILL_1_DFFPOSX1_855 ( );
FILL FILL_2_DFFPOSX1_855 ( );
FILL FILL_3_DFFPOSX1_855 ( );
FILL FILL_4_DFFPOSX1_855 ( );
FILL FILL_5_DFFPOSX1_855 ( );
FILL FILL_0_OAI21X1_1294 ( );
FILL FILL_1_OAI21X1_1294 ( );
FILL FILL_0_DFFPOSX1_903 ( );
FILL FILL_1_DFFPOSX1_903 ( );
FILL FILL_2_DFFPOSX1_903 ( );
FILL FILL_3_DFFPOSX1_903 ( );
FILL FILL_4_DFFPOSX1_903 ( );
FILL FILL_5_DFFPOSX1_903 ( );
FILL FILL_0_OAI21X1_1293 ( );
FILL FILL_1_OAI21X1_1293 ( );
FILL FILL_2_OAI21X1_1293 ( );
FILL FILL_0_BUFX4_140 ( );
FILL FILL_1_BUFX4_140 ( );
FILL FILL_0_OAI21X1_980 ( );
FILL FILL_1_OAI21X1_980 ( );
FILL FILL_2_OAI21X1_980 ( );
FILL FILL_0_BUFX2_383 ( );
FILL FILL_1_BUFX2_383 ( );
FILL FILL_0_CLKBUF1_42 ( );
FILL FILL_1_CLKBUF1_42 ( );
FILL FILL_2_CLKBUF1_42 ( );
FILL FILL_3_CLKBUF1_42 ( );
FILL FILL_4_CLKBUF1_42 ( );
FILL FILL_0_DFFPOSX1_56 ( );
FILL FILL_1_DFFPOSX1_56 ( );
FILL FILL_2_DFFPOSX1_56 ( );
FILL FILL_3_DFFPOSX1_56 ( );
FILL FILL_4_DFFPOSX1_56 ( );
FILL FILL_5_DFFPOSX1_56 ( );
FILL FILL_0_BUFX2_258 ( );
FILL FILL_1_BUFX2_258 ( );
FILL FILL_0_OAI21X1_1686 ( );
FILL FILL_1_OAI21X1_1686 ( );
FILL FILL_2_OAI21X1_1686 ( );
FILL FILL_0_OAI21X1_1687 ( );
FILL FILL_1_OAI21X1_1687 ( );
FILL FILL_0_OAI21X1_1666 ( );
FILL FILL_1_OAI21X1_1666 ( );
FILL FILL_2_OAI21X1_1666 ( );
FILL FILL_0_DFFPOSX1_123 ( );
FILL FILL_1_DFFPOSX1_123 ( );
FILL FILL_2_DFFPOSX1_123 ( );
FILL FILL_3_DFFPOSX1_123 ( );
FILL FILL_4_DFFPOSX1_123 ( );
FILL FILL_5_DFFPOSX1_123 ( );
FILL FILL_0_OAI21X1_1797 ( );
FILL FILL_1_OAI21X1_1797 ( );
FILL FILL_2_OAI21X1_1797 ( );
FILL FILL_0_NAND2X1_738 ( );
FILL FILL_0_OAI21X1_1665 ( );
FILL FILL_1_OAI21X1_1665 ( );
FILL FILL_0_OAI21X1_1664 ( );
FILL FILL_1_OAI21X1_1664 ( );
FILL FILL_0_DFFPOSX1_45 ( );
FILL FILL_1_DFFPOSX1_45 ( );
FILL FILL_2_DFFPOSX1_45 ( );
FILL FILL_3_DFFPOSX1_45 ( );
FILL FILL_4_DFFPOSX1_45 ( );
FILL FILL_5_DFFPOSX1_45 ( );
FILL FILL_0_OAI21X1_910 ( );
FILL FILL_1_OAI21X1_910 ( );
FILL FILL_0_OAI21X1_911 ( );
FILL FILL_1_OAI21X1_911 ( );
FILL FILL_0_DFFPOSX1_681 ( );
FILL FILL_1_DFFPOSX1_681 ( );
FILL FILL_2_DFFPOSX1_681 ( );
FILL FILL_3_DFFPOSX1_681 ( );
FILL FILL_4_DFFPOSX1_681 ( );
FILL FILL_5_DFFPOSX1_681 ( );
FILL FILL_6_DFFPOSX1_681 ( );
FILL FILL_0_BUFX2_793 ( );
FILL FILL_1_BUFX2_793 ( );
FILL FILL_0_BUFX2_792 ( );
FILL FILL_0_BUFX2_264 ( );
FILL FILL_0_BUFX2_744 ( );
FILL FILL_1_BUFX2_744 ( );
FILL FILL_0_DFFPOSX1_632 ( );
FILL FILL_1_DFFPOSX1_632 ( );
FILL FILL_2_DFFPOSX1_632 ( );
FILL FILL_3_DFFPOSX1_632 ( );
FILL FILL_4_DFFPOSX1_632 ( );
FILL FILL_5_DFFPOSX1_632 ( );
FILL FILL_0_OAI21X1_860 ( );
FILL FILL_1_OAI21X1_860 ( );
FILL FILL_0_INVX1_61 ( );
FILL FILL_0_INVX2_177 ( );
FILL FILL_0_INVX1_78 ( );
FILL FILL_0_OAI21X1_877 ( );
FILL FILL_1_OAI21X1_877 ( );
FILL FILL_0_NAND2X1_371 ( );
FILL FILL_1_NAND2X1_371 ( );
FILL FILL_0_NAND2X1_671 ( );
FILL FILL_1_NAND2X1_671 ( );
FILL FILL_0_DFFPOSX1_649 ( );
FILL FILL_1_DFFPOSX1_649 ( );
FILL FILL_2_DFFPOSX1_649 ( );
FILL FILL_3_DFFPOSX1_649 ( );
FILL FILL_4_DFFPOSX1_649 ( );
FILL FILL_5_DFFPOSX1_649 ( );
FILL FILL_0_BUFX4_211 ( );
FILL FILL_1_BUFX4_211 ( );
FILL FILL_0_BUFX2_994 ( );
FILL FILL_1_BUFX2_994 ( );
FILL FILL_0_OAI21X1_263 ( );
FILL FILL_1_OAI21X1_263 ( );
FILL FILL_0_DFFPOSX1_323 ( );
FILL FILL_1_DFFPOSX1_323 ( );
FILL FILL_2_DFFPOSX1_323 ( );
FILL FILL_3_DFFPOSX1_323 ( );
FILL FILL_4_DFFPOSX1_323 ( );
FILL FILL_5_DFFPOSX1_323 ( );
FILL FILL_6_DFFPOSX1_323 ( );
FILL FILL_0_BUFX2_766 ( );
FILL FILL_0_DFFPOSX1_89 ( );
FILL FILL_1_DFFPOSX1_89 ( );
FILL FILL_2_DFFPOSX1_89 ( );
FILL FILL_3_DFFPOSX1_89 ( );
FILL FILL_4_DFFPOSX1_89 ( );
FILL FILL_5_DFFPOSX1_89 ( );
FILL FILL_6_DFFPOSX1_89 ( );
FILL FILL_0_BUFX4_75 ( );
FILL FILL_1_BUFX4_75 ( );
FILL FILL_0_BUFX4_70 ( );
FILL FILL_1_BUFX4_70 ( );
FILL FILL_0_BUFX4_269 ( );
FILL FILL_1_BUFX4_269 ( );
FILL FILL_0_DFFPOSX1_748 ( );
FILL FILL_1_DFFPOSX1_748 ( );
FILL FILL_2_DFFPOSX1_748 ( );
FILL FILL_3_DFFPOSX1_748 ( );
FILL FILL_4_DFFPOSX1_748 ( );
FILL FILL_5_DFFPOSX1_748 ( );
FILL FILL_6_DFFPOSX1_748 ( );
FILL FILL_0_NAND2X1_406 ( );
FILL FILL_1_NAND2X1_406 ( );
FILL FILL_0_OAI21X1_1040 ( );
FILL FILL_1_OAI21X1_1040 ( );
FILL FILL_0_DFFPOSX1_944 ( );
FILL FILL_1_DFFPOSX1_944 ( );
FILL FILL_2_DFFPOSX1_944 ( );
FILL FILL_3_DFFPOSX1_944 ( );
FILL FILL_4_DFFPOSX1_944 ( );
FILL FILL_5_DFFPOSX1_944 ( );
FILL FILL_0_OAI21X1_1408 ( );
FILL FILL_1_OAI21X1_1408 ( );
FILL FILL_0_OAI21X1_626 ( );
FILL FILL_1_OAI21X1_626 ( );
FILL FILL_0_DFFPOSX1_750 ( );
FILL FILL_1_DFFPOSX1_750 ( );
FILL FILL_2_DFFPOSX1_750 ( );
FILL FILL_3_DFFPOSX1_750 ( );
FILL FILL_4_DFFPOSX1_750 ( );
FILL FILL_5_DFFPOSX1_750 ( );
FILL FILL_6_DFFPOSX1_750 ( );
FILL FILL_0_OAI21X1_1406 ( );
FILL FILL_1_OAI21X1_1406 ( );
FILL FILL_0_OAI21X1_1393 ( );
FILL FILL_1_OAI21X1_1393 ( );
FILL FILL_0_XNOR2X1_90 ( );
FILL FILL_1_XNOR2X1_90 ( );
FILL FILL_2_XNOR2X1_90 ( );
FILL FILL_3_XNOR2X1_90 ( );
FILL FILL_0_BUFX4_29 ( );
FILL FILL_1_BUFX4_29 ( );
FILL FILL_0_INVX1_219 ( );
FILL FILL_0_NOR2X1_217 ( );
FILL FILL_1_NOR2X1_217 ( );
FILL FILL_0_NOR2X1_216 ( );
FILL FILL_0_OAI21X1_1409 ( );
FILL FILL_1_OAI21X1_1409 ( );
FILL FILL_0_OAI21X1_1410 ( );
FILL FILL_1_OAI21X1_1410 ( );
FILL FILL_2_OAI21X1_1410 ( );
FILL FILL_0_OAI21X1_1405 ( );
FILL FILL_1_OAI21X1_1405 ( );
FILL FILL_2_OAI21X1_1405 ( );
FILL FILL_0_INVX4_50 ( );
FILL FILL_1_INVX4_50 ( );
FILL FILL_0_OAI21X1_1404 ( );
FILL FILL_1_OAI21X1_1404 ( );
FILL FILL_0_NAND2X1_624 ( );
FILL FILL_1_NAND2X1_624 ( );
FILL FILL_0_DFFPOSX1_311 ( );
FILL FILL_1_DFFPOSX1_311 ( );
FILL FILL_2_DFFPOSX1_311 ( );
FILL FILL_3_DFFPOSX1_311 ( );
FILL FILL_4_DFFPOSX1_311 ( );
FILL FILL_5_DFFPOSX1_311 ( );
FILL FILL_0_BUFX2_135 ( );
FILL FILL_1_BUFX2_135 ( );
FILL FILL_0_BUFX2_632 ( );
FILL FILL_1_BUFX2_632 ( );
FILL FILL_0_OAI21X1_1249 ( );
FILL FILL_1_OAI21X1_1249 ( );
FILL FILL_0_BUFX4_146 ( );
FILL FILL_1_BUFX4_146 ( );
FILL FILL_0_NAND2X1_304 ( );
FILL FILL_1_NAND2X1_304 ( );
FILL FILL_0_INVX4_25 ( );
FILL FILL_1_INVX4_25 ( );
FILL FILL_0_DFFPOSX1_949 ( );
FILL FILL_1_DFFPOSX1_949 ( );
FILL FILL_2_DFFPOSX1_949 ( );
FILL FILL_3_DFFPOSX1_949 ( );
FILL FILL_4_DFFPOSX1_949 ( );
FILL FILL_5_DFFPOSX1_949 ( );
FILL FILL_6_DFFPOSX1_949 ( );
FILL FILL_0_OAI21X1_1423 ( );
FILL FILL_1_OAI21X1_1423 ( );
FILL FILL_0_OAI21X1_1424 ( );
FILL FILL_1_OAI21X1_1424 ( );
FILL FILL_2_OAI21X1_1424 ( );
FILL FILL_0_DFFPOSX1_948 ( );
FILL FILL_1_DFFPOSX1_948 ( );
FILL FILL_2_DFFPOSX1_948 ( );
FILL FILL_3_DFFPOSX1_948 ( );
FILL FILL_4_DFFPOSX1_948 ( );
FILL FILL_5_DFFPOSX1_948 ( );
FILL FILL_0_OAI21X1_1420 ( );
FILL FILL_1_OAI21X1_1420 ( );
FILL FILL_0_CLKBUF1_29 ( );
FILL FILL_1_CLKBUF1_29 ( );
FILL FILL_2_CLKBUF1_29 ( );
FILL FILL_3_CLKBUF1_29 ( );
FILL FILL_4_CLKBUF1_29 ( );
FILL FILL_0_OAI21X1_1418 ( );
FILL FILL_1_OAI21X1_1418 ( );
FILL FILL_0_DFFPOSX1_418 ( );
FILL FILL_1_DFFPOSX1_418 ( );
FILL FILL_2_DFFPOSX1_418 ( );
FILL FILL_3_DFFPOSX1_418 ( );
FILL FILL_4_DFFPOSX1_418 ( );
FILL FILL_5_DFFPOSX1_418 ( );
FILL FILL_0_NAND2X1_306 ( );
FILL FILL_1_NAND2X1_306 ( );
FILL FILL_0_DFFPOSX1_947 ( );
FILL FILL_1_DFFPOSX1_947 ( );
FILL FILL_2_DFFPOSX1_947 ( );
FILL FILL_3_DFFPOSX1_947 ( );
FILL FILL_4_DFFPOSX1_947 ( );
FILL FILL_5_DFFPOSX1_947 ( );
FILL FILL_6_DFFPOSX1_947 ( );
FILL FILL_0_BUFX4_150 ( );
FILL FILL_1_BUFX4_150 ( );
FILL FILL_2_BUFX4_150 ( );
FILL FILL_0_OAI21X1_1425 ( );
FILL FILL_1_OAI21X1_1425 ( );
FILL FILL_2_OAI21X1_1425 ( );
FILL FILL_0_INVX1_220 ( );
FILL FILL_0_OAI21X1_1427 ( );
FILL FILL_1_OAI21X1_1427 ( );
FILL FILL_0_DFFPOSX1_950 ( );
FILL FILL_1_DFFPOSX1_950 ( );
FILL FILL_2_DFFPOSX1_950 ( );
FILL FILL_3_DFFPOSX1_950 ( );
FILL FILL_4_DFFPOSX1_950 ( );
FILL FILL_5_DFFPOSX1_950 ( );
FILL FILL_0_XNOR2X1_57 ( );
FILL FILL_1_XNOR2X1_57 ( );
FILL FILL_2_XNOR2X1_57 ( );
FILL FILL_3_XNOR2X1_57 ( );
FILL FILL_0_OAI21X1_1129 ( );
FILL FILL_1_OAI21X1_1129 ( );
FILL FILL_0_NOR2X1_131 ( );
FILL FILL_0_NAND2X1_497 ( );
FILL FILL_0_NOR2X1_133 ( );
FILL FILL_0_NAND2X1_501 ( );
FILL FILL_1_NAND2X1_501 ( );
FILL FILL_0_OR2X2_16 ( );
FILL FILL_1_OR2X2_16 ( );
FILL FILL_2_OR2X2_16 ( );
FILL FILL_0_DFFPOSX1_953 ( );
FILL FILL_1_DFFPOSX1_953 ( );
FILL FILL_2_DFFPOSX1_953 ( );
FILL FILL_3_DFFPOSX1_953 ( );
FILL FILL_4_DFFPOSX1_953 ( );
FILL FILL_5_DFFPOSX1_953 ( );
FILL FILL_0_NOR2X1_132 ( );
FILL FILL_0_INVX1_221 ( );
FILL FILL_0_XNOR2X1_58 ( );
FILL FILL_1_XNOR2X1_58 ( );
FILL FILL_2_XNOR2X1_58 ( );
FILL FILL_0_DFFPOSX1_825 ( );
FILL FILL_1_DFFPOSX1_825 ( );
FILL FILL_2_DFFPOSX1_825 ( );
FILL FILL_3_DFFPOSX1_825 ( );
FILL FILL_4_DFFPOSX1_825 ( );
FILL FILL_5_DFFPOSX1_825 ( );
FILL FILL_0_NAND2X1_498 ( );
FILL FILL_1_NAND2X1_498 ( );
FILL FILL_0_DFFPOSX1_292 ( );
FILL FILL_1_DFFPOSX1_292 ( );
FILL FILL_2_DFFPOSX1_292 ( );
FILL FILL_3_DFFPOSX1_292 ( );
FILL FILL_4_DFFPOSX1_292 ( );
FILL FILL_5_DFFPOSX1_292 ( );
FILL FILL_0_BUFX4_149 ( );
FILL FILL_1_BUFX4_149 ( );
FILL FILL_0_OAI21X1_1774 ( );
FILL FILL_1_OAI21X1_1774 ( );
FILL FILL_0_DFFPOSX1_100 ( );
FILL FILL_1_DFFPOSX1_100 ( );
FILL FILL_2_DFFPOSX1_100 ( );
FILL FILL_3_DFFPOSX1_100 ( );
FILL FILL_4_DFFPOSX1_100 ( );
FILL FILL_5_DFFPOSX1_100 ( );
FILL FILL_6_DFFPOSX1_100 ( );
FILL FILL_0_DFFPOSX1_60 ( );
FILL FILL_1_DFFPOSX1_60 ( );
FILL FILL_2_DFFPOSX1_60 ( );
FILL FILL_3_DFFPOSX1_60 ( );
FILL FILL_4_DFFPOSX1_60 ( );
FILL FILL_5_DFFPOSX1_60 ( );
FILL FILL_0_OAI21X1_65 ( );
FILL FILL_1_OAI21X1_65 ( );
FILL FILL_0_DFFPOSX1_221 ( );
FILL FILL_1_DFFPOSX1_221 ( );
FILL FILL_2_DFFPOSX1_221 ( );
FILL FILL_3_DFFPOSX1_221 ( );
FILL FILL_4_DFFPOSX1_221 ( );
FILL FILL_5_DFFPOSX1_221 ( );
FILL FILL_6_DFFPOSX1_221 ( );
FILL FILL_0_DFFPOSX1_63 ( );
FILL FILL_1_DFFPOSX1_63 ( );
FILL FILL_2_DFFPOSX1_63 ( );
FILL FILL_3_DFFPOSX1_63 ( );
FILL FILL_4_DFFPOSX1_63 ( );
FILL FILL_5_DFFPOSX1_63 ( );
FILL FILL_6_DFFPOSX1_63 ( );
FILL FILL_0_DFFPOSX1_136 ( );
FILL FILL_1_DFFPOSX1_136 ( );
FILL FILL_2_DFFPOSX1_136 ( );
FILL FILL_3_DFFPOSX1_136 ( );
FILL FILL_4_DFFPOSX1_136 ( );
FILL FILL_5_DFFPOSX1_136 ( );
FILL FILL_0_OAI21X1_1810 ( );
FILL FILL_1_OAI21X1_1810 ( );
FILL FILL_2_OAI21X1_1810 ( );
FILL FILL_0_CLKBUF1_16 ( );
FILL FILL_1_CLKBUF1_16 ( );
FILL FILL_2_CLKBUF1_16 ( );
FILL FILL_3_CLKBUF1_16 ( );
FILL FILL_4_CLKBUF1_16 ( );
FILL FILL_0_BUFX4_106 ( );
FILL FILL_1_BUFX4_106 ( );
FILL FILL_0_BUFX4_279 ( );
FILL FILL_1_BUFX4_279 ( );
FILL FILL_0_INVX1_182 ( );
FILL FILL_0_OAI21X1_1103 ( );
FILL FILL_1_OAI21X1_1103 ( );
FILL FILL_0_NAND2X1_469 ( );
FILL FILL_1_NAND2X1_469 ( );
FILL FILL_0_BUFX2_963 ( );
FILL FILL_0_BUFX2_211 ( );
FILL FILL_1_BUFX2_211 ( );
FILL FILL_0_OAI21X1_1584 ( );
FILL FILL_1_OAI21X1_1584 ( );
FILL FILL_0_NAND2X1_653 ( );
FILL FILL_1_NAND2X1_653 ( );
FILL FILL_0_DFFPOSX1_1007 ( );
FILL FILL_1_DFFPOSX1_1007 ( );
FILL FILL_2_DFFPOSX1_1007 ( );
FILL FILL_3_DFFPOSX1_1007 ( );
FILL FILL_4_DFFPOSX1_1007 ( );
FILL FILL_5_DFFPOSX1_1007 ( );
FILL FILL_0_OAI21X1_1465 ( );
FILL FILL_1_OAI21X1_1465 ( );
FILL FILL_0_BUFX2_750 ( );
FILL FILL_0_BUFX2_150 ( );
FILL FILL_0_OAI21X1_1759 ( );
FILL FILL_1_OAI21X1_1759 ( );
FILL FILL_0_DFFPOSX1_92 ( );
FILL FILL_1_DFFPOSX1_92 ( );
FILL FILL_2_DFFPOSX1_92 ( );
FILL FILL_3_DFFPOSX1_92 ( );
FILL FILL_4_DFFPOSX1_92 ( );
FILL FILL_5_DFFPOSX1_92 ( );
FILL FILL_0_NAND2X1_525 ( );
FILL FILL_0_DFFPOSX1_837 ( );
FILL FILL_1_DFFPOSX1_837 ( );
FILL FILL_2_DFFPOSX1_837 ( );
FILL FILL_3_DFFPOSX1_837 ( );
FILL FILL_4_DFFPOSX1_837 ( );
FILL FILL_5_DFFPOSX1_837 ( );
FILL FILL_6_DFFPOSX1_837 ( );
FILL FILL_0_DFFPOSX1_335 ( );
FILL FILL_1_DFFPOSX1_335 ( );
FILL FILL_2_DFFPOSX1_335 ( );
FILL FILL_3_DFFPOSX1_335 ( );
FILL FILL_4_DFFPOSX1_335 ( );
FILL FILL_5_DFFPOSX1_335 ( );
FILL FILL_0_OAI21X1_1744 ( );
FILL FILL_1_OAI21X1_1744 ( );
FILL FILL_0_OAI21X1_287 ( );
FILL FILL_1_OAI21X1_287 ( );
FILL FILL_0_BUFX4_55 ( );
FILL FILL_1_BUFX4_55 ( );
FILL FILL_0_BUFX4_50 ( );
FILL FILL_1_BUFX4_50 ( );
FILL FILL_0_OAI21X1_1155 ( );
FILL FILL_1_OAI21X1_1155 ( );
FILL FILL_0_DFFPOSX1_838 ( );
FILL FILL_1_DFFPOSX1_838 ( );
FILL FILL_2_DFFPOSX1_838 ( );
FILL FILL_3_DFFPOSX1_838 ( );
FILL FILL_4_DFFPOSX1_838 ( );
FILL FILL_5_DFFPOSX1_838 ( );
FILL FILL_0_NOR2X1_148 ( );
FILL FILL_0_DFFPOSX1_851 ( );
FILL FILL_1_DFFPOSX1_851 ( );
FILL FILL_2_DFFPOSX1_851 ( );
FILL FILL_3_DFFPOSX1_851 ( );
FILL FILL_4_DFFPOSX1_851 ( );
FILL FILL_5_DFFPOSX1_851 ( );
FILL FILL_0_BUFX4_301 ( );
FILL FILL_1_BUFX4_301 ( );
FILL FILL_0_BUFX2_90 ( );
FILL FILL_0_BUFX4_293 ( );
FILL FILL_1_BUFX4_293 ( );
FILL FILL_0_DFFPOSX1_968 ( );
FILL FILL_1_DFFPOSX1_968 ( );
FILL FILL_2_DFFPOSX1_968 ( );
FILL FILL_3_DFFPOSX1_968 ( );
FILL FILL_4_DFFPOSX1_968 ( );
FILL FILL_5_DFFPOSX1_968 ( );
FILL FILL_0_BUFX4_341 ( );
FILL FILL_1_BUFX4_341 ( );
FILL FILL_0_OAI21X1_1067 ( );
FILL FILL_1_OAI21X1_1067 ( );
FILL FILL_2_OAI21X1_1067 ( );
FILL FILL_0_DFFPOSX1_775 ( );
FILL FILL_1_DFFPOSX1_775 ( );
FILL FILL_2_DFFPOSX1_775 ( );
FILL FILL_3_DFFPOSX1_775 ( );
FILL FILL_4_DFFPOSX1_775 ( );
FILL FILL_5_DFFPOSX1_775 ( );
FILL FILL_0_DFFPOSX1_333 ( );
FILL FILL_1_DFFPOSX1_333 ( );
FILL FILL_2_DFFPOSX1_333 ( );
FILL FILL_3_DFFPOSX1_333 ( );
FILL FILL_4_DFFPOSX1_333 ( );
FILL FILL_5_DFFPOSX1_333 ( );
FILL FILL_0_OAI21X1_981 ( );
FILL FILL_1_OAI21X1_981 ( );
FILL FILL_0_DFFPOSX1_967 ( );
FILL FILL_1_DFFPOSX1_967 ( );
FILL FILL_2_DFFPOSX1_967 ( );
FILL FILL_3_DFFPOSX1_967 ( );
FILL FILL_4_DFFPOSX1_967 ( );
FILL FILL_5_DFFPOSX1_967 ( );
FILL FILL_6_DFFPOSX1_967 ( );
FILL FILL_0_BUFX4_128 ( );
FILL FILL_1_BUFX4_128 ( );
FILL FILL_0_BUFX4_272 ( );
FILL FILL_1_BUFX4_272 ( );
FILL FILL_0_DFFPOSX1_149 ( );
FILL FILL_1_DFFPOSX1_149 ( );
FILL FILL_2_DFFPOSX1_149 ( );
FILL FILL_3_DFFPOSX1_149 ( );
FILL FILL_4_DFFPOSX1_149 ( );
FILL FILL_5_DFFPOSX1_149 ( );
FILL FILL_0_BUFX4_103 ( );
FILL FILL_1_BUFX4_103 ( );
FILL FILL_0_OAI21X1_1667 ( );
FILL FILL_1_OAI21X1_1667 ( );
FILL FILL_0_DFFPOSX1_46 ( );
FILL FILL_1_DFFPOSX1_46 ( );
FILL FILL_2_DFFPOSX1_46 ( );
FILL FILL_3_DFFPOSX1_46 ( );
FILL FILL_4_DFFPOSX1_46 ( );
FILL FILL_5_DFFPOSX1_46 ( );
FILL FILL_6_DFFPOSX1_46 ( );
FILL FILL_0_BUFX2_171 ( );
FILL FILL_1_BUFX2_171 ( );
FILL FILL_0_OAI21X1_31 ( );
FILL FILL_1_OAI21X1_31 ( );
FILL FILL_0_NAND2X1_31 ( );
FILL FILL_1_NAND2X1_31 ( );
FILL FILL_0_INVX1_145 ( );
FILL FILL_0_BUFX2_154 ( );
FILL FILL_1_BUFX2_154 ( );
FILL FILL_0_DFFPOSX1_186 ( );
FILL FILL_1_DFFPOSX1_186 ( );
FILL FILL_2_DFFPOSX1_186 ( );
FILL FILL_3_DFFPOSX1_186 ( );
FILL FILL_4_DFFPOSX1_186 ( );
FILL FILL_5_DFFPOSX1_186 ( );
FILL FILL_0_OAI21X1_30 ( );
FILL FILL_1_OAI21X1_30 ( );
FILL FILL_0_NAND2X1_30 ( );
FILL FILL_1_NAND2X1_30 ( );
FILL FILL_0_OAI21X1_1624 ( );
FILL FILL_1_OAI21X1_1624 ( );
FILL FILL_0_DFFPOSX1_14 ( );
FILL FILL_1_DFFPOSX1_14 ( );
FILL FILL_2_DFFPOSX1_14 ( );
FILL FILL_3_DFFPOSX1_14 ( );
FILL FILL_4_DFFPOSX1_14 ( );
FILL FILL_5_DFFPOSX1_14 ( );
FILL FILL_0_INVX2_168 ( );
FILL FILL_0_NAND2X1_343 ( );
FILL FILL_0_NAND2X1_354 ( );
FILL FILL_1_NAND2X1_354 ( );
FILL FILL_0_BUFX2_294 ( );
FILL FILL_1_BUFX2_294 ( );
FILL FILL_0_BUFX2_663 ( );
FILL FILL_1_BUFX2_663 ( );
FILL FILL_0_INVX2_128 ( );
FILL FILL_0_DFFPOSX1_1025 ( );
FILL FILL_1_DFFPOSX1_1025 ( );
FILL FILL_2_DFFPOSX1_1025 ( );
FILL FILL_3_DFFPOSX1_1025 ( );
FILL FILL_4_DFFPOSX1_1025 ( );
FILL FILL_5_DFFPOSX1_1025 ( );
FILL FILL_6_DFFPOSX1_1025 ( );
FILL FILL_0_OAI21X1_1602 ( );
FILL FILL_1_OAI21X1_1602 ( );
FILL FILL_0_DFFPOSX1_737 ( );
FILL FILL_1_DFFPOSX1_737 ( );
FILL FILL_2_DFFPOSX1_737 ( );
FILL FILL_3_DFFPOSX1_737 ( );
FILL FILL_4_DFFPOSX1_737 ( );
FILL FILL_5_DFFPOSX1_737 ( );
FILL FILL_6_DFFPOSX1_737 ( );
FILL FILL_0_NAND2X1_703 ( );
FILL FILL_1_NAND2X1_703 ( );
FILL FILL_0_OAI21X1_1635 ( );
FILL FILL_1_OAI21X1_1635 ( );
FILL FILL_0_DFFPOSX1_25 ( );
FILL FILL_1_DFFPOSX1_25 ( );
FILL FILL_2_DFFPOSX1_25 ( );
FILL FILL_3_DFFPOSX1_25 ( );
FILL FILL_4_DFFPOSX1_25 ( );
FILL FILL_5_DFFPOSX1_25 ( );
FILL FILL_0_BUFX2_855 ( );
FILL FILL_1_BUFX2_855 ( );
FILL FILL_0_BUFX4_352 ( );
FILL FILL_1_BUFX4_352 ( );
FILL FILL_0_OAI21X1_1753 ( );
FILL FILL_1_OAI21X1_1753 ( );
FILL FILL_0_DFFPOSX1_47 ( );
FILL FILL_1_DFFPOSX1_47 ( );
FILL FILL_2_DFFPOSX1_47 ( );
FILL FILL_3_DFFPOSX1_47 ( );
FILL FILL_4_DFFPOSX1_47 ( );
FILL FILL_5_DFFPOSX1_47 ( );
FILL FILL_0_OAI21X1_1669 ( );
FILL FILL_1_OAI21X1_1669 ( );
FILL FILL_0_BUFX2_35 ( );
FILL FILL_0_BUFX2_255 ( );
FILL FILL_1_BUFX2_255 ( );
FILL FILL_0_OAI21X1_1668 ( );
FILL FILL_1_OAI21X1_1668 ( );
FILL FILL_0_BUFX2_570 ( );
FILL FILL_1_BUFX2_570 ( );
FILL FILL_0_OAI21X1_1400 ( );
FILL FILL_1_OAI21X1_1400 ( );
FILL FILL_0_BUFX2_440 ( );
FILL FILL_1_BUFX2_440 ( );
FILL FILL_0_OAI21X1_1401 ( );
FILL FILL_1_OAI21X1_1401 ( );
FILL FILL_0_DFFPOSX1_749 ( );
FILL FILL_1_DFFPOSX1_749 ( );
FILL FILL_2_DFFPOSX1_749 ( );
FILL FILL_3_DFFPOSX1_749 ( );
FILL FILL_4_DFFPOSX1_749 ( );
FILL FILL_5_DFFPOSX1_749 ( );
FILL FILL_0_DFFPOSX1_941 ( );
FILL FILL_1_DFFPOSX1_941 ( );
FILL FILL_2_DFFPOSX1_941 ( );
FILL FILL_3_DFFPOSX1_941 ( );
FILL FILL_4_DFFPOSX1_941 ( );
FILL FILL_5_DFFPOSX1_941 ( );
FILL FILL_6_DFFPOSX1_941 ( );
FILL FILL_0_NAND2X1_408 ( );
FILL FILL_0_OAI21X1_1042 ( );
FILL FILL_1_OAI21X1_1042 ( );
FILL FILL_2_OAI21X1_1042 ( );
FILL FILL_0_INVX2_57 ( );
FILL FILL_0_BUFX2_584 ( );
FILL FILL_0_OAI21X1_1392 ( );
FILL FILL_1_OAI21X1_1392 ( );
FILL FILL_2_OAI21X1_1392 ( );
FILL FILL_0_BUFX2_623 ( );
FILL FILL_0_NOR2X1_122 ( );
FILL FILL_1_NOR2X1_122 ( );
FILL FILL_0_NOR2X1_215 ( );
FILL FILL_0_OAI21X1_1112 ( );
FILL FILL_1_OAI21X1_1112 ( );
FILL FILL_0_OAI21X1_1113 ( );
FILL FILL_1_OAI21X1_1113 ( );
FILL FILL_0_OAI21X1_1402 ( );
FILL FILL_1_OAI21X1_1402 ( );
FILL FILL_0_OAI21X1_1403 ( );
FILL FILL_1_OAI21X1_1403 ( );
FILL FILL_0_OAI21X1_1115 ( );
FILL FILL_1_OAI21X1_1115 ( );
FILL FILL_2_OAI21X1_1115 ( );
FILL FILL_0_INVX1_185 ( );
FILL FILL_1_INVX1_185 ( );
FILL FILL_0_NAND2X1_476 ( );
FILL FILL_0_NAND3X1_38 ( );
FILL FILL_1_NAND3X1_38 ( );
FILL FILL_0_OAI21X1_1118 ( );
FILL FILL_1_OAI21X1_1118 ( );
FILL FILL_0_INVX2_94 ( );
FILL FILL_0_NOR2X1_123 ( );
FILL FILL_0_BUFX2_639 ( );
FILL FILL_1_BUFX2_639 ( );
FILL FILL_0_OAI21X1_1413 ( );
FILL FILL_1_OAI21X1_1413 ( );
FILL FILL_0_DFFPOSX1_541 ( );
FILL FILL_1_DFFPOSX1_541 ( );
FILL FILL_2_DFFPOSX1_541 ( );
FILL FILL_3_DFFPOSX1_541 ( );
FILL FILL_4_DFFPOSX1_541 ( );
FILL FILL_5_DFFPOSX1_541 ( );
FILL FILL_0_OAI21X1_643 ( );
FILL FILL_1_OAI21X1_643 ( );
FILL FILL_0_NAND2X1_303 ( );
FILL FILL_0_INVX2_63 ( );
FILL FILL_0_OAI21X1_645 ( );
FILL FILL_1_OAI21X1_645 ( );
FILL FILL_0_NAND2X1_648 ( );
FILL FILL_0_NAND2X1_625 ( );
FILL FILL_1_NAND2X1_625 ( );
FILL FILL_0_BUFX2_643 ( );
FILL FILL_1_BUFX2_643 ( );
FILL FILL_0_INVX2_108 ( );
FILL FILL_0_NOR2X1_218 ( );
FILL FILL_0_NOR2X1_128 ( );
FILL FILL_0_DFFPOSX1_818 ( );
FILL FILL_1_DFFPOSX1_818 ( );
FILL FILL_2_DFFPOSX1_818 ( );
FILL FILL_3_DFFPOSX1_818 ( );
FILL FILL_4_DFFPOSX1_818 ( );
FILL FILL_5_DFFPOSX1_818 ( );
FILL FILL_0_AOI21X1_60 ( );
FILL FILL_1_AOI21X1_60 ( );
FILL FILL_2_AOI21X1_60 ( );
FILL FILL_0_OAI21X1_1121 ( );
FILL FILL_1_OAI21X1_1121 ( );
FILL FILL_0_OAI21X1_1120 ( );
FILL FILL_1_OAI21X1_1120 ( );
FILL FILL_0_OAI21X1_1422 ( );
FILL FILL_1_OAI21X1_1422 ( );
FILL FILL_0_OAI21X1_1421 ( );
FILL FILL_1_OAI21X1_1421 ( );
FILL FILL_0_NAND2X1_134 ( );
FILL FILL_1_NAND2X1_134 ( );
FILL FILL_0_XNOR2X1_91 ( );
FILL FILL_1_XNOR2X1_91 ( );
FILL FILL_2_XNOR2X1_91 ( );
FILL FILL_3_XNOR2X1_91 ( );
FILL FILL_0_OAI21X1_653 ( );
FILL FILL_1_OAI21X1_653 ( );
FILL FILL_0_OAI21X1_656 ( );
FILL FILL_1_OAI21X1_656 ( );
FILL FILL_0_OAI21X1_1247 ( );
FILL FILL_1_OAI21X1_1247 ( );
FILL FILL_0_OAI21X1_1246 ( );
FILL FILL_1_OAI21X1_1246 ( );
FILL FILL_0_OAI21X1_274 ( );
FILL FILL_1_OAI21X1_274 ( );
FILL FILL_0_NAND2X1_494 ( );
FILL FILL_0_NOR2X1_130 ( );
FILL FILL_1_NOR2X1_130 ( );
FILL FILL_0_NOR2X1_219 ( );
FILL FILL_0_DFFPOSX1_248 ( );
FILL FILL_1_DFFPOSX1_248 ( );
FILL FILL_2_DFFPOSX1_248 ( );
FILL FILL_3_DFFPOSX1_248 ( );
FILL FILL_4_DFFPOSX1_248 ( );
FILL FILL_5_DFFPOSX1_248 ( );
FILL FILL_0_OAI21X1_113 ( );
FILL FILL_1_OAI21X1_113 ( );
FILL FILL_0_INVX1_186 ( );
FILL FILL_1_INVX1_186 ( );
FILL FILL_0_NAND2X1_495 ( );
FILL FILL_1_NAND2X1_495 ( );
FILL FILL_0_NAND2X1_496 ( );
FILL FILL_1_NAND2X1_496 ( );
FILL FILL_0_NOR2X1_185 ( );
FILL FILL_0_NAND2X1_500 ( );
FILL FILL_1_NAND2X1_500 ( );
FILL FILL_0_NAND3X1_52 ( );
FILL FILL_1_NAND3X1_52 ( );
FILL FILL_0_NAND2X1_626 ( );
FILL FILL_0_XNOR2X1_93 ( );
FILL FILL_1_XNOR2X1_93 ( );
FILL FILL_2_XNOR2X1_93 ( );
FILL FILL_3_XNOR2X1_93 ( );
FILL FILL_0_BUFX2_74 ( );
FILL FILL_0_XNOR2X1_59 ( );
FILL FILL_1_XNOR2X1_59 ( );
FILL FILL_2_XNOR2X1_59 ( );
FILL FILL_3_XNOR2X1_59 ( );
FILL FILL_0_OAI21X1_1131 ( );
FILL FILL_1_OAI21X1_1131 ( );
FILL FILL_0_NAND2X1_499 ( );
FILL FILL_1_NAND2X1_499 ( );
FILL FILL_0_OAI21X1_1130 ( );
FILL FILL_1_OAI21X1_1130 ( );
FILL FILL_0_DFFPOSX1_824 ( );
FILL FILL_1_DFFPOSX1_824 ( );
FILL FILL_2_DFFPOSX1_824 ( );
FILL FILL_3_DFFPOSX1_824 ( );
FILL FILL_4_DFFPOSX1_824 ( );
FILL FILL_5_DFFPOSX1_824 ( );
FILL FILL_6_DFFPOSX1_824 ( );
FILL FILL_0_OAI21X1_201 ( );
FILL FILL_1_OAI21X1_201 ( );
FILL FILL_2_OAI21X1_201 ( );
FILL FILL_0_OAI21X1_200 ( );
FILL FILL_1_OAI21X1_200 ( );
FILL FILL_0_BUFX2_481 ( );
FILL FILL_1_BUFX2_481 ( );
FILL FILL_0_BUFX4_379 ( );
FILL FILL_1_BUFX4_379 ( );
FILL FILL_0_BUFX2_546 ( );
FILL FILL_1_BUFX2_546 ( );
FILL FILL_0_NAND2X1_715 ( );
FILL FILL_1_NAND2X1_715 ( );
FILL FILL_0_BUFX4_168 ( );
FILL FILL_1_BUFX4_168 ( );
FILL FILL_0_BUFX2_785 ( );
FILL FILL_1_BUFX2_785 ( );
FILL FILL_0_BUFX2_777 ( );
FILL FILL_1_BUFX2_777 ( );
FILL FILL_0_OAI21X1_1391 ( );
FILL FILL_1_OAI21X1_1391 ( );
FILL FILL_0_OAI21X1_1695 ( );
FILL FILL_1_OAI21X1_1695 ( );
FILL FILL_0_OAI21X1_1437 ( );
FILL FILL_1_OAI21X1_1437 ( );
FILL FILL_2_OAI21X1_1437 ( );
FILL FILL_0_NAND2X1_65 ( );
FILL FILL_1_NAND2X1_65 ( );
FILL FILL_0_BUFX2_894 ( );
FILL FILL_1_BUFX2_894 ( );
FILL FILL_0_OAI21X1_1701 ( );
FILL FILL_1_OAI21X1_1701 ( );
FILL FILL_0_OAI21X1_1700 ( );
FILL FILL_1_OAI21X1_1700 ( );
FILL FILL_0_DFFPOSX1_90 ( );
FILL FILL_1_DFFPOSX1_90 ( );
FILL FILL_2_DFFPOSX1_90 ( );
FILL FILL_3_DFFPOSX1_90 ( );
FILL FILL_4_DFFPOSX1_90 ( );
FILL FILL_5_DFFPOSX1_90 ( );
FILL FILL_0_OAI21X1_1459 ( );
FILL FILL_1_OAI21X1_1459 ( );
FILL FILL_0_CLKBUF1_93 ( );
FILL FILL_1_CLKBUF1_93 ( );
FILL FILL_2_CLKBUF1_93 ( );
FILL FILL_3_CLKBUF1_93 ( );
FILL FILL_4_CLKBUF1_93 ( );
FILL FILL_0_BUFX4_36 ( );
FILL FILL_1_BUFX4_36 ( );
FILL FILL_0_NAND2X1_751 ( );
FILL FILL_0_CLKBUF1_7 ( );
FILL FILL_1_CLKBUF1_7 ( );
FILL FILL_2_CLKBUF1_7 ( );
FILL FILL_3_CLKBUF1_7 ( );
FILL FILL_4_CLKBUF1_7 ( );
FILL FILL_0_BUFX2_212 ( );
FILL FILL_0_DFFPOSX1_811 ( );
FILL FILL_1_DFFPOSX1_811 ( );
FILL FILL_2_DFFPOSX1_811 ( );
FILL FILL_3_DFFPOSX1_811 ( );
FILL FILL_4_DFFPOSX1_811 ( );
FILL FILL_5_DFFPOSX1_811 ( );
FILL FILL_6_DFFPOSX1_811 ( );
FILL FILL_0_OAI21X1_1653 ( );
FILL FILL_1_OAI21X1_1653 ( );
FILL FILL_2_OAI21X1_1653 ( );
FILL FILL_0_DFFPOSX1_39 ( );
FILL FILL_1_DFFPOSX1_39 ( );
FILL FILL_2_DFFPOSX1_39 ( );
FILL FILL_3_DFFPOSX1_39 ( );
FILL FILL_4_DFFPOSX1_39 ( );
FILL FILL_5_DFFPOSX1_39 ( );
FILL FILL_6_DFFPOSX1_39 ( );
FILL FILL_0_OAI21X1_296 ( );
FILL FILL_1_OAI21X1_296 ( );
FILL FILL_0_DFFPOSX1_773 ( );
FILL FILL_1_DFFPOSX1_773 ( );
FILL FILL_2_DFFPOSX1_773 ( );
FILL FILL_3_DFFPOSX1_773 ( );
FILL FILL_4_DFFPOSX1_773 ( );
FILL FILL_5_DFFPOSX1_773 ( );
FILL FILL_0_OAI21X1_1065 ( );
FILL FILL_1_OAI21X1_1065 ( );
FILL FILL_0_OAI21X1_1758 ( );
FILL FILL_1_OAI21X1_1758 ( );
FILL FILL_0_OAI21X1_108 ( );
FILL FILL_1_OAI21X1_108 ( );
FILL FILL_0_OAI21X1_109 ( );
FILL FILL_1_OAI21X1_109 ( );
FILL FILL_0_DFFPOSX1_246 ( );
FILL FILL_1_DFFPOSX1_246 ( );
FILL FILL_2_DFFPOSX1_246 ( );
FILL FILL_3_DFFPOSX1_246 ( );
FILL FILL_4_DFFPOSX1_246 ( );
FILL FILL_5_DFFPOSX1_246 ( );
FILL FILL_0_CLKBUF1_14 ( );
FILL FILL_1_CLKBUF1_14 ( );
FILL FILL_2_CLKBUF1_14 ( );
FILL FILL_3_CLKBUF1_14 ( );
FILL FILL_4_CLKBUF1_14 ( );
FILL FILL_0_DFFPOSX1_85 ( );
FILL FILL_1_DFFPOSX1_85 ( );
FILL FILL_2_DFFPOSX1_85 ( );
FILL FILL_3_DFFPOSX1_85 ( );
FILL FILL_4_DFFPOSX1_85 ( );
FILL FILL_5_DFFPOSX1_85 ( );
FILL FILL_6_DFFPOSX1_85 ( );
FILL FILL_0_BUFX2_214 ( );
FILL FILL_1_BUFX2_214 ( );
FILL FILL_0_BUFX2_923 ( );
FILL FILL_1_BUFX2_923 ( );
FILL FILL_0_OAI21X1_1792 ( );
FILL FILL_1_OAI21X1_1792 ( );
FILL FILL_0_OAI21X1_1156 ( );
FILL FILL_1_OAI21X1_1156 ( );
FILL FILL_0_CLKBUF1_95 ( );
FILL FILL_1_CLKBUF1_95 ( );
FILL FILL_2_CLKBUF1_95 ( );
FILL FILL_3_CLKBUF1_95 ( );
FILL FILL_0_AOI21X1_38 ( );
FILL FILL_1_AOI21X1_38 ( );
FILL FILL_0_BUFX2_89 ( );
FILL FILL_1_BUFX2_89 ( );
FILL FILL_0_NOR2X1_149 ( );
FILL FILL_1_NOR2X1_149 ( );
FILL FILL_0_OAI21X1_1154 ( );
FILL FILL_1_OAI21X1_1154 ( );
FILL FILL_0_CLKBUF1_86 ( );
FILL FILL_1_CLKBUF1_86 ( );
FILL FILL_2_CLKBUF1_86 ( );
FILL FILL_3_CLKBUF1_86 ( );
FILL FILL_4_CLKBUF1_86 ( );
FILL FILL_0_BUFX4_170 ( );
FILL FILL_1_BUFX4_170 ( );
FILL FILL_2_BUFX4_170 ( );
FILL FILL_0_OAI21X1_1533 ( );
FILL FILL_1_OAI21X1_1533 ( );
FILL FILL_0_BUFX2_27 ( );
FILL FILL_0_OAI21X1_1738 ( );
FILL FILL_1_OAI21X1_1738 ( );
FILL FILL_0_DFFPOSX1_985 ( );
FILL FILL_1_DFFPOSX1_985 ( );
FILL FILL_2_DFFPOSX1_985 ( );
FILL FILL_3_DFFPOSX1_985 ( );
FILL FILL_4_DFFPOSX1_985 ( );
FILL FILL_5_DFFPOSX1_985 ( );
FILL FILL_0_NAND2X1_433 ( );
FILL FILL_0_BUFX2_103 ( );
FILL FILL_0_BUFX2_155 ( );
FILL FILL_0_BUFX2_26 ( );
FILL FILL_1_BUFX2_26 ( );
FILL FILL_0_OAI21X1_283 ( );
FILL FILL_1_OAI21X1_283 ( );
FILL FILL_0_OAI21X1_282 ( );
FILL FILL_1_OAI21X1_282 ( );
FILL FILL_0_BUFX4_203 ( );
FILL FILL_1_BUFX4_203 ( );
FILL FILL_0_CLKBUF1_8 ( );
FILL FILL_1_CLKBUF1_8 ( );
FILL FILL_2_CLKBUF1_8 ( );
FILL FILL_3_CLKBUF1_8 ( );
FILL FILL_4_CLKBUF1_8 ( );
FILL FILL_0_BUFX4_313 ( );
FILL FILL_1_BUFX4_313 ( );
FILL FILL_0_BUFX2_218 ( );
FILL FILL_1_BUFX2_218 ( );
FILL FILL_0_OAI21X1_1823 ( );
FILL FILL_1_OAI21X1_1823 ( );
FILL FILL_2_OAI21X1_1823 ( );
FILL FILL_0_NAND2X1_764 ( );
FILL FILL_0_DFFPOSX1_62 ( );
FILL FILL_1_DFFPOSX1_62 ( );
FILL FILL_2_DFFPOSX1_62 ( );
FILL FILL_3_DFFPOSX1_62 ( );
FILL FILL_4_DFFPOSX1_62 ( );
FILL FILL_5_DFFPOSX1_62 ( );
FILL FILL_0_OAI21X1_1698 ( );
FILL FILL_1_OAI21X1_1698 ( );
FILL FILL_0_OAI21X1_1699 ( );
FILL FILL_1_OAI21X1_1699 ( );
FILL FILL_2_OAI21X1_1699 ( );
FILL FILL_0_BUFX2_821 ( );
FILL FILL_1_BUFX2_821 ( );
FILL FILL_0_BUFX2_715 ( );
FILL FILL_1_BUFX2_715 ( );
FILL FILL_0_DFFPOSX1_187 ( );
FILL FILL_1_DFFPOSX1_187 ( );
FILL FILL_2_DFFPOSX1_187 ( );
FILL FILL_3_DFFPOSX1_187 ( );
FILL FILL_4_DFFPOSX1_187 ( );
FILL FILL_5_DFFPOSX1_187 ( );
FILL FILL_6_DFFPOSX1_187 ( );
FILL FILL_0_DFFPOSX1_1024 ( );
FILL FILL_1_DFFPOSX1_1024 ( );
FILL FILL_2_DFFPOSX1_1024 ( );
FILL FILL_3_DFFPOSX1_1024 ( );
FILL FILL_4_DFFPOSX1_1024 ( );
FILL FILL_5_DFFPOSX1_1024 ( );
FILL FILL_0_OAI21X1_1601 ( );
FILL FILL_1_OAI21X1_1601 ( );
FILL FILL_0_NAND2X1_670 ( );
FILL FILL_1_NAND2X1_670 ( );
FILL FILL_0_BUFX4_193 ( );
FILL FILL_1_BUFX4_193 ( );
FILL FILL_0_BUFX2_662 ( );
FILL FILL_0_BUFX2_857 ( );
FILL FILL_0_BUFX2_726 ( );
FILL FILL_1_BUFX2_726 ( );
FILL FILL_0_NAND2X1_692 ( );
FILL FILL_1_NAND2X1_692 ( );
FILL FILL_0_INVX2_137 ( );
FILL FILL_0_BUFX2_885 ( );
FILL FILL_0_BUFX2_856 ( );
FILL FILL_1_BUFX2_856 ( );
FILL FILL_0_NAND2X1_349 ( );
FILL FILL_0_INVX1_90 ( );
FILL FILL_1_INVX1_90 ( );
FILL FILL_0_BUFX2_269 ( );
FILL FILL_0_OAI21X1_861 ( );
FILL FILL_1_OAI21X1_861 ( );
FILL FILL_2_OAI21X1_861 ( );
FILL FILL_0_INVX1_62 ( );
FILL FILL_0_DFFPOSX1_633 ( );
FILL FILL_1_DFFPOSX1_633 ( );
FILL FILL_2_DFFPOSX1_633 ( );
FILL FILL_3_DFFPOSX1_633 ( );
FILL FILL_4_DFFPOSX1_633 ( );
FILL FILL_5_DFFPOSX1_633 ( );
FILL FILL_6_DFFPOSX1_633 ( );
FILL FILL_0_BUFX2_375 ( );
FILL FILL_1_BUFX2_375 ( );
FILL FILL_0_DFFPOSX1_57 ( );
FILL FILL_1_DFFPOSX1_57 ( );
FILL FILL_2_DFFPOSX1_57 ( );
FILL FILL_3_DFFPOSX1_57 ( );
FILL FILL_4_DFFPOSX1_57 ( );
FILL FILL_5_DFFPOSX1_57 ( );
FILL FILL_6_DFFPOSX1_57 ( );
FILL FILL_0_OAI21X1_1023 ( );
FILL FILL_1_OAI21X1_1023 ( );
FILL FILL_0_OAI21X1_1022 ( );
FILL FILL_1_OAI21X1_1022 ( );
FILL FILL_0_BUFX2_695 ( );
FILL FILL_1_BUFX2_695 ( );
FILL FILL_0_DFFPOSX1_722 ( );
FILL FILL_1_DFFPOSX1_722 ( );
FILL FILL_2_DFFPOSX1_722 ( );
FILL FILL_3_DFFPOSX1_722 ( );
FILL FILL_4_DFFPOSX1_722 ( );
FILL FILL_5_DFFPOSX1_722 ( );
FILL FILL_6_DFFPOSX1_722 ( );
FILL FILL_0_DFFPOSX1_201 ( );
FILL FILL_1_DFFPOSX1_201 ( );
FILL FILL_2_DFFPOSX1_201 ( );
FILL FILL_3_DFFPOSX1_201 ( );
FILL FILL_4_DFFPOSX1_201 ( );
FILL FILL_5_DFFPOSX1_201 ( );
FILL FILL_0_NAND2X1_45 ( );
FILL FILL_0_OAI21X1_45 ( );
FILL FILL_1_OAI21X1_45 ( );
FILL FILL_2_OAI21X1_45 ( );
FILL FILL_0_BUFX2_759 ( );
FILL FILL_1_BUFX2_759 ( );
FILL FILL_0_OAI21X1_1752 ( );
FILL FILL_1_OAI21X1_1752 ( );
FILL FILL_0_OAI21X1_27 ( );
FILL FILL_1_OAI21X1_27 ( );
FILL FILL_0_BUFX4_136 ( );
FILL FILL_1_BUFX4_136 ( );
FILL FILL_0_OAI21X1_309 ( );
FILL FILL_1_OAI21X1_309 ( );
FILL FILL_0_OAI21X1_308 ( );
FILL FILL_1_OAI21X1_308 ( );
FILL FILL_0_DFFPOSX1_942 ( );
FILL FILL_1_DFFPOSX1_942 ( );
FILL FILL_2_DFFPOSX1_942 ( );
FILL FILL_3_DFFPOSX1_942 ( );
FILL FILL_4_DFFPOSX1_942 ( );
FILL FILL_5_DFFPOSX1_942 ( );
FILL FILL_0_BUFX2_46 ( );
FILL FILL_0_CLKBUF1_98 ( );
FILL FILL_1_CLKBUF1_98 ( );
FILL FILL_2_CLKBUF1_98 ( );
FILL FILL_3_CLKBUF1_98 ( );
FILL FILL_4_CLKBUF1_98 ( );
FILL FILL_0_BUFX2_57 ( );
FILL FILL_1_BUFX2_57 ( );
FILL FILL_0_OAI21X1_1613 ( );
FILL FILL_1_OAI21X1_1613 ( );
FILL FILL_2_OAI21X1_1613 ( );
FILL FILL_0_OAI21X1_1399 ( );
FILL FILL_1_OAI21X1_1399 ( );
FILL FILL_2_OAI21X1_1399 ( );
FILL FILL_0_NAND2X1_407 ( );
FILL FILL_1_NAND2X1_407 ( );
FILL FILL_0_OAI21X1_1041 ( );
FILL FILL_1_OAI21X1_1041 ( );
FILL FILL_0_OAI21X1_1221 ( );
FILL FILL_1_OAI21X1_1221 ( );
FILL FILL_0_NAND2X1_590 ( );
FILL FILL_1_NAND2X1_590 ( );
FILL FILL_0_OAI21X1_1104 ( );
FILL FILL_1_OAI21X1_1104 ( );
FILL FILL_0_OAI21X1_1218 ( );
FILL FILL_1_OAI21X1_1218 ( );
FILL FILL_2_OAI21X1_1218 ( );
FILL FILL_0_NAND2X1_472 ( );
FILL FILL_1_NAND2X1_472 ( );
FILL FILL_0_INVX2_58 ( );
FILL FILL_0_OAI21X1_1396 ( );
FILL FILL_1_OAI21X1_1396 ( );
FILL FILL_0_OAI21X1_1397 ( );
FILL FILL_1_OAI21X1_1397 ( );
FILL FILL_0_INVX2_59 ( );
FILL FILL_0_OAI21X1_1109 ( );
FILL FILL_1_OAI21X1_1109 ( );
FILL FILL_2_OAI21X1_1109 ( );
FILL FILL_0_INVX1_184 ( );
FILL FILL_0_DFFPOSX1_753 ( );
FILL FILL_1_DFFPOSX1_753 ( );
FILL FILL_2_DFFPOSX1_753 ( );
FILL FILL_3_DFFPOSX1_753 ( );
FILL FILL_4_DFFPOSX1_753 ( );
FILL FILL_5_DFFPOSX1_753 ( );
FILL FILL_0_NOR2X1_127 ( );
FILL FILL_1_NOR2X1_127 ( );
FILL FILL_0_OAI21X1_1117 ( );
FILL FILL_1_OAI21X1_1117 ( );
FILL FILL_0_NOR2X1_179 ( );
FILL FILL_1_NOR2X1_179 ( );
FILL FILL_0_NAND2X1_481 ( );
FILL FILL_0_XNOR2X1_75 ( );
FILL FILL_1_XNOR2X1_75 ( );
FILL FILL_2_XNOR2X1_75 ( );
FILL FILL_3_XNOR2X1_75 ( );
FILL FILL_0_OAI21X1_641 ( );
FILL FILL_1_OAI21X1_641 ( );
FILL FILL_0_DFFPOSX1_946 ( );
FILL FILL_1_DFFPOSX1_946 ( );
FILL FILL_2_DFFPOSX1_946 ( );
FILL FILL_3_DFFPOSX1_946 ( );
FILL FILL_4_DFFPOSX1_946 ( );
FILL FILL_5_DFFPOSX1_946 ( );
FILL FILL_0_OAI21X1_1415 ( );
FILL FILL_1_OAI21X1_1415 ( );
FILL FILL_0_OAI21X1_1046 ( );
FILL FILL_1_OAI21X1_1046 ( );
FILL FILL_0_BUFX2_982 ( );
FILL FILL_0_BUFX4_231 ( );
FILL FILL_1_BUFX4_231 ( );
FILL FILL_0_OAI21X1_490 ( );
FILL FILL_1_OAI21X1_490 ( );
FILL FILL_2_OAI21X1_490 ( );
FILL FILL_0_DFFPOSX1_819 ( );
FILL FILL_1_DFFPOSX1_819 ( );
FILL FILL_2_DFFPOSX1_819 ( );
FILL FILL_3_DFFPOSX1_819 ( );
FILL FILL_4_DFFPOSX1_819 ( );
FILL FILL_5_DFFPOSX1_819 ( );
FILL FILL_6_DFFPOSX1_819 ( );
FILL FILL_0_NAND2X1_484 ( );
FILL FILL_0_XNOR2X1_56 ( );
FILL FILL_1_XNOR2X1_56 ( );
FILL FILL_2_XNOR2X1_56 ( );
FILL FILL_3_XNOR2X1_56 ( );
FILL FILL_0_AND2X2_16 ( );
FILL FILL_1_AND2X2_16 ( );
FILL FILL_0_NAND2X1_305 ( );
FILL FILL_1_NAND2X1_305 ( );
FILL FILL_0_NAND2X1_487 ( );
FILL FILL_0_DFFPOSX1_544 ( );
FILL FILL_1_DFFPOSX1_544 ( );
FILL FILL_2_DFFPOSX1_544 ( );
FILL FILL_3_DFFPOSX1_544 ( );
FILL FILL_4_DFFPOSX1_544 ( );
FILL FILL_5_DFFPOSX1_544 ( );
FILL FILL_6_DFFPOSX1_544 ( );
FILL FILL_0_NAND2X1_307 ( );
FILL FILL_1_NAND2X1_307 ( );
FILL FILL_0_AND2X2_17 ( );
FILL FILL_1_AND2X2_17 ( );
FILL FILL_0_OAI21X1_275 ( );
FILL FILL_1_OAI21X1_275 ( );
FILL FILL_0_DFFPOSX1_329 ( );
FILL FILL_1_DFFPOSX1_329 ( );
FILL FILL_2_DFFPOSX1_329 ( );
FILL FILL_3_DFFPOSX1_329 ( );
FILL FILL_4_DFFPOSX1_329 ( );
FILL FILL_5_DFFPOSX1_329 ( );
FILL FILL_0_NAND3X1_63 ( );
FILL FILL_1_NAND3X1_63 ( );
FILL FILL_0_NAND2X1_594 ( );
FILL FILL_0_INVX2_96 ( );
FILL FILL_0_NAND3X1_39 ( );
FILL FILL_1_NAND3X1_39 ( );
FILL FILL_0_OAI21X1_1242 ( );
FILL FILL_1_OAI21X1_1242 ( );
FILL FILL_0_OAI21X1_1243 ( );
FILL FILL_1_OAI21X1_1243 ( );
FILL FILL_0_NOR2X1_183 ( );
FILL FILL_0_BUFX4_210 ( );
FILL FILL_1_BUFX4_210 ( );
FILL FILL_0_INVX2_66 ( );
FILL FILL_0_NAND2X1_595 ( );
FILL FILL_1_NAND2X1_595 ( );
FILL FILL_0_INVX4_34 ( );
FILL FILL_0_NOR2X1_182 ( );
FILL FILL_1_NOR2X1_182 ( );
FILL FILL_0_DFFPOSX1_890 ( );
FILL FILL_1_DFFPOSX1_890 ( );
FILL FILL_2_DFFPOSX1_890 ( );
FILL FILL_3_DFFPOSX1_890 ( );
FILL FILL_4_DFFPOSX1_890 ( );
FILL FILL_5_DFFPOSX1_890 ( );
FILL FILL_0_INVX1_200 ( );
FILL FILL_0_OAI21X1_1252 ( );
FILL FILL_1_OAI21X1_1252 ( );
FILL FILL_0_INVX2_105 ( );
FILL FILL_0_OAI21X1_1430 ( );
FILL FILL_1_OAI21X1_1430 ( );
FILL FILL_0_OAI21X1_1253 ( );
FILL FILL_1_OAI21X1_1253 ( );
FILL FILL_0_DFFPOSX1_952 ( );
FILL FILL_1_DFFPOSX1_952 ( );
FILL FILL_2_DFFPOSX1_952 ( );
FILL FILL_3_DFFPOSX1_952 ( );
FILL FILL_4_DFFPOSX1_952 ( );
FILL FILL_5_DFFPOSX1_952 ( );
FILL FILL_6_DFFPOSX1_952 ( );
FILL FILL_0_BUFX4_44 ( );
FILL FILL_1_BUFX4_44 ( );
FILL FILL_0_OAI21X1_1255 ( );
FILL FILL_1_OAI21X1_1255 ( );
FILL FILL_0_DFFPOSX1_888 ( );
FILL FILL_1_DFFPOSX1_888 ( );
FILL FILL_2_DFFPOSX1_888 ( );
FILL FILL_3_DFFPOSX1_888 ( );
FILL FILL_4_DFFPOSX1_888 ( );
FILL FILL_5_DFFPOSX1_888 ( );
FILL FILL_0_OAI21X1_1254 ( );
FILL FILL_1_OAI21X1_1254 ( );
FILL FILL_2_OAI21X1_1254 ( );
FILL FILL_0_BUFX4_65 ( );
FILL FILL_1_BUFX4_65 ( );
FILL FILL_0_OAI21X1_1694 ( );
FILL FILL_1_OAI21X1_1694 ( );
FILL FILL_0_DFFPOSX1_939 ( );
FILL FILL_1_DFFPOSX1_939 ( );
FILL FILL_2_DFFPOSX1_939 ( );
FILL FILL_3_DFFPOSX1_939 ( );
FILL FILL_4_DFFPOSX1_939 ( );
FILL FILL_5_DFFPOSX1_939 ( );
FILL FILL_6_DFFPOSX1_939 ( );
FILL FILL_0_OAI21X1_1390 ( );
FILL FILL_1_OAI21X1_1390 ( );
FILL FILL_0_BUFX4_97 ( );
FILL FILL_1_BUFX4_97 ( );
FILL FILL_0_DFFPOSX1_26 ( );
FILL FILL_1_DFFPOSX1_26 ( );
FILL FILL_2_DFFPOSX1_26 ( );
FILL FILL_3_DFFPOSX1_26 ( );
FILL FILL_4_DFFPOSX1_26 ( );
FILL FILL_5_DFFPOSX1_26 ( );
FILL FILL_6_DFFPOSX1_26 ( );
FILL FILL_0_OAI21X1_1755 ( );
FILL FILL_1_OAI21X1_1755 ( );
FILL FILL_2_OAI21X1_1755 ( );
FILL FILL_0_OAI21X1_1754 ( );
FILL FILL_1_OAI21X1_1754 ( );
FILL FILL_0_BUFX2_83 ( );
FILL FILL_1_BUFX2_83 ( );
FILL FILL_0_DFFPOSX1_835 ( );
FILL FILL_1_DFFPOSX1_835 ( );
FILL FILL_2_DFFPOSX1_835 ( );
FILL FILL_3_DFFPOSX1_835 ( );
FILL FILL_4_DFFPOSX1_835 ( );
FILL FILL_5_DFFPOSX1_835 ( );
FILL FILL_6_DFFPOSX1_835 ( );
FILL FILL_0_BUFX4_229 ( );
FILL FILL_1_BUFX4_229 ( );
FILL FILL_0_XNOR2X1_64 ( );
FILL FILL_1_XNOR2X1_64 ( );
FILL FILL_2_XNOR2X1_64 ( );
FILL FILL_3_XNOR2X1_64 ( );
FILL FILL_0_OAI21X1_1147 ( );
FILL FILL_1_OAI21X1_1147 ( );
FILL FILL_0_BUFX4_377 ( );
FILL FILL_1_BUFX4_377 ( );
FILL FILL_0_OAI21X1_1652 ( );
FILL FILL_1_OAI21X1_1652 ( );
FILL FILL_0_OAI21X1_273 ( );
FILL FILL_1_OAI21X1_273 ( );
FILL FILL_0_DFFPOSX1_340 ( );
FILL FILL_1_DFFPOSX1_340 ( );
FILL FILL_2_DFFPOSX1_340 ( );
FILL FILL_3_DFFPOSX1_340 ( );
FILL FILL_4_DFFPOSX1_340 ( );
FILL FILL_5_DFFPOSX1_340 ( );
FILL FILL_0_BUFX2_22 ( );
FILL FILL_0_OAI21X1_297 ( );
FILL FILL_1_OAI21X1_297 ( );
FILL FILL_0_DFFPOSX1_239 ( );
FILL FILL_1_DFFPOSX1_239 ( );
FILL FILL_2_DFFPOSX1_239 ( );
FILL FILL_3_DFFPOSX1_239 ( );
FILL FILL_4_DFFPOSX1_239 ( );
FILL FILL_5_DFFPOSX1_239 ( );
FILL FILL_6_DFFPOSX1_239 ( );
FILL FILL_0_NAND2X1_431 ( );
FILL FILL_0_BUFX2_23 ( );
FILL FILL_1_BUFX2_23 ( );
FILL FILL_0_DFFPOSX1_303 ( );
FILL FILL_1_DFFPOSX1_303 ( );
FILL FILL_2_DFFPOSX1_303 ( );
FILL FILL_3_DFFPOSX1_303 ( );
FILL FILL_4_DFFPOSX1_303 ( );
FILL FILL_5_DFFPOSX1_303 ( );
FILL FILL_0_BUFX4_202 ( );
FILL FILL_1_BUFX4_202 ( );
FILL FILL_2_BUFX4_202 ( );
FILL FILL_0_DFFPOSX1_53 ( );
FILL FILL_1_DFFPOSX1_53 ( );
FILL FILL_2_DFFPOSX1_53 ( );
FILL FILL_3_DFFPOSX1_53 ( );
FILL FILL_4_DFFPOSX1_53 ( );
FILL FILL_5_DFFPOSX1_53 ( );
FILL FILL_0_DFFPOSX1_841 ( );
FILL FILL_1_DFFPOSX1_841 ( );
FILL FILL_2_DFFPOSX1_841 ( );
FILL FILL_3_DFFPOSX1_841 ( );
FILL FILL_4_DFFPOSX1_841 ( );
FILL FILL_5_DFFPOSX1_841 ( );
FILL FILL_6_DFFPOSX1_841 ( );
FILL FILL_0_OAI21X1_1745 ( );
FILL FILL_1_OAI21X1_1745 ( );
FILL FILL_0_DFFPOSX1_118 ( );
FILL FILL_1_DFFPOSX1_118 ( );
FILL FILL_2_DFFPOSX1_118 ( );
FILL FILL_3_DFFPOSX1_118 ( );
FILL FILL_4_DFFPOSX1_118 ( );
FILL FILL_5_DFFPOSX1_118 ( );
FILL FILL_0_NAND2X1_532 ( );
FILL FILL_1_NAND2X1_532 ( );
FILL FILL_0_BUFX2_232 ( );
FILL FILL_1_BUFX2_232 ( );
FILL FILL_0_DFFPOSX1_840 ( );
FILL FILL_1_DFFPOSX1_840 ( );
FILL FILL_2_DFFPOSX1_840 ( );
FILL FILL_3_DFFPOSX1_840 ( );
FILL FILL_4_DFFPOSX1_840 ( );
FILL FILL_5_DFFPOSX1_840 ( );
FILL FILL_0_DFFPOSX1_51 ( );
FILL FILL_1_DFFPOSX1_51 ( );
FILL FILL_2_DFFPOSX1_51 ( );
FILL FILL_3_DFFPOSX1_51 ( );
FILL FILL_4_DFFPOSX1_51 ( );
FILL FILL_5_DFFPOSX1_51 ( );
FILL FILL_0_DFFPOSX1_82 ( );
FILL FILL_1_DFFPOSX1_82 ( );
FILL FILL_2_DFFPOSX1_82 ( );
FILL FILL_3_DFFPOSX1_82 ( );
FILL FILL_4_DFFPOSX1_82 ( );
FILL FILL_5_DFFPOSX1_82 ( );
FILL FILL_0_OAI21X1_1532 ( );
FILL FILL_1_OAI21X1_1532 ( );
FILL FILL_0_BUFX2_28 ( );
FILL FILL_1_BUFX2_28 ( );
FILL FILL_0_OAI21X1_1739 ( );
FILL FILL_1_OAI21X1_1739 ( );
FILL FILL_0_BUFX2_219 ( );
FILL FILL_1_BUFX2_219 ( );
FILL FILL_0_BUFX2_751 ( );
FILL FILL_1_BUFX2_751 ( );
FILL FILL_0_BUFX2_108 ( );
FILL FILL_0_DFFPOSX1_18 ( );
FILL FILL_1_DFFPOSX1_18 ( );
FILL FILL_2_DFFPOSX1_18 ( );
FILL FILL_3_DFFPOSX1_18 ( );
FILL FILL_4_DFFPOSX1_18 ( );
FILL FILL_5_DFFPOSX1_18 ( );
FILL FILL_6_DFFPOSX1_18 ( );
FILL FILL_0_DFFPOSX1_341 ( );
FILL FILL_1_DFFPOSX1_341 ( );
FILL FILL_2_DFFPOSX1_341 ( );
FILL FILL_3_DFFPOSX1_341 ( );
FILL FILL_4_DFFPOSX1_341 ( );
FILL FILL_5_DFFPOSX1_341 ( );
FILL FILL_6_DFFPOSX1_341 ( );
FILL FILL_0_OAI21X1_1595 ( );
FILL FILL_1_OAI21X1_1595 ( );
FILL FILL_0_DFFPOSX1_143 ( );
FILL FILL_1_DFFPOSX1_143 ( );
FILL FILL_2_DFFPOSX1_143 ( );
FILL FILL_3_DFFPOSX1_143 ( );
FILL FILL_4_DFFPOSX1_143 ( );
FILL FILL_5_DFFPOSX1_143 ( );
FILL FILL_6_DFFPOSX1_143 ( );
FILL FILL_0_OAI21X1_299 ( );
FILL FILL_1_OAI21X1_299 ( );
FILL FILL_0_DFFPOSX1_1012 ( );
FILL FILL_1_DFFPOSX1_1012 ( );
FILL FILL_2_DFFPOSX1_1012 ( );
FILL FILL_3_DFFPOSX1_1012 ( );
FILL FILL_4_DFFPOSX1_1012 ( );
FILL FILL_5_DFFPOSX1_1012 ( );
FILL FILL_6_DFFPOSX1_1012 ( );
FILL FILL_0_OAI21X1_1589 ( );
FILL FILL_1_OAI21X1_1589 ( );
FILL FILL_0_NAND2X1_658 ( );
FILL FILL_1_NAND2X1_658 ( );
FILL FILL_0_OAI21X1_1662 ( );
FILL FILL_1_OAI21X1_1662 ( );
FILL FILL_0_OAI21X1_1663 ( );
FILL FILL_1_OAI21X1_1663 ( );
FILL FILL_0_DFFPOSX1_44 ( );
FILL FILL_1_DFFPOSX1_44 ( );
FILL FILL_2_DFFPOSX1_44 ( );
FILL FILL_3_DFFPOSX1_44 ( );
FILL FILL_4_DFFPOSX1_44 ( );
FILL FILL_5_DFFPOSX1_44 ( );
FILL FILL_6_DFFPOSX1_44 ( );
FILL FILL_0_INVX2_164 ( );
FILL FILL_0_DFFPOSX1_207 ( );
FILL FILL_1_DFFPOSX1_207 ( );
FILL FILL_2_DFFPOSX1_207 ( );
FILL FILL_3_DFFPOSX1_207 ( );
FILL FILL_4_DFFPOSX1_207 ( );
FILL FILL_5_DFFPOSX1_207 ( );
FILL FILL_0_OAI21X1_51 ( );
FILL FILL_1_OAI21X1_51 ( );
FILL FILL_0_OAI21X1_1622 ( );
FILL FILL_1_OAI21X1_1622 ( );
FILL FILL_0_NAND2X1_690 ( );
FILL FILL_1_NAND2X1_690 ( );
FILL FILL_0_DFFPOSX1_12 ( );
FILL FILL_1_DFFPOSX1_12 ( );
FILL FILL_2_DFFPOSX1_12 ( );
FILL FILL_3_DFFPOSX1_12 ( );
FILL FILL_4_DFFPOSX1_12 ( );
FILL FILL_5_DFFPOSX1_12 ( );
FILL FILL_0_DFFPOSX1_660 ( );
FILL FILL_1_DFFPOSX1_660 ( );
FILL FILL_2_DFFPOSX1_660 ( );
FILL FILL_3_DFFPOSX1_660 ( );
FILL FILL_4_DFFPOSX1_660 ( );
FILL FILL_5_DFFPOSX1_660 ( );
FILL FILL_0_NAND2X1_355 ( );
FILL FILL_0_DFFPOSX1_624 ( );
FILL FILL_1_DFFPOSX1_624 ( );
FILL FILL_2_DFFPOSX1_624 ( );
FILL FILL_3_DFFPOSX1_624 ( );
FILL FILL_4_DFFPOSX1_624 ( );
FILL FILL_5_DFFPOSX1_624 ( );
FILL FILL_6_DFFPOSX1_624 ( );
FILL FILL_0_OAI21X1_852 ( );
FILL FILL_1_OAI21X1_852 ( );
FILL FILL_0_INVX1_53 ( );
FILL FILL_0_BUFX2_359 ( );
FILL FILL_1_BUFX2_359 ( );
FILL FILL_0_DFFPOSX1_736 ( );
FILL FILL_1_DFFPOSX1_736 ( );
FILL FILL_2_DFFPOSX1_736 ( );
FILL FILL_3_DFFPOSX1_736 ( );
FILL FILL_4_DFFPOSX1_736 ( );
FILL FILL_5_DFFPOSX1_736 ( );
FILL FILL_0_OAI21X1_1021 ( );
FILL FILL_1_OAI21X1_1021 ( );
FILL FILL_0_OAI21X1_1020 ( );
FILL FILL_1_OAI21X1_1020 ( );
FILL FILL_0_OAI21X1_993 ( );
FILL FILL_1_OAI21X1_993 ( );
FILL FILL_0_OAI21X1_992 ( );
FILL FILL_1_OAI21X1_992 ( );
FILL FILL_0_OAI21X1_990 ( );
FILL FILL_1_OAI21X1_990 ( );
FILL FILL_2_OAI21X1_990 ( );
FILL FILL_0_OAI21X1_991 ( );
FILL FILL_1_OAI21X1_991 ( );
FILL FILL_0_BUFX2_872 ( );
FILL FILL_0_DFFPOSX1_721 ( );
FILL FILL_1_DFFPOSX1_721 ( );
FILL FILL_2_DFFPOSX1_721 ( );
FILL FILL_3_DFFPOSX1_721 ( );
FILL FILL_4_DFFPOSX1_721 ( );
FILL FILL_5_DFFPOSX1_721 ( );
FILL FILL_0_OAI21X1_266 ( );
FILL FILL_1_OAI21X1_266 ( );
FILL FILL_2_OAI21X1_266 ( );
FILL FILL_0_NAND2X1_27 ( );
FILL FILL_1_NAND2X1_27 ( );
FILL FILL_0_DFFPOSX1_183 ( );
FILL FILL_1_DFFPOSX1_183 ( );
FILL FILL_2_DFFPOSX1_183 ( );
FILL FILL_3_DFFPOSX1_183 ( );
FILL FILL_4_DFFPOSX1_183 ( );
FILL FILL_5_DFFPOSX1_183 ( );
FILL FILL_0_BUFX2_1019 ( );
FILL FILL_1_BUFX2_1019 ( );
FILL FILL_0_DFFPOSX1_346 ( );
FILL FILL_1_DFFPOSX1_346 ( );
FILL FILL_2_DFFPOSX1_346 ( );
FILL FILL_3_DFFPOSX1_346 ( );
FILL FILL_4_DFFPOSX1_346 ( );
FILL FILL_5_DFFPOSX1_346 ( );
FILL FILL_0_CLKBUF1_96 ( );
FILL FILL_1_CLKBUF1_96 ( );
FILL FILL_2_CLKBUF1_96 ( );
FILL FILL_3_CLKBUF1_96 ( );
FILL FILL_4_CLKBUF1_96 ( );
FILL FILL_0_DFFPOSX1_52 ( );
FILL FILL_1_DFFPOSX1_52 ( );
FILL FILL_2_DFFPOSX1_52 ( );
FILL FILL_3_DFFPOSX1_52 ( );
FILL FILL_4_DFFPOSX1_52 ( );
FILL FILL_5_DFFPOSX1_52 ( );
FILL FILL_6_DFFPOSX1_52 ( );
FILL FILL_0_BUFX2_567 ( );
FILL FILL_1_BUFX2_567 ( );
FILL FILL_0_BUFX4_100 ( );
FILL FILL_1_BUFX4_100 ( );
FILL FILL_0_OAI21X1_1219 ( );
FILL FILL_1_OAI21X1_1219 ( );
FILL FILL_0_DFFPOSX1_877 ( );
FILL FILL_1_DFFPOSX1_877 ( );
FILL FILL_2_DFFPOSX1_877 ( );
FILL FILL_3_DFFPOSX1_877 ( );
FILL FILL_4_DFFPOSX1_877 ( );
FILL FILL_5_DFFPOSX1_877 ( );
FILL FILL_0_OAI21X1_1220 ( );
FILL FILL_1_OAI21X1_1220 ( );
FILL FILL_0_NAND2X1_470 ( );
FILL FILL_1_NAND2X1_470 ( );
FILL FILL_0_INVX2_56 ( );
FILL FILL_0_NOR2X1_177 ( );
FILL FILL_0_INVX1_183 ( );
FILL FILL_0_AOI21X1_36 ( );
FILL FILL_1_AOI21X1_36 ( );
FILL FILL_0_INVX4_32 ( );
FILL FILL_0_NAND2X1_477 ( );
FILL FILL_1_NAND2X1_477 ( );
FILL FILL_0_OAI21X1_1108 ( );
FILL FILL_1_OAI21X1_1108 ( );
FILL FILL_2_OAI21X1_1108 ( );
FILL FILL_0_OAI21X1_1107 ( );
FILL FILL_1_OAI21X1_1107 ( );
FILL FILL_0_NAND2X1_411 ( );
FILL FILL_1_NAND2X1_411 ( );
FILL FILL_0_OAI21X1_1045 ( );
FILL FILL_1_OAI21X1_1045 ( );
FILL FILL_0_OAI21X1_230 ( );
FILL FILL_1_OAI21X1_230 ( );
FILL FILL_0_NAND2X1_482 ( );
FILL FILL_1_NAND2X1_482 ( );
FILL FILL_0_NOR2X1_121 ( );
FILL FILL_1_NOR2X1_121 ( );
FILL FILL_0_INVX2_62 ( );
FILL FILL_0_OAI21X1_1234 ( );
FILL FILL_1_OAI21X1_1234 ( );
FILL FILL_0_OAI21X1_1235 ( );
FILL FILL_1_OAI21X1_1235 ( );
FILL FILL_0_DFFPOSX1_882 ( );
FILL FILL_1_DFFPOSX1_882 ( );
FILL FILL_2_DFFPOSX1_882 ( );
FILL FILL_3_DFFPOSX1_882 ( );
FILL FILL_4_DFFPOSX1_882 ( );
FILL FILL_5_DFFPOSX1_882 ( );
FILL FILL_6_DFFPOSX1_882 ( );
FILL FILL_0_BUFX4_251 ( );
FILL FILL_1_BUFX4_251 ( );
FILL FILL_0_OAI21X1_1414 ( );
FILL FILL_1_OAI21X1_1414 ( );
FILL FILL_0_NAND2X1_412 ( );
FILL FILL_1_NAND2X1_412 ( );
FILL FILL_0_DFFPOSX1_754 ( );
FILL FILL_1_DFFPOSX1_754 ( );
FILL FILL_2_DFFPOSX1_754 ( );
FILL FILL_3_DFFPOSX1_754 ( );
FILL FILL_4_DFFPOSX1_754 ( );
FILL FILL_5_DFFPOSX1_754 ( );
FILL FILL_6_DFFPOSX1_754 ( );
FILL FILL_0_NAND2X1_256 ( );
FILL FILL_0_DFFPOSX1_478 ( );
FILL FILL_1_DFFPOSX1_478 ( );
FILL FILL_2_DFFPOSX1_478 ( );
FILL FILL_3_DFFPOSX1_478 ( );
FILL FILL_4_DFFPOSX1_478 ( );
FILL FILL_5_DFFPOSX1_478 ( );
FILL FILL_0_BUFX2_1032 ( );
FILL FILL_1_BUFX2_1032 ( );
FILL FILL_0_OAI21X1_1122 ( );
FILL FILL_1_OAI21X1_1122 ( );
FILL FILL_0_NAND2X1_485 ( );
FILL FILL_1_NAND2X1_485 ( );
FILL FILL_0_NAND2X1_486 ( );
FILL FILL_1_NAND2X1_486 ( );
FILL FILL_0_OAI21X1_1124 ( );
FILL FILL_1_OAI21X1_1124 ( );
FILL FILL_0_NAND2X1_488 ( );
FILL FILL_1_NAND2X1_488 ( );
FILL FILL_0_INVX2_95 ( );
FILL FILL_0_AOI21X1_25 ( );
FILL FILL_1_AOI21X1_25 ( );
FILL FILL_0_OAI21X1_651 ( );
FILL FILL_1_OAI21X1_651 ( );
FILL FILL_0_OAI21X1_650 ( );
FILL FILL_1_OAI21X1_650 ( );
FILL FILL_2_OAI21X1_650 ( );
FILL FILL_0_BUFX4_3 ( );
FILL FILL_1_BUFX4_3 ( );
FILL FILL_0_OAI21X1_146 ( );
FILL FILL_1_OAI21X1_146 ( );
FILL FILL_0_OAI21X1_147 ( );
FILL FILL_1_OAI21X1_147 ( );
FILL FILL_0_DFFPOSX1_265 ( );
FILL FILL_1_DFFPOSX1_265 ( );
FILL FILL_2_DFFPOSX1_265 ( );
FILL FILL_3_DFFPOSX1_265 ( );
FILL FILL_4_DFFPOSX1_265 ( );
FILL FILL_5_DFFPOSX1_265 ( );
FILL FILL_6_DFFPOSX1_265 ( );
FILL FILL_0_INVX2_65 ( );
FILL FILL_0_NOR2X1_129 ( );
FILL FILL_1_NOR2X1_129 ( );
FILL FILL_0_NAND2X1_489 ( );
FILL FILL_1_NAND2X1_489 ( );
FILL FILL_0_OAI21X1_1127 ( );
FILL FILL_1_OAI21X1_1127 ( );
FILL FILL_0_NAND2X1_492 ( );
FILL FILL_1_NAND2X1_492 ( );
FILL FILL_0_OAI21X1_1049 ( );
FILL FILL_1_OAI21X1_1049 ( );
FILL FILL_0_DFFPOSX1_757 ( );
FILL FILL_1_DFFPOSX1_757 ( );
FILL FILL_2_DFFPOSX1_757 ( );
FILL FILL_3_DFFPOSX1_757 ( );
FILL FILL_4_DFFPOSX1_757 ( );
FILL FILL_5_DFFPOSX1_757 ( );
FILL FILL_6_DFFPOSX1_757 ( );
FILL FILL_0_OAI21X1_1050 ( );
FILL FILL_1_OAI21X1_1050 ( );
FILL FILL_0_OAI21X1_1259 ( );
FILL FILL_1_OAI21X1_1259 ( );
FILL FILL_0_NOR2X1_181 ( );
FILL FILL_1_NOR2X1_181 ( );
FILL FILL_0_BUFX4_340 ( );
FILL FILL_1_BUFX4_340 ( );
FILL FILL_0_OAI21X1_1260 ( );
FILL FILL_1_OAI21X1_1260 ( );
FILL FILL_2_OAI21X1_1260 ( );
FILL FILL_0_OAI21X1_1261 ( );
FILL FILL_1_OAI21X1_1261 ( );
FILL FILL_0_AOI21X1_46 ( );
FILL FILL_1_AOI21X1_46 ( );
FILL FILL_0_INVX2_68 ( );
FILL FILL_0_NOR2X1_184 ( );
FILL FILL_0_OAI21X1_1256 ( );
FILL FILL_1_OAI21X1_1256 ( );
FILL FILL_0_OAI21X1_1431 ( );
FILL FILL_1_OAI21X1_1431 ( );
FILL FILL_0_OAI21X1_1433 ( );
FILL FILL_1_OAI21X1_1433 ( );
FILL FILL_0_OAI21X1_1432 ( );
FILL FILL_1_OAI21X1_1432 ( );
FILL FILL_2_OAI21X1_1432 ( );
FILL FILL_0_BUFX2_605 ( );
FILL FILL_0_OAI21X1_73 ( );
FILL FILL_1_OAI21X1_73 ( );
FILL FILL_0_OAI21X1_72 ( );
FILL FILL_1_OAI21X1_72 ( );
FILL FILL_0_DFFPOSX1_228 ( );
FILL FILL_1_DFFPOSX1_228 ( );
FILL FILL_2_DFFPOSX1_228 ( );
FILL FILL_3_DFFPOSX1_228 ( );
FILL FILL_4_DFFPOSX1_228 ( );
FILL FILL_5_DFFPOSX1_228 ( );
FILL FILL_6_DFFPOSX1_228 ( );
FILL FILL_0_OAI21X1_1765 ( );
FILL FILL_1_OAI21X1_1765 ( );
FILL FILL_0_DFFPOSX1_95 ( );
FILL FILL_1_DFFPOSX1_95 ( );
FILL FILL_2_DFFPOSX1_95 ( );
FILL FILL_3_DFFPOSX1_95 ( );
FILL FILL_4_DFFPOSX1_95 ( );
FILL FILL_5_DFFPOSX1_95 ( );
FILL FILL_0_NAND2X1_24 ( );
FILL FILL_0_OAI21X1_24 ( );
FILL FILL_1_OAI21X1_24 ( );
FILL FILL_0_OAI21X1_1608 ( );
FILL FILL_1_OAI21X1_1608 ( );
FILL FILL_0_OAI21X1_1636 ( );
FILL FILL_1_OAI21X1_1636 ( );
FILL FILL_0_NAND2X1_704 ( );
FILL FILL_1_NAND2X1_704 ( );
FILL FILL_0_BUFX2_730 ( );
FILL FILL_1_BUFX2_730 ( );
FILL FILL_0_BUFX2_733 ( );
FILL FILL_1_BUFX2_733 ( );
FILL FILL_0_NAND2X1_44 ( );
FILL FILL_1_NAND2X1_44 ( );
FILL FILL_0_DFFPOSX1_200 ( );
FILL FILL_1_DFFPOSX1_200 ( );
FILL FILL_2_DFFPOSX1_200 ( );
FILL FILL_3_DFFPOSX1_200 ( );
FILL FILL_4_DFFPOSX1_200 ( );
FILL FILL_5_DFFPOSX1_200 ( );
FILL FILL_6_DFFPOSX1_200 ( );
FILL FILL_0_OAI21X1_44 ( );
FILL FILL_1_OAI21X1_44 ( );
FILL FILL_0_DFFPOSX1_339 ( );
FILL FILL_1_DFFPOSX1_339 ( );
FILL FILL_2_DFFPOSX1_339 ( );
FILL FILL_3_DFFPOSX1_339 ( );
FILL FILL_4_DFFPOSX1_339 ( );
FILL FILL_5_DFFPOSX1_339 ( );
FILL FILL_0_NAND2X1_522 ( );
FILL FILL_1_NAND2X1_522 ( );
FILL FILL_0_OAI21X1_288 ( );
FILL FILL_1_OAI21X1_288 ( );
FILL FILL_0_DFFPOSX1_328 ( );
FILL FILL_1_DFFPOSX1_328 ( );
FILL FILL_2_DFFPOSX1_328 ( );
FILL FILL_3_DFFPOSX1_328 ( );
FILL FILL_4_DFFPOSX1_328 ( );
FILL FILL_5_DFFPOSX1_328 ( );
FILL FILL_6_DFFPOSX1_328 ( );
FILL FILL_0_OAI21X1_272 ( );
FILL FILL_1_OAI21X1_272 ( );
FILL FILL_2_OAI21X1_272 ( );
FILL FILL_0_BUFX2_807 ( );
FILL FILL_0_BUFX2_148 ( );
FILL FILL_1_BUFX2_148 ( );
FILL FILL_0_BUFX2_84 ( );
FILL FILL_1_BUFX2_84 ( );
FILL FILL_0_DFFPOSX1_148 ( );
FILL FILL_1_DFFPOSX1_148 ( );
FILL FILL_2_DFFPOSX1_148 ( );
FILL FILL_3_DFFPOSX1_148 ( );
FILL FILL_4_DFFPOSX1_148 ( );
FILL FILL_5_DFFPOSX1_148 ( );
FILL FILL_6_DFFPOSX1_148 ( );
FILL FILL_0_OAI21X1_169 ( );
FILL FILL_1_OAI21X1_169 ( );
FILL FILL_0_OAI21X1_168 ( );
FILL FILL_1_OAI21X1_168 ( );
FILL FILL_2_OAI21X1_168 ( );
FILL FILL_0_BUFX4_148 ( );
FILL FILL_1_BUFX4_148 ( );
FILL FILL_0_BUFX2_1012 ( );
FILL FILL_1_BUFX2_1012 ( );
FILL FILL_0_BUFX2_672 ( );
FILL FILL_0_OAI21X1_1143 ( );
FILL FILL_1_OAI21X1_1143 ( );
FILL FILL_0_OAI21X1_222 ( );
FILL FILL_1_OAI21X1_222 ( );
FILL FILL_0_OAI21X1_223 ( );
FILL FILL_1_OAI21X1_223 ( );
FILL FILL_0_OAI21X1_95 ( );
FILL FILL_1_OAI21X1_95 ( );
FILL FILL_0_OAI21X1_94 ( );
FILL FILL_1_OAI21X1_94 ( );
FILL FILL_0_BUFX4_178 ( );
FILL FILL_1_BUFX4_178 ( );
FILL FILL_0_DFFPOSX1_711 ( );
FILL FILL_1_DFFPOSX1_711 ( );
FILL FILL_2_DFFPOSX1_711 ( );
FILL FILL_3_DFFPOSX1_711 ( );
FILL FILL_4_DFFPOSX1_711 ( );
FILL FILL_5_DFFPOSX1_711 ( );
FILL FILL_6_DFFPOSX1_711 ( );
FILL FILL_0_OAI21X1_970 ( );
FILL FILL_1_OAI21X1_970 ( );
FILL FILL_0_NAND2X1_733 ( );
FILL FILL_0_OAI21X1_971 ( );
FILL FILL_1_OAI21X1_971 ( );
FILL FILL_0_DFFPOSX1_77 ( );
FILL FILL_1_DFFPOSX1_77 ( );
FILL FILL_2_DFFPOSX1_77 ( );
FILL FILL_3_DFFPOSX1_77 ( );
FILL FILL_4_DFFPOSX1_77 ( );
FILL FILL_5_DFFPOSX1_77 ( );
FILL FILL_0_OAI21X1_1728 ( );
FILL FILL_1_OAI21X1_1728 ( );
FILL FILL_0_OAI21X1_1729 ( );
FILL FILL_1_OAI21X1_1729 ( );
FILL FILL_2_OAI21X1_1729 ( );
FILL FILL_0_NAND2X1_531 ( );
FILL FILL_1_NAND2X1_531 ( );
FILL FILL_0_OAI21X1_1740 ( );
FILL FILL_1_OAI21X1_1740 ( );
FILL FILL_0_OAI21X1_1677 ( );
FILL FILL_1_OAI21X1_1677 ( );
FILL FILL_0_OAI21X1_1676 ( );
FILL FILL_1_OAI21X1_1676 ( );
FILL FILL_0_DFFPOSX1_234 ( );
FILL FILL_1_DFFPOSX1_234 ( );
FILL FILL_2_DFFPOSX1_234 ( );
FILL FILL_3_DFFPOSX1_234 ( );
FILL FILL_4_DFFPOSX1_234 ( );
FILL FILL_5_DFFPOSX1_234 ( );
FILL FILL_6_DFFPOSX1_234 ( );
FILL FILL_0_OAI21X1_85 ( );
FILL FILL_1_OAI21X1_85 ( );
FILL FILL_0_OAI21X1_84 ( );
FILL FILL_1_OAI21X1_84 ( );
FILL FILL_2_OAI21X1_84 ( );
FILL FILL_0_OAI21X1_1646 ( );
FILL FILL_1_OAI21X1_1646 ( );
FILL FILL_0_DFFPOSX1_36 ( );
FILL FILL_1_DFFPOSX1_36 ( );
FILL FILL_2_DFFPOSX1_36 ( );
FILL FILL_3_DFFPOSX1_36 ( );
FILL FILL_4_DFFPOSX1_36 ( );
FILL FILL_5_DFFPOSX1_36 ( );
FILL FILL_0_OAI21X1_1628 ( );
FILL FILL_1_OAI21X1_1628 ( );
FILL FILL_0_NAND2X1_696 ( );
FILL FILL_1_NAND2X1_696 ( );
FILL FILL_0_BUFX2_40 ( );
FILL FILL_0_BUFX2_1005 ( );
FILL FILL_0_NAND2X1_664 ( );
FILL FILL_0_DFFPOSX1_1018 ( );
FILL FILL_1_DFFPOSX1_1018 ( );
FILL FILL_2_DFFPOSX1_1018 ( );
FILL FILL_3_DFFPOSX1_1018 ( );
FILL FILL_4_DFFPOSX1_1018 ( );
FILL FILL_5_DFFPOSX1_1018 ( );
FILL FILL_0_OAI21X1_298 ( );
FILL FILL_1_OAI21X1_298 ( );
FILL FILL_2_OAI21X1_298 ( );
FILL FILL_0_OAI21X1_1817 ( );
FILL FILL_1_OAI21X1_1817 ( );
FILL FILL_2_OAI21X1_1817 ( );
FILL FILL_0_NAND2X1_758 ( );
FILL FILL_0_BUFX2_687 ( );
FILL FILL_1_BUFX2_687 ( );
FILL FILL_0_OAI21X1_1714 ( );
FILL FILL_1_OAI21X1_1714 ( );
FILL FILL_0_DFFPOSX1_70 ( );
FILL FILL_1_DFFPOSX1_70 ( );
FILL FILL_2_DFFPOSX1_70 ( );
FILL FILL_3_DFFPOSX1_70 ( );
FILL FILL_4_DFFPOSX1_70 ( );
FILL FILL_5_DFFPOSX1_70 ( );
FILL FILL_6_DFFPOSX1_70 ( );
FILL FILL_0_OAI21X1_1715 ( );
FILL FILL_1_OAI21X1_1715 ( );
FILL FILL_0_BUFX4_349 ( );
FILL FILL_1_BUFX4_349 ( );
FILL FILL_0_BUFX2_732 ( );
FILL FILL_0_NAND2X1_652 ( );
FILL FILL_1_NAND2X1_652 ( );
FILL FILL_0_OAI21X1_1583 ( );
FILL FILL_1_OAI21X1_1583 ( );
FILL FILL_0_DFFPOSX1_1006 ( );
FILL FILL_1_DFFPOSX1_1006 ( );
FILL FILL_2_DFFPOSX1_1006 ( );
FILL FILL_3_DFFPOSX1_1006 ( );
FILL FILL_4_DFFPOSX1_1006 ( );
FILL FILL_5_DFFPOSX1_1006 ( );
FILL FILL_6_DFFPOSX1_1006 ( );
FILL FILL_0_NAND2X1_51 ( );
FILL FILL_1_NAND2X1_51 ( );
FILL FILL_0_DFFPOSX1_176 ( );
FILL FILL_1_DFFPOSX1_176 ( );
FILL FILL_2_DFFPOSX1_176 ( );
FILL FILL_3_DFFPOSX1_176 ( );
FILL FILL_4_DFFPOSX1_176 ( );
FILL FILL_5_DFFPOSX1_176 ( );
FILL FILL_6_DFFPOSX1_176 ( );
FILL FILL_0_INVX2_184 ( );
FILL FILL_1_INVX2_184 ( );
FILL FILL_0_BUFX2_879 ( );
FILL FILL_1_BUFX2_879 ( );
FILL FILL_0_BUFX2_679 ( );
FILL FILL_1_BUFX2_679 ( );
FILL FILL_0_OAI21X1_888 ( );
FILL FILL_1_OAI21X1_888 ( );
FILL FILL_0_NAND2X1_382 ( );
FILL FILL_0_BUFX2_291 ( );
FILL FILL_1_BUFX2_291 ( );
FILL FILL_0_BUFX2_270 ( );
FILL FILL_1_BUFX2_270 ( );
FILL FILL_0_DFFPOSX1_630 ( );
FILL FILL_1_DFFPOSX1_630 ( );
FILL FILL_2_DFFPOSX1_630 ( );
FILL FILL_3_DFFPOSX1_630 ( );
FILL FILL_4_DFFPOSX1_630 ( );
FILL FILL_5_DFFPOSX1_630 ( );
FILL FILL_0_INVX2_138 ( );
FILL FILL_0_BUFX2_727 ( );
FILL FILL_0_INVX1_151 ( );
FILL FILL_0_INVX1_165 ( );
FILL FILL_0_OAI21X1_1688 ( );
FILL FILL_1_OAI21X1_1688 ( );
FILL FILL_0_OAI21X1_1689 ( );
FILL FILL_1_OAI21X1_1689 ( );
FILL FILL_0_INVX1_150 ( );
FILL FILL_0_BUFX2_388 ( );
FILL FILL_1_BUFX2_388 ( );
FILL FILL_0_DFFPOSX1_154 ( );
FILL FILL_1_DFFPOSX1_154 ( );
FILL FILL_2_DFFPOSX1_154 ( );
FILL FILL_3_DFFPOSX1_154 ( );
FILL FILL_4_DFFPOSX1_154 ( );
FILL FILL_5_DFFPOSX1_154 ( );
FILL FILL_6_DFFPOSX1_154 ( );
FILL FILL_0_NAND2X1_769 ( );
FILL FILL_1_NAND2X1_769 ( );
FILL FILL_0_OAI21X1_1828 ( );
FILL FILL_1_OAI21X1_1828 ( );
FILL FILL_0_BUFX2_716 ( );
FILL FILL_0_BUFX2_852 ( );
FILL FILL_0_DFFPOSX1_325 ( );
FILL FILL_1_DFFPOSX1_325 ( );
FILL FILL_2_DFFPOSX1_325 ( );
FILL FILL_3_DFFPOSX1_325 ( );
FILL FILL_4_DFFPOSX1_325 ( );
FILL FILL_5_DFFPOSX1_325 ( );
FILL FILL_6_DFFPOSX1_325 ( );
FILL FILL_0_OAI21X1_267 ( );
FILL FILL_1_OAI21X1_267 ( );
FILL FILL_0_BUFX4_368 ( );
FILL FILL_1_BUFX4_368 ( );
FILL FILL_0_OAI21X1_115 ( );
FILL FILL_1_OAI21X1_115 ( );
FILL FILL_0_DFFPOSX1_249 ( );
FILL FILL_1_DFFPOSX1_249 ( );
FILL FILL_2_DFFPOSX1_249 ( );
FILL FILL_3_DFFPOSX1_249 ( );
FILL FILL_4_DFFPOSX1_249 ( );
FILL FILL_5_DFFPOSX1_249 ( );
FILL FILL_0_CLKBUF1_101 ( );
FILL FILL_1_CLKBUF1_101 ( );
FILL FILL_2_CLKBUF1_101 ( );
FILL FILL_3_CLKBUF1_101 ( );
FILL FILL_0_DFFPOSX1_878 ( );
FILL FILL_1_DFFPOSX1_878 ( );
FILL FILL_2_DFFPOSX1_878 ( );
FILL FILL_3_DFFPOSX1_878 ( );
FILL FILL_4_DFFPOSX1_878 ( );
FILL FILL_5_DFFPOSX1_878 ( );
FILL FILL_6_DFFPOSX1_878 ( );
FILL FILL_0_OAI21X1_1678 ( );
FILL FILL_1_OAI21X1_1678 ( );
FILL FILL_0_OAI21X1_1679 ( );
FILL FILL_1_OAI21X1_1679 ( );
FILL FILL_2_OAI21X1_1679 ( );
FILL FILL_0_BUFX4_126 ( );
FILL FILL_1_BUFX4_126 ( );
FILL FILL_0_OAI21X1_1398 ( );
FILL FILL_1_OAI21X1_1398 ( );
FILL FILL_0_OAI21X1_1224 ( );
FILL FILL_1_OAI21X1_1224 ( );
FILL FILL_2_OAI21X1_1224 ( );
FILL FILL_0_OAI21X1_1222 ( );
FILL FILL_1_OAI21X1_1222 ( );
FILL FILL_0_NAND2X1_591 ( );
FILL FILL_1_NAND2X1_591 ( );
FILL FILL_0_NOR2X1_124 ( );
FILL FILL_1_NOR2X1_124 ( );
FILL FILL_0_OAI21X1_1105 ( );
FILL FILL_1_OAI21X1_1105 ( );
FILL FILL_0_DFFPOSX1_813 ( );
FILL FILL_1_DFFPOSX1_813 ( );
FILL FILL_2_DFFPOSX1_813 ( );
FILL FILL_3_DFFPOSX1_813 ( );
FILL FILL_4_DFFPOSX1_813 ( );
FILL FILL_5_DFFPOSX1_813 ( );
FILL FILL_6_DFFPOSX1_813 ( );
FILL FILL_0_INVX2_61 ( );
FILL FILL_1_INVX2_61 ( );
FILL FILL_0_INVX4_47 ( );
FILL FILL_0_OAI21X1_1110 ( );
FILL FILL_1_OAI21X1_1110 ( );
FILL FILL_0_BUFX4_132 ( );
FILL FILL_1_BUFX4_132 ( );
FILL FILL_0_OAI21X1_231 ( );
FILL FILL_1_OAI21X1_231 ( );
FILL FILL_0_DFFPOSX1_307 ( );
FILL FILL_1_DFFPOSX1_307 ( );
FILL FILL_2_DFFPOSX1_307 ( );
FILL FILL_3_DFFPOSX1_307 ( );
FILL FILL_4_DFFPOSX1_307 ( );
FILL FILL_5_DFFPOSX1_307 ( );
FILL FILL_0_NAND2X1_592 ( );
FILL FILL_1_NAND2X1_592 ( );
FILL FILL_0_INVX2_93 ( );
FILL FILL_0_BUFX4_382 ( );
FILL FILL_1_BUFX4_382 ( );
FILL FILL_2_BUFX4_382 ( );
FILL FILL_0_BUFX2_389 ( );
FILL FILL_0_DFFPOSX1_542 ( );
FILL FILL_1_DFFPOSX1_542 ( );
FILL FILL_2_DFFPOSX1_542 ( );
FILL FILL_3_DFFPOSX1_542 ( );
FILL FILL_4_DFFPOSX1_542 ( );
FILL FILL_5_DFFPOSX1_542 ( );
FILL FILL_6_DFFPOSX1_542 ( );
FILL FILL_0_OAI21X1_644 ( );
FILL FILL_1_OAI21X1_644 ( );
FILL FILL_0_OAI21X1_646 ( );
FILL FILL_1_OAI21X1_646 ( );
FILL FILL_2_OAI21X1_646 ( );
FILL FILL_0_AOI21X1_24 ( );
FILL FILL_1_AOI21X1_24 ( );
FILL FILL_0_DFFPOSX1_820 ( );
FILL FILL_1_DFFPOSX1_820 ( );
FILL FILL_2_DFFPOSX1_820 ( );
FILL FILL_3_DFFPOSX1_820 ( );
FILL FILL_4_DFFPOSX1_820 ( );
FILL FILL_5_DFFPOSX1_820 ( );
FILL FILL_0_DFFPOSX1_884 ( );
FILL FILL_1_DFFPOSX1_884 ( );
FILL FILL_2_DFFPOSX1_884 ( );
FILL FILL_3_DFFPOSX1_884 ( );
FILL FILL_4_DFFPOSX1_884 ( );
FILL FILL_5_DFFPOSX1_884 ( );
FILL FILL_6_DFFPOSX1_884 ( );
FILL FILL_0_OAI21X1_1241 ( );
FILL FILL_1_OAI21X1_1241 ( );
FILL FILL_2_OAI21X1_1241 ( );
FILL FILL_0_OAI21X1_1239 ( );
FILL FILL_1_OAI21X1_1239 ( );
FILL FILL_0_INVX4_33 ( );
FILL FILL_1_INVX4_33 ( );
FILL FILL_0_OAI21X1_1238 ( );
FILL FILL_1_OAI21X1_1238 ( );
FILL FILL_0_NOR2X1_98 ( );
FILL FILL_0_BUFX4_246 ( );
FILL FILL_1_BUFX4_246 ( );
FILL FILL_0_OAI21X1_1123 ( );
FILL FILL_1_OAI21X1_1123 ( );
FILL FILL_0_BUFX2_1000 ( );
FILL FILL_0_NOR2X1_100 ( );
FILL FILL_1_NOR2X1_100 ( );
FILL FILL_0_OAI21X1_654 ( );
FILL FILL_1_OAI21X1_654 ( );
FILL FILL_0_BUFX2_199 ( );
FILL FILL_0_AOI21X1_26 ( );
FILL FILL_1_AOI21X1_26 ( );
FILL FILL_0_CLKBUF1_70 ( );
FILL FILL_1_CLKBUF1_70 ( );
FILL FILL_2_CLKBUF1_70 ( );
FILL FILL_3_CLKBUF1_70 ( );
FILL FILL_4_CLKBUF1_70 ( );
FILL FILL_0_DFFPOSX1_822 ( );
FILL FILL_1_DFFPOSX1_822 ( );
FILL FILL_2_DFFPOSX1_822 ( );
FILL FILL_3_DFFPOSX1_822 ( );
FILL FILL_4_DFFPOSX1_822 ( );
FILL FILL_5_DFFPOSX1_822 ( );
FILL FILL_6_DFFPOSX1_822 ( );
FILL FILL_0_OAI21X1_1125 ( );
FILL FILL_1_OAI21X1_1125 ( );
FILL FILL_0_NAND2X1_490 ( );
FILL FILL_0_OAI21X1_112 ( );
FILL FILL_1_OAI21X1_112 ( );
FILL FILL_0_XNOR2X1_77 ( );
FILL FILL_1_XNOR2X1_77 ( );
FILL FILL_2_XNOR2X1_77 ( );
FILL FILL_3_XNOR2X1_77 ( );
FILL FILL_0_NAND2X1_415 ( );
FILL FILL_1_NAND2X1_415 ( );
FILL FILL_0_BUFX4_385 ( );
FILL FILL_1_BUFX4_385 ( );
FILL FILL_0_INVX2_67 ( );
FILL FILL_0_DFFPOSX1_758 ( );
FILL FILL_1_DFFPOSX1_758 ( );
FILL FILL_2_DFFPOSX1_758 ( );
FILL FILL_3_DFFPOSX1_758 ( );
FILL FILL_4_DFFPOSX1_758 ( );
FILL FILL_5_DFFPOSX1_758 ( );
FILL FILL_0_BUFX2_904 ( );
FILL FILL_0_OAI21X1_1051 ( );
FILL FILL_1_OAI21X1_1051 ( );
FILL FILL_0_NAND2X1_417 ( );
FILL FILL_1_NAND2X1_417 ( );
FILL FILL_0_BUFX2_616 ( );
FILL FILL_1_BUFX2_616 ( );
FILL FILL_0_NAND2X1_597 ( );
FILL FILL_1_NAND2X1_597 ( );
FILL FILL_0_NAND2X1_596 ( );
FILL FILL_1_NAND2X1_596 ( );
FILL FILL_0_NAND2X1_8 ( );
FILL FILL_1_NAND2X1_8 ( );
FILL FILL_0_OAI21X1_8 ( );
FILL FILL_1_OAI21X1_8 ( );
FILL FILL_0_OAI21X1_1053 ( );
FILL FILL_1_OAI21X1_1053 ( );
FILL FILL_0_NAND2X1_419 ( );
FILL FILL_1_NAND2X1_419 ( );
FILL FILL_0_BUFX4_359 ( );
FILL FILL_1_BUFX4_359 ( );
FILL FILL_0_DFFPOSX1_258 ( );
FILL FILL_1_DFFPOSX1_258 ( );
FILL FILL_2_DFFPOSX1_258 ( );
FILL FILL_3_DFFPOSX1_258 ( );
FILL FILL_4_DFFPOSX1_258 ( );
FILL FILL_5_DFFPOSX1_258 ( );
FILL FILL_6_DFFPOSX1_258 ( );
FILL FILL_0_BUFX4_164 ( );
FILL FILL_1_BUFX4_164 ( );
FILL FILL_0_NAND2X1_672 ( );
FILL FILL_0_OAI21X1_1603 ( );
FILL FILL_1_OAI21X1_1603 ( );
FILL FILL_0_BUFX2_905 ( );
FILL FILL_1_BUFX2_905 ( );
FILL FILL_0_OAI21X1_1764 ( );
FILL FILL_1_OAI21X1_1764 ( );
FILL FILL_0_DFFPOSX1_180 ( );
FILL FILL_1_DFFPOSX1_180 ( );
FILL FILL_2_DFFPOSX1_180 ( );
FILL FILL_3_DFFPOSX1_180 ( );
FILL FILL_4_DFFPOSX1_180 ( );
FILL FILL_5_DFFPOSX1_180 ( );
FILL FILL_6_DFFPOSX1_180 ( );
FILL FILL_0_BUFX2_216 ( );
FILL FILL_1_BUFX2_216 ( );
FILL FILL_0_DFFPOSX1_1031 ( );
FILL FILL_1_DFFPOSX1_1031 ( );
FILL FILL_2_DFFPOSX1_1031 ( );
FILL FILL_3_DFFPOSX1_1031 ( );
FILL FILL_4_DFFPOSX1_1031 ( );
FILL FILL_5_DFFPOSX1_1031 ( );
FILL FILL_0_BUFX2_696 ( );
FILL FILL_0_DFFPOSX1_275 ( );
FILL FILL_1_DFFPOSX1_275 ( );
FILL FILL_2_DFFPOSX1_275 ( );
FILL FILL_3_DFFPOSX1_275 ( );
FILL FILL_4_DFFPOSX1_275 ( );
FILL FILL_5_DFFPOSX1_275 ( );
FILL FILL_0_OAI21X1_167 ( );
FILL FILL_1_OAI21X1_167 ( );
FILL FILL_0_DFFPOSX1_147 ( );
FILL FILL_1_DFFPOSX1_147 ( );
FILL FILL_2_DFFPOSX1_147 ( );
FILL FILL_3_DFFPOSX1_147 ( );
FILL FILL_4_DFFPOSX1_147 ( );
FILL FILL_5_DFFPOSX1_147 ( );
FILL FILL_0_OAI21X1_295 ( );
FILL FILL_1_OAI21X1_295 ( );
FILL FILL_0_OAI21X1_294 ( );
FILL FILL_1_OAI21X1_294 ( );
FILL FILL_0_BUFX4_361 ( );
FILL FILL_1_BUFX4_361 ( );
FILL FILL_0_BUFX2_85 ( );
FILL FILL_0_OAI21X1_289 ( );
FILL FILL_1_OAI21X1_289 ( );
FILL FILL_0_NAND2X1_759 ( );
FILL FILL_0_DFFPOSX1_336 ( );
FILL FILL_1_DFFPOSX1_336 ( );
FILL FILL_2_DFFPOSX1_336 ( );
FILL FILL_3_DFFPOSX1_336 ( );
FILL FILL_4_DFFPOSX1_336 ( );
FILL FILL_5_DFFPOSX1_336 ( );
FILL FILL_6_DFFPOSX1_336 ( );
FILL FILL_0_DFFPOSX1_318 ( );
FILL FILL_1_DFFPOSX1_318 ( );
FILL FILL_2_DFFPOSX1_318 ( );
FILL FILL_3_DFFPOSX1_318 ( );
FILL FILL_4_DFFPOSX1_318 ( );
FILL FILL_5_DFFPOSX1_318 ( );
FILL FILL_0_NAND2X1_763 ( );
FILL FILL_1_NAND2X1_763 ( );
FILL FILL_0_OAI21X1_1822 ( );
FILL FILL_1_OAI21X1_1822 ( );
FILL FILL_0_DFFPOSX1_276 ( );
FILL FILL_1_DFFPOSX1_276 ( );
FILL FILL_2_DFFPOSX1_276 ( );
FILL FILL_3_DFFPOSX1_276 ( );
FILL FILL_4_DFFPOSX1_276 ( );
FILL FILL_5_DFFPOSX1_276 ( );
FILL FILL_6_DFFPOSX1_276 ( );
FILL FILL_0_OAI21X1_1066 ( );
FILL FILL_1_OAI21X1_1066 ( );
FILL FILL_0_NAND2X1_432 ( );
FILL FILL_1_NAND2X1_432 ( );
FILL FILL_0_BUFX4_220 ( );
FILL FILL_1_BUFX4_220 ( );
FILL FILL_0_NAND2X1_515 ( );
FILL FILL_1_NAND2X1_515 ( );
FILL FILL_0_BUFX2_948 ( );
FILL FILL_0_BUFX2_906 ( );
FILL FILL_0_BUFX2_87 ( );
FILL FILL_0_OAI21X1_1681 ( );
FILL FILL_1_OAI21X1_1681 ( );
FILL FILL_0_OAI21X1_1680 ( );
FILL FILL_1_OAI21X1_1680 ( );
FILL FILL_0_BUFX2_1007 ( );
FILL FILL_1_BUFX2_1007 ( );
FILL FILL_0_DFFPOSX1_345 ( );
FILL FILL_1_DFFPOSX1_345 ( );
FILL FILL_2_DFFPOSX1_345 ( );
FILL FILL_3_DFFPOSX1_345 ( );
FILL FILL_4_DFFPOSX1_345 ( );
FILL FILL_5_DFFPOSX1_345 ( );
FILL FILL_6_DFFPOSX1_345 ( );
FILL FILL_0_DFFPOSX1_281 ( );
FILL FILL_1_DFFPOSX1_281 ( );
FILL FILL_2_DFFPOSX1_281 ( );
FILL FILL_3_DFFPOSX1_281 ( );
FILL FILL_4_DFFPOSX1_281 ( );
FILL FILL_5_DFFPOSX1_281 ( );
FILL FILL_0_DFFPOSX1_936 ( );
FILL FILL_1_DFFPOSX1_936 ( );
FILL FILL_2_DFFPOSX1_936 ( );
FILL FILL_3_DFFPOSX1_936 ( );
FILL FILL_4_DFFPOSX1_936 ( );
FILL FILL_5_DFFPOSX1_936 ( );
FILL FILL_6_DFFPOSX1_936 ( );
FILL FILL_0_BUFX4_172 ( );
FILL FILL_1_BUFX4_172 ( );
FILL FILL_0_OAI21X1_1741 ( );
FILL FILL_1_OAI21X1_1741 ( );
FILL FILL_0_DFFPOSX1_83 ( );
FILL FILL_1_DFFPOSX1_83 ( );
FILL FILL_2_DFFPOSX1_83 ( );
FILL FILL_3_DFFPOSX1_83 ( );
FILL FILL_4_DFFPOSX1_83 ( );
FILL FILL_5_DFFPOSX1_83 ( );
FILL FILL_6_DFFPOSX1_83 ( );
FILL FILL_0_BUFX2_105 ( );
FILL FILL_0_DFFPOSX1_4 ( );
FILL FILL_1_DFFPOSX1_4 ( );
FILL FILL_2_DFFPOSX1_4 ( );
FILL FILL_3_DFFPOSX1_4 ( );
FILL FILL_4_DFFPOSX1_4 ( );
FILL FILL_5_DFFPOSX1_4 ( );
FILL FILL_0_OAI21X1_1614 ( );
FILL FILL_1_OAI21X1_1614 ( );
FILL FILL_0_BUFX2_157 ( );
FILL FILL_0_OAI21X1_1647 ( );
FILL FILL_1_OAI21X1_1647 ( );
FILL FILL_2_OAI21X1_1647 ( );
FILL FILL_0_DFFPOSX1_251 ( );
FILL FILL_1_DFFPOSX1_251 ( );
FILL FILL_2_DFFPOSX1_251 ( );
FILL FILL_3_DFFPOSX1_251 ( );
FILL FILL_4_DFFPOSX1_251 ( );
FILL FILL_5_DFFPOSX1_251 ( );
FILL FILL_0_DFFPOSX1_138 ( );
FILL FILL_1_DFFPOSX1_138 ( );
FILL FILL_2_DFFPOSX1_138 ( );
FILL FILL_3_DFFPOSX1_138 ( );
FILL FILL_4_DFFPOSX1_138 ( );
FILL FILL_5_DFFPOSX1_138 ( );
FILL FILL_0_OAI21X1_1581 ( );
FILL FILL_1_OAI21X1_1581 ( );
FILL FILL_2_OAI21X1_1581 ( );
FILL FILL_0_NAND2X1_650 ( );
FILL FILL_0_OAI21X1_1812 ( );
FILL FILL_1_OAI21X1_1812 ( );
FILL FILL_0_NAND2X1_753 ( );
FILL FILL_0_DFFPOSX1_266 ( );
FILL FILL_1_DFFPOSX1_266 ( );
FILL FILL_2_DFFPOSX1_266 ( );
FILL FILL_3_DFFPOSX1_266 ( );
FILL FILL_4_DFFPOSX1_266 ( );
FILL FILL_5_DFFPOSX1_266 ( );
FILL FILL_0_DFFPOSX1_1014 ( );
FILL FILL_1_DFFPOSX1_1014 ( );
FILL FILL_2_DFFPOSX1_1014 ( );
FILL FILL_3_DFFPOSX1_1014 ( );
FILL FILL_4_DFFPOSX1_1014 ( );
FILL FILL_5_DFFPOSX1_1014 ( );
FILL FILL_6_DFFPOSX1_1014 ( );
FILL FILL_0_OAI21X1_1591 ( );
FILL FILL_1_OAI21X1_1591 ( );
FILL FILL_0_NAND2X1_660 ( );
FILL FILL_1_NAND2X1_660 ( );
FILL FILL_0_CLKBUF1_99 ( );
FILL FILL_1_CLKBUF1_99 ( );
FILL FILL_2_CLKBUF1_99 ( );
FILL FILL_3_CLKBUF1_99 ( );
FILL FILL_4_CLKBUF1_99 ( );
FILL FILL_0_OAI21X1_1607 ( );
FILL FILL_1_OAI21X1_1607 ( );
FILL FILL_2_OAI21X1_1607 ( );
FILL FILL_0_NAND2X1_676 ( );
FILL FILL_0_DFFPOSX1_1030 ( );
FILL FILL_1_DFFPOSX1_1030 ( );
FILL FILL_2_DFFPOSX1_1030 ( );
FILL FILL_3_DFFPOSX1_1030 ( );
FILL FILL_4_DFFPOSX1_1030 ( );
FILL FILL_5_DFFPOSX1_1030 ( );
FILL FILL_6_DFFPOSX1_1030 ( );
FILL FILL_0_BUFX2_815 ( );
FILL FILL_0_OAI21X1_20 ( );
FILL FILL_1_OAI21X1_20 ( );
FILL FILL_0_NAND2X1_20 ( );
FILL FILL_0_OAI21X1_46 ( );
FILL FILL_1_OAI21X1_46 ( );
FILL FILL_0_NAND2X1_46 ( );
FILL FILL_0_DFFPOSX1_202 ( );
FILL FILL_1_DFFPOSX1_202 ( );
FILL FILL_2_DFFPOSX1_202 ( );
FILL FILL_3_DFFPOSX1_202 ( );
FILL FILL_4_DFFPOSX1_202 ( );
FILL FILL_5_DFFPOSX1_202 ( );
FILL FILL_6_DFFPOSX1_202 ( );
FILL FILL_0_BUFX2_1013 ( );
FILL FILL_0_BUFX2_328 ( );
FILL FILL_1_BUFX2_328 ( );
FILL FILL_0_BUFX2_267 ( );
FILL FILL_0_INVX1_59 ( );
FILL FILL_0_OAI21X1_858 ( );
FILL FILL_1_OAI21X1_858 ( );
FILL FILL_0_BUFX2_374 ( );
FILL FILL_1_BUFX2_374 ( );
FILL FILL_0_DFFPOSX1_688 ( );
FILL FILL_1_DFFPOSX1_688 ( );
FILL FILL_2_DFFPOSX1_688 ( );
FILL FILL_3_DFFPOSX1_688 ( );
FILL FILL_4_DFFPOSX1_688 ( );
FILL FILL_5_DFFPOSX1_688 ( );
FILL FILL_0_OAI21X1_925 ( );
FILL FILL_1_OAI21X1_925 ( );
FILL FILL_0_OAI21X1_924 ( );
FILL FILL_1_OAI21X1_924 ( );
FILL FILL_0_OAI21X1_933 ( );
FILL FILL_1_OAI21X1_933 ( );
FILL FILL_2_OAI21X1_933 ( );
FILL FILL_0_OAI21X1_932 ( );
FILL FILL_1_OAI21X1_932 ( );
FILL FILL_0_DFFPOSX1_692 ( );
FILL FILL_1_DFFPOSX1_692 ( );
FILL FILL_2_DFFPOSX1_692 ( );
FILL FILL_3_DFFPOSX1_692 ( );
FILL FILL_4_DFFPOSX1_692 ( );
FILL FILL_5_DFFPOSX1_692 ( );
FILL FILL_6_DFFPOSX1_692 ( );
FILL FILL_0_DFFPOSX1_197 ( );
FILL FILL_1_DFFPOSX1_197 ( );
FILL FILL_2_DFFPOSX1_197 ( );
FILL FILL_3_DFFPOSX1_197 ( );
FILL FILL_4_DFFPOSX1_197 ( );
FILL FILL_5_DFFPOSX1_197 ( );
FILL FILL_0_NAND2X1_41 ( );
FILL FILL_0_OAI21X1_41 ( );
FILL FILL_1_OAI21X1_41 ( );
FILL FILL_2_OAI21X1_41 ( );
FILL FILL_0_BUFX2_891 ( );
FILL FILL_0_BUFX4_143 ( );
FILL FILL_1_BUFX4_143 ( );
FILL FILL_0_BUFX4_329 ( );
FILL FILL_1_BUFX4_329 ( );
FILL FILL_0_NAND2X1_62 ( );
FILL FILL_1_NAND2X1_62 ( );
FILL FILL_0_OAI21X1_62 ( );
FILL FILL_1_OAI21X1_62 ( );
FILL FILL_0_OAI21X1_114 ( );
FILL FILL_1_OAI21X1_114 ( );
FILL FILL_0_DFFPOSX1_218 ( );
FILL FILL_1_DFFPOSX1_218 ( );
FILL FILL_2_DFFPOSX1_218 ( );
FILL FILL_3_DFFPOSX1_218 ( );
FILL FILL_4_DFFPOSX1_218 ( );
FILL FILL_5_DFFPOSX1_218 ( );
FILL FILL_0_OAI21X1_951 ( );
FILL FILL_1_OAI21X1_951 ( );
FILL FILL_0_OAI21X1_950 ( );
FILL FILL_1_OAI21X1_950 ( );
FILL FILL_0_DFFPOSX1_701 ( );
FILL FILL_1_DFFPOSX1_701 ( );
FILL FILL_2_DFFPOSX1_701 ( );
FILL FILL_3_DFFPOSX1_701 ( );
FILL FILL_4_DFFPOSX1_701 ( );
FILL FILL_5_DFFPOSX1_701 ( );
FILL FILL_0_BUFX2_174 ( );
FILL FILL_1_BUFX2_174 ( );
FILL FILL_0_BUFX4_8 ( );
FILL FILL_1_BUFX4_8 ( );
FILL FILL_0_OAI21X1_1743 ( );
FILL FILL_1_OAI21X1_1743 ( );
FILL FILL_0_OAI21X1_1216 ( );
FILL FILL_1_OAI21X1_1216 ( );
FILL FILL_0_OAI21X1_1223 ( );
FILL FILL_1_OAI21X1_1223 ( );
FILL FILL_0_OAI21X1_1217 ( );
FILL FILL_1_OAI21X1_1217 ( );
FILL FILL_0_NAND2X1_474 ( );
FILL FILL_0_BUFX4_249 ( );
FILL FILL_1_BUFX4_249 ( );
FILL FILL_0_DFFPOSX1_879 ( );
FILL FILL_1_DFFPOSX1_879 ( );
FILL FILL_2_DFFPOSX1_879 ( );
FILL FILL_3_DFFPOSX1_879 ( );
FILL FILL_4_DFFPOSX1_879 ( );
FILL FILL_5_DFFPOSX1_879 ( );
FILL FILL_0_OAI21X1_1227 ( );
FILL FILL_1_OAI21X1_1227 ( );
FILL FILL_2_OAI21X1_1227 ( );
FILL FILL_0_NOR2X1_178 ( );
FILL FILL_0_OAI21X1_1225 ( );
FILL FILL_1_OAI21X1_1225 ( );
FILL FILL_0_NAND2X1_473 ( );
FILL FILL_0_NAND2X1_480 ( );
FILL FILL_1_NAND2X1_480 ( );
FILL FILL_0_OAI21X1_1229 ( );
FILL FILL_1_OAI21X1_1229 ( );
FILL FILL_0_OAI21X1_1228 ( );
FILL FILL_1_OAI21X1_1228 ( );
FILL FILL_0_BUFX2_254 ( );
FILL FILL_0_NOR2X1_125 ( );
FILL FILL_1_NOR2X1_125 ( );
FILL FILL_0_BUFX2_131 ( );
FILL FILL_0_NOR2X1_180 ( );
FILL FILL_0_NAND2X1_593 ( );
FILL FILL_1_NAND2X1_593 ( );
FILL FILL_0_NOR2X1_126 ( );
FILL FILL_0_OAI21X1_1116 ( );
FILL FILL_1_OAI21X1_1116 ( );
FILL FILL_0_BUFX2_574 ( );
FILL FILL_1_BUFX2_574 ( );
FILL FILL_0_DFFPOSX1_816 ( );
FILL FILL_1_DFFPOSX1_816 ( );
FILL FILL_2_DFFPOSX1_816 ( );
FILL FILL_3_DFFPOSX1_816 ( );
FILL FILL_4_DFFPOSX1_816 ( );
FILL FILL_5_DFFPOSX1_816 ( );
FILL FILL_0_BUFX2_390 ( );
FILL FILL_1_BUFX2_390 ( );
FILL FILL_0_CLKBUF1_74 ( );
FILL FILL_1_CLKBUF1_74 ( );
FILL FILL_2_CLKBUF1_74 ( );
FILL FILL_3_CLKBUF1_74 ( );
FILL FILL_4_CLKBUF1_74 ( );
FILL FILL_0_BUFX2_69 ( );
FILL FILL_0_BUFX4_198 ( );
FILL FILL_1_BUFX4_198 ( );
FILL FILL_0_OAI21X1_1630 ( );
FILL FILL_1_OAI21X1_1630 ( );
FILL FILL_0_NAND2X1_698 ( );
FILL FILL_1_NAND2X1_698 ( );
FILL FILL_0_DFFPOSX1_20 ( );
FILL FILL_1_DFFPOSX1_20 ( );
FILL FILL_2_DFFPOSX1_20 ( );
FILL FILL_3_DFFPOSX1_20 ( );
FILL FILL_4_DFFPOSX1_20 ( );
FILL FILL_5_DFFPOSX1_20 ( );
FILL FILL_6_DFFPOSX1_20 ( );
FILL FILL_0_OAI21X1_1240 ( );
FILL FILL_1_OAI21X1_1240 ( );
FILL FILL_0_OAI21X1_647 ( );
FILL FILL_1_OAI21X1_647 ( );
FILL FILL_0_OAI21X1_649 ( );
FILL FILL_1_OAI21X1_649 ( );
FILL FILL_0_OAI21X1_648 ( );
FILL FILL_1_OAI21X1_648 ( );
FILL FILL_0_INVX2_64 ( );
FILL FILL_0_BUFX2_452 ( );
FILL FILL_1_BUFX2_452 ( );
FILL FILL_0_INVX1_4 ( );
FILL FILL_0_XNOR2X1_76 ( );
FILL FILL_1_XNOR2X1_76 ( );
FILL FILL_2_XNOR2X1_76 ( );
FILL FILL_3_XNOR2X1_76 ( );
FILL FILL_0_OAI21X1_652 ( );
FILL FILL_1_OAI21X1_652 ( );
FILL FILL_0_DFFPOSX1_545 ( );
FILL FILL_1_DFFPOSX1_545 ( );
FILL FILL_2_DFFPOSX1_545 ( );
FILL FILL_3_DFFPOSX1_545 ( );
FILL FILL_4_DFFPOSX1_545 ( );
FILL FILL_5_DFFPOSX1_545 ( );
FILL FILL_0_OAI21X1_657 ( );
FILL FILL_1_OAI21X1_657 ( );
FILL FILL_2_OAI21X1_657 ( );
FILL FILL_0_DFFPOSX1_546 ( );
FILL FILL_1_DFFPOSX1_546 ( );
FILL FILL_2_DFFPOSX1_546 ( );
FILL FILL_3_DFFPOSX1_546 ( );
FILL FILL_4_DFFPOSX1_546 ( );
FILL FILL_5_DFFPOSX1_546 ( );
FILL FILL_6_DFFPOSX1_546 ( );
FILL FILL_0_NAND2X1_493 ( );
FILL FILL_1_NAND2X1_493 ( );
FILL FILL_0_OAI21X1_1128 ( );
FILL FILL_1_OAI21X1_1128 ( );
FILL FILL_0_BUFX2_918 ( );
FILL FILL_1_BUFX2_918 ( );
FILL FILL_0_BUFX2_72 ( );
FILL FILL_0_BUFX4_235 ( );
FILL FILL_1_BUFX4_235 ( );
FILL FILL_2_BUFX4_235 ( );
FILL FILL_0_BUFX2_468 ( );
FILL FILL_1_BUFX2_468 ( );
FILL FILL_0_BUFX2_6 ( );
FILL FILL_1_BUFX2_6 ( );
FILL FILL_0_OAI21X1_1258 ( );
FILL FILL_1_OAI21X1_1258 ( );
FILL FILL_0_BUFX2_9 ( );
FILL FILL_0_NAND2X1_416 ( );
FILL FILL_1_NAND2X1_416 ( );
FILL FILL_0_DFFPOSX1_759 ( );
FILL FILL_1_DFFPOSX1_759 ( );
FILL FILL_2_DFFPOSX1_759 ( );
FILL FILL_3_DFFPOSX1_759 ( );
FILL FILL_4_DFFPOSX1_759 ( );
FILL FILL_5_DFFPOSX1_759 ( );
FILL FILL_6_DFFPOSX1_759 ( );
FILL FILL_0_DFFPOSX1_164 ( );
FILL FILL_1_DFFPOSX1_164 ( );
FILL FILL_2_DFFPOSX1_164 ( );
FILL FILL_3_DFFPOSX1_164 ( );
FILL FILL_4_DFFPOSX1_164 ( );
FILL FILL_5_DFFPOSX1_164 ( );
FILL FILL_0_DFFPOSX1_761 ( );
FILL FILL_1_DFFPOSX1_761 ( );
FILL FILL_2_DFFPOSX1_761 ( );
FILL FILL_3_DFFPOSX1_761 ( );
FILL FILL_4_DFFPOSX1_761 ( );
FILL FILL_5_DFFPOSX1_761 ( );
FILL FILL_6_DFFPOSX1_761 ( );
FILL FILL_0_BUFX2_73 ( );
FILL FILL_1_BUFX2_73 ( );
FILL FILL_0_OAI21X1_133 ( );
FILL FILL_1_OAI21X1_133 ( );
FILL FILL_0_OAI21X1_132 ( );
FILL FILL_1_OAI21X1_132 ( );
FILL FILL_0_BUFX4_110 ( );
FILL FILL_1_BUFX4_110 ( );
FILL FILL_0_DFFPOSX1_1026 ( );
FILL FILL_1_DFFPOSX1_1026 ( );
FILL FILL_2_DFFPOSX1_1026 ( );
FILL FILL_3_DFFPOSX1_1026 ( );
FILL FILL_4_DFFPOSX1_1026 ( );
FILL FILL_5_DFFPOSX1_1026 ( );
FILL FILL_0_BUFX2_763 ( );
FILL FILL_0_DFFPOSX1_725 ( );
FILL FILL_1_DFFPOSX1_725 ( );
FILL FILL_2_DFFPOSX1_725 ( );
FILL FILL_3_DFFPOSX1_725 ( );
FILL FILL_4_DFFPOSX1_725 ( );
FILL FILL_5_DFFPOSX1_725 ( );
FILL FILL_0_BUFX2_765 ( );
FILL FILL_1_BUFX2_765 ( );
FILL FILL_0_OAI21X1_1691 ( );
FILL FILL_1_OAI21X1_1691 ( );
FILL FILL_0_NAND2X1_356 ( );
FILL FILL_0_NAND2X1_677 ( );
FILL FILL_0_DFFPOSX1_58 ( );
FILL FILL_1_DFFPOSX1_58 ( );
FILL FILL_2_DFFPOSX1_58 ( );
FILL FILL_3_DFFPOSX1_58 ( );
FILL FILL_4_DFFPOSX1_58 ( );
FILL FILL_5_DFFPOSX1_58 ( );
FILL FILL_0_BUFX2_669 ( );
FILL FILL_1_BUFX2_669 ( );
FILL FILL_0_BUFX2_760 ( );
FILL FILL_1_BUFX2_760 ( );
FILL FILL_0_OAI21X1_166 ( );
FILL FILL_1_OAI21X1_166 ( );
FILL FILL_0_BUFX2_871 ( );
FILL FILL_1_BUFX2_871 ( );
FILL FILL_0_OAI21X1_1821 ( );
FILL FILL_1_OAI21X1_1821 ( );
FILL FILL_0_NAND2X1_762 ( );
FILL FILL_1_NAND2X1_762 ( );
FILL FILL_0_OAI21X1_1208 ( );
FILL FILL_1_OAI21X1_1208 ( );
FILL FILL_0_DFFPOSX1_872 ( );
FILL FILL_1_DFFPOSX1_872 ( );
FILL FILL_2_DFFPOSX1_872 ( );
FILL FILL_3_DFFPOSX1_872 ( );
FILL FILL_4_DFFPOSX1_872 ( );
FILL FILL_5_DFFPOSX1_872 ( );
FILL FILL_0_OAI21X1_1209 ( );
FILL FILL_1_OAI21X1_1209 ( );
FILL FILL_0_OAI21X1_160 ( );
FILL FILL_1_OAI21X1_160 ( );
FILL FILL_0_OAI21X1_1818 ( );
FILL FILL_1_OAI21X1_1818 ( );
FILL FILL_0_DFFPOSX1_144 ( );
FILL FILL_1_DFFPOSX1_144 ( );
FILL FILL_2_DFFPOSX1_144 ( );
FILL FILL_3_DFFPOSX1_144 ( );
FILL FILL_4_DFFPOSX1_144 ( );
FILL FILL_5_DFFPOSX1_144 ( );
FILL FILL_0_OAI21X1_252 ( );
FILL FILL_1_OAI21X1_252 ( );
FILL FILL_0_OAI21X1_124 ( );
FILL FILL_1_OAI21X1_124 ( );
FILL FILL_0_OAI21X1_125 ( );
FILL FILL_1_OAI21X1_125 ( );
FILL FILL_0_OAI21X1_253 ( );
FILL FILL_1_OAI21X1_253 ( );
FILL FILL_2_OAI21X1_253 ( );
FILL FILL_0_BUFX2_1008 ( );
FILL FILL_0_DFFPOSX1_774 ( );
FILL FILL_1_DFFPOSX1_774 ( );
FILL FILL_2_DFFPOSX1_774 ( );
FILL FILL_3_DFFPOSX1_774 ( );
FILL FILL_4_DFFPOSX1_774 ( );
FILL FILL_5_DFFPOSX1_774 ( );
FILL FILL_6_DFFPOSX1_774 ( );
FILL FILL_0_DFFPOSX1_832 ( );
FILL FILL_1_DFFPOSX1_832 ( );
FILL FILL_2_DFFPOSX1_832 ( );
FILL FILL_3_DFFPOSX1_832 ( );
FILL FILL_4_DFFPOSX1_832 ( );
FILL FILL_5_DFFPOSX1_832 ( );
FILL FILL_6_DFFPOSX1_832 ( );
FILL FILL_0_BUFX2_213 ( );
FILL FILL_1_BUFX2_213 ( );
FILL FILL_0_BUFX2_972 ( );
FILL FILL_1_BUFX2_972 ( );
FILL FILL_0_OAI21X1_862 ( );
FILL FILL_1_OAI21X1_862 ( );
FILL FILL_0_BUFX2_762 ( );
FILL FILL_1_BUFX2_762 ( );
FILL FILL_0_BUFX2_722 ( );
FILL FILL_0_BUFX2_754 ( );
FILL FILL_1_BUFX2_754 ( );
FILL FILL_0_OAI21X1_307 ( );
FILL FILL_1_OAI21X1_307 ( );
FILL FILL_0_OAI21X1_306 ( );
FILL FILL_1_OAI21X1_306 ( );
FILL FILL_0_OAI21X1_179 ( );
FILL FILL_1_OAI21X1_179 ( );
FILL FILL_0_OAI21X1_178 ( );
FILL FILL_1_OAI21X1_178 ( );
FILL FILL_0_BUFX2_787 ( );
FILL FILL_0_BUFX2_954 ( );
FILL FILL_1_BUFX2_954 ( );
FILL FILL_0_OAI21X1_1384 ( );
FILL FILL_1_OAI21X1_1384 ( );
FILL FILL_0_OAI21X1_1385 ( );
FILL FILL_1_OAI21X1_1385 ( );
FILL FILL_0_OAI21X1_246 ( );
FILL FILL_1_OAI21X1_246 ( );
FILL FILL_2_OAI21X1_246 ( );
FILL FILL_0_BUFX2_776 ( );
FILL FILL_0_DFFPOSX1_315 ( );
FILL FILL_1_DFFPOSX1_315 ( );
FILL FILL_2_DFFPOSX1_315 ( );
FILL FILL_3_DFFPOSX1_315 ( );
FILL FILL_4_DFFPOSX1_315 ( );
FILL FILL_5_DFFPOSX1_315 ( );
FILL FILL_6_DFFPOSX1_315 ( );
FILL FILL_0_OAI21X1_247 ( );
FILL FILL_1_OAI21X1_247 ( );
FILL FILL_0_BUFX2_91 ( );
FILL FILL_1_BUFX2_91 ( );
FILL FILL_0_CLKBUF1_25 ( );
FILL FILL_1_CLKBUF1_25 ( );
FILL FILL_2_CLKBUF1_25 ( );
FILL FILL_3_CLKBUF1_25 ( );
FILL FILL_4_CLKBUF1_25 ( );
FILL FILL_0_BUFX2_237 ( );
FILL FILL_1_BUFX2_237 ( );
FILL FILL_0_NAND2X1_682 ( );
FILL FILL_0_BUFX2_681 ( );
FILL FILL_1_BUFX2_681 ( );
FILL FILL_0_CLKBUF1_17 ( );
FILL FILL_1_CLKBUF1_17 ( );
FILL FILL_2_CLKBUF1_17 ( );
FILL FILL_3_CLKBUF1_17 ( );
FILL FILL_0_OAI21X1_119 ( );
FILL FILL_1_OAI21X1_119 ( );
FILL FILL_0_OAI21X1_118 ( );
FILL FILL_1_OAI21X1_118 ( );
FILL FILL_0_BUFX4_322 ( );
FILL FILL_1_BUFX4_322 ( );
FILL FILL_0_BUFX2_713 ( );
FILL FILL_1_BUFX2_713 ( );
FILL FILL_0_DFFPOSX1_1004 ( );
FILL FILL_1_DFFPOSX1_1004 ( );
FILL FILL_2_DFFPOSX1_1004 ( );
FILL FILL_3_DFFPOSX1_1004 ( );
FILL FILL_4_DFFPOSX1_1004 ( );
FILL FILL_5_DFFPOSX1_1004 ( );
FILL FILL_6_DFFPOSX1_1004 ( );
FILL FILL_0_BUFX2_655 ( );
FILL FILL_1_BUFX2_655 ( );
FILL FILL_0_OAI21X1_148 ( );
FILL FILL_1_OAI21X1_148 ( );
FILL FILL_0_OAI21X1_149 ( );
FILL FILL_1_OAI21X1_149 ( );
FILL FILL_2_OAI21X1_149 ( );
FILL FILL_0_OAI21X1_1730 ( );
FILL FILL_1_OAI21X1_1730 ( );
FILL FILL_0_DFFPOSX1_78 ( );
FILL FILL_1_DFFPOSX1_78 ( );
FILL FILL_2_DFFPOSX1_78 ( );
FILL FILL_3_DFFPOSX1_78 ( );
FILL FILL_4_DFFPOSX1_78 ( );
FILL FILL_5_DFFPOSX1_78 ( );
FILL FILL_6_DFFPOSX1_78 ( );
FILL FILL_0_OAI21X1_1731 ( );
FILL FILL_1_OAI21X1_1731 ( );
FILL FILL_0_BUFX2_747 ( );
FILL FILL_1_BUFX2_747 ( );
FILL FILL_0_CLKBUF1_32 ( );
FILL FILL_1_CLKBUF1_32 ( );
FILL FILL_2_CLKBUF1_32 ( );
FILL FILL_3_CLKBUF1_32 ( );
FILL FILL_4_CLKBUF1_32 ( );
FILL FILL_0_BUFX2_757 ( );
FILL FILL_1_BUFX2_757 ( );
FILL FILL_0_BUFX4_227 ( );
FILL FILL_1_BUFX4_227 ( );
FILL FILL_0_BUFX2_661 ( );
FILL FILL_1_BUFX2_661 ( );
FILL FILL_0_OAI21X1_1640 ( );
FILL FILL_1_OAI21X1_1640 ( );
FILL FILL_0_NAND2X1_708 ( );
FILL FILL_0_DFFPOSX1_30 ( );
FILL FILL_1_DFFPOSX1_30 ( );
FILL FILL_2_DFFPOSX1_30 ( );
FILL FILL_3_DFFPOSX1_30 ( );
FILL FILL_4_DFFPOSX1_30 ( );
FILL FILL_5_DFFPOSX1_30 ( );
FILL FILL_0_DFFPOSX1_640 ( );
FILL FILL_1_DFFPOSX1_640 ( );
FILL FILL_2_DFFPOSX1_640 ( );
FILL FILL_3_DFFPOSX1_640 ( );
FILL FILL_4_DFFPOSX1_640 ( );
FILL FILL_5_DFFPOSX1_640 ( );
FILL FILL_6_DFFPOSX1_640 ( );
FILL FILL_0_OAI21X1_868 ( );
FILL FILL_1_OAI21X1_868 ( );
FILL FILL_2_OAI21X1_868 ( );
FILL FILL_0_INVX1_69 ( );
FILL FILL_0_INVX2_127 ( );
FILL FILL_0_NAND2X1_362 ( );
FILL FILL_0_BUFX2_873 ( );
FILL FILL_1_BUFX2_873 ( );
FILL FILL_0_BUFX2_355 ( );
FILL FILL_0_INVX1_97 ( );
FILL FILL_0_INVX1_117 ( );
FILL FILL_0_OAI21X1_896 ( );
FILL FILL_1_OAI21X1_896 ( );
FILL FILL_0_NAND2X1_390 ( );
FILL FILL_1_NAND2X1_390 ( );
FILL FILL_0_DFFPOSX1_668 ( );
FILL FILL_1_DFFPOSX1_668 ( );
FILL FILL_2_DFFPOSX1_668 ( );
FILL FILL_3_DFFPOSX1_668 ( );
FILL FILL_4_DFFPOSX1_668 ( );
FILL FILL_5_DFFPOSX1_668 ( );
FILL FILL_6_DFFPOSX1_668 ( );
FILL FILL_0_INVX1_121 ( );
FILL FILL_0_INVX2_183 ( );
FILL FILL_0_INVX1_166 ( );
FILL FILL_1_INVX1_166 ( );
FILL FILL_0_BUFX4_184 ( );
FILL FILL_1_BUFX4_184 ( );
FILL FILL_0_OAI21X1_884 ( );
FILL FILL_1_OAI21X1_884 ( );
FILL FILL_0_DFFPOSX1_656 ( );
FILL FILL_1_DFFPOSX1_656 ( );
FILL FILL_2_DFFPOSX1_656 ( );
FILL FILL_3_DFFPOSX1_656 ( );
FILL FILL_4_DFFPOSX1_656 ( );
FILL FILL_5_DFFPOSX1_656 ( );
FILL FILL_0_OAI21X1_1811 ( );
FILL FILL_1_OAI21X1_1811 ( );
FILL FILL_0_NAND2X1_752 ( );
FILL FILL_0_DFFPOSX1_137 ( );
FILL FILL_1_DFFPOSX1_137 ( );
FILL FILL_2_DFFPOSX1_137 ( );
FILL FILL_3_DFFPOSX1_137 ( );
FILL FILL_4_DFFPOSX1_137 ( );
FILL FILL_5_DFFPOSX1_137 ( );
FILL FILL_6_DFFPOSX1_137 ( );
FILL FILL_0_INVX1_130 ( );
FILL FILL_0_DFFPOSX1_121 ( );
FILL FILL_1_DFFPOSX1_121 ( );
FILL FILL_2_DFFPOSX1_121 ( );
FILL FILL_3_DFFPOSX1_121 ( );
FILL FILL_4_DFFPOSX1_121 ( );
FILL FILL_5_DFFPOSX1_121 ( );
FILL FILL_0_OAI21X1_1795 ( );
FILL FILL_1_OAI21X1_1795 ( );
FILL FILL_0_BUFX4_247 ( );
FILL FILL_1_BUFX4_247 ( );
FILL FILL_0_BUFX2_339 ( );
FILL FILL_0_OAI21X1_1789 ( );
FILL FILL_1_OAI21X1_1789 ( );
FILL FILL_0_NAND2X1_730 ( );
FILL FILL_1_NAND2X1_730 ( );
FILL FILL_0_OAI21X1_1609 ( );
FILL FILL_1_OAI21X1_1609 ( );
FILL FILL_0_NAND2X1_678 ( );
FILL FILL_1_NAND2X1_678 ( );
FILL FILL_0_CLKBUF1_39 ( );
FILL FILL_1_CLKBUF1_39 ( );
FILL FILL_2_CLKBUF1_39 ( );
FILL FILL_3_CLKBUF1_39 ( );
FILL FILL_4_CLKBUF1_39 ( );
FILL FILL_0_INVX8_5 ( );
FILL FILL_1_INVX8_5 ( );
FILL FILL_2_INVX8_5 ( );
FILL FILL_0_DFFPOSX1_84 ( );
FILL FILL_1_DFFPOSX1_84 ( );
FILL FILL_2_DFFPOSX1_84 ( );
FILL FILL_3_DFFPOSX1_84 ( );
FILL FILL_4_DFFPOSX1_84 ( );
FILL FILL_5_DFFPOSX1_84 ( );
FILL FILL_0_OAI21X1_1742 ( );
FILL FILL_1_OAI21X1_1742 ( );
FILL FILL_2_OAI21X1_1742 ( );
FILL FILL_0_BUFX2_190 ( );
FILL FILL_1_BUFX2_190 ( );
FILL FILL_0_OAI21X1_1226 ( );
FILL FILL_1_OAI21X1_1226 ( );
FILL FILL_0_OAI21X1_908 ( );
FILL FILL_1_OAI21X1_908 ( );
FILL FILL_0_OAI21X1_1230 ( );
FILL FILL_1_OAI21X1_1230 ( );
FILL FILL_0_DFFPOSX1_880 ( );
FILL FILL_1_DFFPOSX1_880 ( );
FILL FILL_2_DFFPOSX1_880 ( );
FILL FILL_3_DFFPOSX1_880 ( );
FILL FILL_4_DFFPOSX1_880 ( );
FILL FILL_5_DFFPOSX1_880 ( );
FILL FILL_6_DFFPOSX1_880 ( );
FILL FILL_0_OAI21X1_1231 ( );
FILL FILL_1_OAI21X1_1231 ( );
FILL FILL_0_INVX2_60 ( );
FILL FILL_0_NAND2X1_410 ( );
FILL FILL_0_OAI21X1_1044 ( );
FILL FILL_1_OAI21X1_1044 ( );
FILL FILL_0_OAI21X1_102 ( );
FILL FILL_1_OAI21X1_102 ( );
FILL FILL_0_OAI21X1_103 ( );
FILL FILL_1_OAI21X1_103 ( );
FILL FILL_2_OAI21X1_103 ( );
FILL FILL_0_DFFPOSX1_243 ( );
FILL FILL_1_DFFPOSX1_243 ( );
FILL FILL_2_DFFPOSX1_243 ( );
FILL FILL_3_DFFPOSX1_243 ( );
FILL FILL_4_DFFPOSX1_243 ( );
FILL FILL_5_DFFPOSX1_243 ( );
FILL FILL_6_DFFPOSX1_243 ( );
FILL FILL_0_BUFX4_353 ( );
FILL FILL_1_BUFX4_353 ( );
FILL FILL_0_NAND2X1_479 ( );
FILL FILL_0_OAI21X1_1039 ( );
FILL FILL_1_OAI21X1_1039 ( );
FILL FILL_0_NAND2X1_405 ( );
FILL FILL_1_NAND2X1_405 ( );
FILL FILL_0_DFFPOSX1_747 ( );
FILL FILL_1_DFFPOSX1_747 ( );
FILL FILL_2_DFFPOSX1_747 ( );
FILL FILL_3_DFFPOSX1_747 ( );
FILL FILL_4_DFFPOSX1_747 ( );
FILL FILL_5_DFFPOSX1_747 ( );
FILL FILL_0_BUFX2_3 ( );
FILL FILL_1_BUFX2_3 ( );
FILL FILL_0_INVX4_26 ( );
FILL FILL_0_BUFX4_312 ( );
FILL FILL_1_BUFX4_312 ( );
FILL FILL_0_OAI21X1_1236 ( );
FILL FILL_1_OAI21X1_1236 ( );
FILL FILL_0_DFFPOSX1_883 ( );
FILL FILL_1_DFFPOSX1_883 ( );
FILL FILL_2_DFFPOSX1_883 ( );
FILL FILL_3_DFFPOSX1_883 ( );
FILL FILL_4_DFFPOSX1_883 ( );
FILL FILL_5_DFFPOSX1_883 ( );
FILL FILL_0_OAI21X1_1237 ( );
FILL FILL_1_OAI21X1_1237 ( );
FILL FILL_0_CLKBUF1_11 ( );
FILL FILL_1_CLKBUF1_11 ( );
FILL FILL_2_CLKBUF1_11 ( );
FILL FILL_3_CLKBUF1_11 ( );
FILL FILL_4_CLKBUF1_11 ( );
FILL FILL_0_DFFPOSX1_543 ( );
FILL FILL_1_DFFPOSX1_543 ( );
FILL FILL_2_DFFPOSX1_543 ( );
FILL FILL_3_DFFPOSX1_543 ( );
FILL FILL_4_DFFPOSX1_543 ( );
FILL FILL_5_DFFPOSX1_543 ( );
FILL FILL_0_BUFX4_386 ( );
FILL FILL_1_BUFX4_386 ( );
FILL FILL_0_OAI21X1_1048 ( );
FILL FILL_1_OAI21X1_1048 ( );
FILL FILL_0_NAND2X1_414 ( );
FILL FILL_1_NAND2X1_414 ( );
FILL FILL_0_BUFX2_936 ( );
FILL FILL_1_BUFX2_936 ( );
FILL FILL_0_OAI21X1_1047 ( );
FILL FILL_1_OAI21X1_1047 ( );
FILL FILL_0_NAND2X1_413 ( );
FILL FILL_0_NAND2X1_265 ( );
FILL FILL_1_NAND2X1_265 ( );
FILL FILL_0_NAND2X1_264 ( );
FILL FILL_1_NAND2X1_264 ( );
FILL FILL_0_CLKBUF1_65 ( );
FILL FILL_1_CLKBUF1_65 ( );
FILL FILL_2_CLKBUF1_65 ( );
FILL FILL_3_CLKBUF1_65 ( );
FILL FILL_4_CLKBUF1_65 ( );
FILL FILL_0_BUFX4_101 ( );
FILL FILL_1_BUFX4_101 ( );
FILL FILL_0_OAI21X1_655 ( );
FILL FILL_1_OAI21X1_655 ( );
FILL FILL_0_BUFX4_10 ( );
FILL FILL_1_BUFX4_10 ( );
FILL FILL_0_BUFX4_250 ( );
FILL FILL_1_BUFX4_250 ( );
FILL FILL_0_OAI21X1_1250 ( );
FILL FILL_1_OAI21X1_1250 ( );
FILL FILL_0_OAI21X1_1251 ( );
FILL FILL_1_OAI21X1_1251 ( );
FILL FILL_0_OAI21X1_1257 ( );
FILL FILL_1_OAI21X1_1257 ( );
FILL FILL_0_DFFPOSX1_889 ( );
FILL FILL_1_DFFPOSX1_889 ( );
FILL FILL_2_DFFPOSX1_889 ( );
FILL FILL_3_DFFPOSX1_889 ( );
FILL FILL_4_DFFPOSX1_889 ( );
FILL FILL_5_DFFPOSX1_889 ( );
FILL FILL_6_DFFPOSX1_889 ( );
FILL FILL_0_DFFPOSX1_278 ( );
FILL FILL_1_DFFPOSX1_278 ( );
FILL FILL_2_DFFPOSX1_278 ( );
FILL FILL_3_DFFPOSX1_278 ( );
FILL FILL_4_DFFPOSX1_278 ( );
FILL FILL_5_DFFPOSX1_278 ( );
FILL FILL_6_DFFPOSX1_278 ( );
FILL FILL_0_DFFPOSX1_194 ( );
FILL FILL_1_DFFPOSX1_194 ( );
FILL FILL_2_DFFPOSX1_194 ( );
FILL FILL_3_DFFPOSX1_194 ( );
FILL FILL_4_DFFPOSX1_194 ( );
FILL FILL_5_DFFPOSX1_194 ( );
FILL FILL_0_BUFX2_10 ( );
FILL FILL_1_BUFX2_10 ( );
FILL FILL_0_BUFX2_412 ( );
FILL FILL_0_DFFPOSX1_150 ( );
FILL FILL_1_DFFPOSX1_150 ( );
FILL FILL_2_DFFPOSX1_150 ( );
FILL FILL_3_DFFPOSX1_150 ( );
FILL FILL_4_DFFPOSX1_150 ( );
FILL FILL_5_DFFPOSX1_150 ( );
FILL FILL_6_DFFPOSX1_150 ( );
FILL FILL_0_OAI21X1_184 ( );
FILL FILL_1_OAI21X1_184 ( );
FILL FILL_0_DFFPOSX1_284 ( );
FILL FILL_1_DFFPOSX1_284 ( );
FILL FILL_2_DFFPOSX1_284 ( );
FILL FILL_3_DFFPOSX1_284 ( );
FILL FILL_4_DFFPOSX1_284 ( );
FILL FILL_5_DFFPOSX1_284 ( );
FILL FILL_6_DFFPOSX1_284 ( );
FILL FILL_0_OAI21X1_185 ( );
FILL FILL_1_OAI21X1_185 ( );
FILL FILL_0_DFFPOSX1_252 ( );
FILL FILL_1_DFFPOSX1_252 ( );
FILL FILL_2_DFFPOSX1_252 ( );
FILL FILL_3_DFFPOSX1_252 ( );
FILL FILL_4_DFFPOSX1_252 ( );
FILL FILL_5_DFFPOSX1_252 ( );
FILL FILL_6_DFFPOSX1_252 ( );
FILL FILL_0_BUFX4_248 ( );
FILL FILL_1_BUFX4_248 ( );
FILL FILL_2_BUFX4_248 ( );
FILL FILL_0_OAI21X1_998 ( );
FILL FILL_1_OAI21X1_998 ( );
FILL FILL_0_OAI21X1_999 ( );
FILL FILL_1_OAI21X1_999 ( );
FILL FILL_0_OAI21X1_1690 ( );
FILL FILL_1_OAI21X1_1690 ( );
FILL FILL_0_DFFPOSX1_43 ( );
FILL FILL_1_DFFPOSX1_43 ( );
FILL FILL_2_DFFPOSX1_43 ( );
FILL FILL_3_DFFPOSX1_43 ( );
FILL FILL_4_DFFPOSX1_43 ( );
FILL FILL_5_DFFPOSX1_43 ( );
FILL FILL_0_BUFX2_819 ( );
FILL FILL_1_BUFX2_819 ( );
FILL FILL_0_OAI21X1_1804 ( );
FILL FILL_1_OAI21X1_1804 ( );
FILL FILL_2_OAI21X1_1804 ( );
FILL FILL_0_NAND2X1_745 ( );
FILL FILL_0_DFFPOSX1_130 ( );
FILL FILL_1_DFFPOSX1_130 ( );
FILL FILL_2_DFFPOSX1_130 ( );
FILL FILL_3_DFFPOSX1_130 ( );
FILL FILL_4_DFFPOSX1_130 ( );
FILL FILL_5_DFFPOSX1_130 ( );
FILL FILL_6_DFFPOSX1_130 ( );
FILL FILL_0_OAI21X1_1725 ( );
FILL FILL_1_OAI21X1_1725 ( );
FILL FILL_0_OAI21X1_1724 ( );
FILL FILL_1_OAI21X1_1724 ( );
FILL FILL_0_DFFPOSX1_75 ( );
FILL FILL_1_DFFPOSX1_75 ( );
FILL FILL_2_DFFPOSX1_75 ( );
FILL FILL_3_DFFPOSX1_75 ( );
FILL FILL_4_DFFPOSX1_75 ( );
FILL FILL_5_DFFPOSX1_75 ( );
FILL FILL_0_NAND2X1_33 ( );
FILL FILL_0_OAI21X1_33 ( );
FILL FILL_1_OAI21X1_33 ( );
FILL FILL_0_OAI21X1_161 ( );
FILL FILL_1_OAI21X1_161 ( );
FILL FILL_0_DFFPOSX1_1017 ( );
FILL FILL_1_DFFPOSX1_1017 ( );
FILL FILL_2_DFFPOSX1_1017 ( );
FILL FILL_3_DFFPOSX1_1017 ( );
FILL FILL_4_DFFPOSX1_1017 ( );
FILL FILL_5_DFFPOSX1_1017 ( );
FILL FILL_6_DFFPOSX1_1017 ( );
FILL FILL_0_INVX2_182 ( );
FILL FILL_0_DFFPOSX1_254 ( );
FILL FILL_1_DFFPOSX1_254 ( );
FILL FILL_2_DFFPOSX1_254 ( );
FILL FILL_3_DFFPOSX1_254 ( );
FILL FILL_4_DFFPOSX1_254 ( );
FILL FILL_5_DFFPOSX1_254 ( );
FILL FILL_6_DFFPOSX1_254 ( );
FILL FILL_0_BUFX4_363 ( );
FILL FILL_1_BUFX4_363 ( );
FILL FILL_2_BUFX4_363 ( );
FILL FILL_0_BUFX4_191 ( );
FILL FILL_1_BUFX4_191 ( );
FILL FILL_0_OAI21X1_56 ( );
FILL FILL_1_OAI21X1_56 ( );
FILL FILL_0_NAND2X1_56 ( );
FILL FILL_1_NAND2X1_56 ( );
FILL FILL_0_DFFPOSX1_212 ( );
FILL FILL_1_DFFPOSX1_212 ( );
FILL FILL_2_DFFPOSX1_212 ( );
FILL FILL_3_DFFPOSX1_212 ( );
FILL FILL_4_DFFPOSX1_212 ( );
FILL FILL_5_DFFPOSX1_212 ( );
FILL FILL_0_BUFX2_25 ( );
FILL FILL_0_INVX1_63 ( );
FILL FILL_0_DFFPOSX1_634 ( );
FILL FILL_1_DFFPOSX1_634 ( );
FILL FILL_2_DFFPOSX1_634 ( );
FILL FILL_3_DFFPOSX1_634 ( );
FILL FILL_4_DFFPOSX1_634 ( );
FILL FILL_5_DFFPOSX1_634 ( );
FILL FILL_0_OAI21X1_1598 ( );
FILL FILL_1_OAI21X1_1598 ( );
FILL FILL_2_OAI21X1_1598 ( );
FILL FILL_0_DFFPOSX1_1021 ( );
FILL FILL_1_DFFPOSX1_1021 ( );
FILL FILL_2_DFFPOSX1_1021 ( );
FILL FILL_3_DFFPOSX1_1021 ( );
FILL FILL_4_DFFPOSX1_1021 ( );
FILL FILL_5_DFFPOSX1_1021 ( );
FILL FILL_6_DFFPOSX1_1021 ( );
FILL FILL_0_DFFPOSX1_271 ( );
FILL FILL_1_DFFPOSX1_271 ( );
FILL FILL_2_DFFPOSX1_271 ( );
FILL FILL_3_DFFPOSX1_271 ( );
FILL FILL_4_DFFPOSX1_271 ( );
FILL FILL_5_DFFPOSX1_271 ( );
FILL FILL_6_DFFPOSX1_271 ( );
FILL FILL_0_DFFPOSX1_214 ( );
FILL FILL_1_DFFPOSX1_214 ( );
FILL FILL_2_DFFPOSX1_214 ( );
FILL FILL_3_DFFPOSX1_214 ( );
FILL FILL_4_DFFPOSX1_214 ( );
FILL FILL_5_DFFPOSX1_214 ( );
FILL FILL_0_BUFX4_218 ( );
FILL FILL_1_BUFX4_218 ( );
FILL FILL_0_BUFX2_193 ( );
FILL FILL_1_BUFX2_193 ( );
FILL FILL_0_BUFX2_985 ( );
FILL FILL_1_BUFX2_985 ( );
FILL FILL_0_BUFX2_752 ( );
FILL FILL_1_BUFX2_752 ( );
FILL FILL_0_DFFPOSX1_326 ( );
FILL FILL_1_DFFPOSX1_326 ( );
FILL FILL_2_DFFPOSX1_326 ( );
FILL FILL_3_DFFPOSX1_326 ( );
FILL FILL_4_DFFPOSX1_326 ( );
FILL FILL_5_DFFPOSX1_326 ( );
FILL FILL_0_BUFX4_165 ( );
FILL FILL_1_BUFX4_165 ( );
FILL FILL_0_BUFX2_720 ( );
FILL FILL_1_BUFX2_720 ( );
FILL FILL_0_BUFX4_234 ( );
FILL FILL_1_BUFX4_234 ( );
FILL FILL_0_DFFPOSX1_68 ( );
FILL FILL_1_DFFPOSX1_68 ( );
FILL FILL_2_DFFPOSX1_68 ( );
FILL FILL_3_DFFPOSX1_68 ( );
FILL FILL_4_DFFPOSX1_68 ( );
FILL FILL_5_DFFPOSX1_68 ( );
FILL FILL_6_DFFPOSX1_68 ( );
FILL FILL_0_DFFPOSX1_240 ( );
FILL FILL_1_DFFPOSX1_240 ( );
FILL FILL_2_DFFPOSX1_240 ( );
FILL FILL_3_DFFPOSX1_240 ( );
FILL FILL_4_DFFPOSX1_240 ( );
FILL FILL_5_DFFPOSX1_240 ( );
FILL FILL_0_BUFX2_961 ( );
FILL FILL_0_OAI21X1_1036 ( );
FILL FILL_1_OAI21X1_1036 ( );
FILL FILL_0_NAND2X1_402 ( );
FILL FILL_1_NAND2X1_402 ( );
FILL FILL_0_DFFPOSX1_744 ( );
FILL FILL_1_DFFPOSX1_744 ( );
FILL FILL_2_DFFPOSX1_744 ( );
FILL FILL_3_DFFPOSX1_744 ( );
FILL FILL_4_DFFPOSX1_744 ( );
FILL FILL_5_DFFPOSX1_744 ( );
FILL FILL_6_DFFPOSX1_744 ( );
FILL FILL_0_INVX2_54 ( );
FILL FILL_0_OAI21X1_1100 ( );
FILL FILL_1_OAI21X1_1100 ( );
FILL FILL_0_DFFPOSX1_808 ( );
FILL FILL_1_DFFPOSX1_808 ( );
FILL FILL_2_DFFPOSX1_808 ( );
FILL FILL_3_DFFPOSX1_808 ( );
FILL FILL_4_DFFPOSX1_808 ( );
FILL FILL_5_DFFPOSX1_808 ( );
FILL FILL_0_BUFX4_137 ( );
FILL FILL_1_BUFX4_137 ( );
FILL FILL_2_BUFX4_137 ( );
FILL FILL_0_BUFX4_123 ( );
FILL FILL_1_BUFX4_123 ( );
FILL FILL_0_BUFX4_332 ( );
FILL FILL_1_BUFX4_332 ( );
FILL FILL_0_DFFPOSX1_38 ( );
FILL FILL_1_DFFPOSX1_38 ( );
FILL FILL_2_DFFPOSX1_38 ( );
FILL FILL_3_DFFPOSX1_38 ( );
FILL FILL_4_DFFPOSX1_38 ( );
FILL FILL_5_DFFPOSX1_38 ( );
FILL FILL_0_OAI21X1_1651 ( );
FILL FILL_1_OAI21X1_1651 ( );
FILL FILL_0_OAI21X1_1650 ( );
FILL FILL_1_OAI21X1_1650 ( );
FILL FILL_0_BUFX2_725 ( );
FILL FILL_1_BUFX2_725 ( );
FILL FILL_0_BUFX4_205 ( );
FILL FILL_1_BUFX4_205 ( );
FILL FILL_0_INVX2_169 ( );
FILL FILL_0_INVX2_152 ( );
FILL FILL_0_DFFPOSX1_6 ( );
FILL FILL_1_DFFPOSX1_6 ( );
FILL FILL_2_DFFPOSX1_6 ( );
FILL FILL_3_DFFPOSX1_6 ( );
FILL FILL_4_DFFPOSX1_6 ( );
FILL FILL_5_DFFPOSX1_6 ( );
FILL FILL_0_OAI21X1_1616 ( );
FILL FILL_1_OAI21X1_1616 ( );
FILL FILL_0_NAND2X1_684 ( );
FILL FILL_1_NAND2X1_684 ( );
FILL FILL_0_INVX2_119 ( );
FILL FILL_0_BUFX2_925 ( );
FILL FILL_1_BUFX2_925 ( );
FILL FILL_0_OAI21X1_889 ( );
FILL FILL_1_OAI21X1_889 ( );
FILL FILL_0_BUFX2_877 ( );
FILL FILL_1_BUFX2_877 ( );
FILL FILL_0_INVX1_110 ( );
FILL FILL_0_BUFX2_274 ( );
FILL FILL_0_NAND2X1_352 ( );
FILL FILL_1_NAND2X1_352 ( );
FILL FILL_0_OAI21X1_864 ( );
FILL FILL_1_OAI21X1_864 ( );
FILL FILL_0_INVX1_65 ( );
FILL FILL_0_BUFX2_306 ( );
FILL FILL_0_NAND2X1_346 ( );
FILL FILL_1_NAND2X1_346 ( );
FILL FILL_0_DFFPOSX1_636 ( );
FILL FILL_1_DFFPOSX1_636 ( );
FILL FILL_2_DFFPOSX1_636 ( );
FILL FILL_3_DFFPOSX1_636 ( );
FILL FILL_4_DFFPOSX1_636 ( );
FILL FILL_5_DFFPOSX1_636 ( );
FILL FILL_0_BUFX2_329 ( );
FILL FILL_0_BUFX2_323 ( );
FILL FILL_1_BUFX2_323 ( );
FILL FILL_0_BUFX2_335 ( );
FILL FILL_1_BUFX2_335 ( );
FILL FILL_0_NAND2X1_378 ( );
FILL FILL_1_NAND2X1_378 ( );
FILL FILL_0_BUFX2_827 ( );
FILL FILL_1_BUFX2_827 ( );
FILL FILL_0_BUFX2_808 ( );
FILL FILL_1_BUFX2_808 ( );
FILL FILL_0_OAI21X1_945 ( );
FILL FILL_1_OAI21X1_945 ( );
FILL FILL_0_OAI21X1_944 ( );
FILL FILL_1_OAI21X1_944 ( );
FILL FILL_0_DFFPOSX1_698 ( );
FILL FILL_1_DFFPOSX1_698 ( );
FILL FILL_2_DFFPOSX1_698 ( );
FILL FILL_3_DFFPOSX1_698 ( );
FILL FILL_4_DFFPOSX1_698 ( );
FILL FILL_5_DFFPOSX1_698 ( );
FILL FILL_6_DFFPOSX1_698 ( );
FILL FILL_0_OAI21X1_180 ( );
FILL FILL_1_OAI21X1_180 ( );
FILL FILL_0_BUFX2_791 ( );
FILL FILL_1_BUFX2_791 ( );
FILL FILL_0_NAND2X1_736 ( );
FILL FILL_1_NAND2X1_736 ( );
FILL FILL_0_BUFX2_919 ( );
FILL FILL_0_OAI21X1_181 ( );
FILL FILL_1_OAI21X1_181 ( );
FILL FILL_2_OAI21X1_181 ( );
FILL FILL_0_DFFPOSX1_282 ( );
FILL FILL_1_DFFPOSX1_282 ( );
FILL FILL_2_DFFPOSX1_282 ( );
FILL FILL_3_DFFPOSX1_282 ( );
FILL FILL_4_DFFPOSX1_282 ( );
FILL FILL_5_DFFPOSX1_282 ( );
FILL FILL_6_DFFPOSX1_282 ( );
FILL FILL_0_BUFX2_784 ( );
FILL FILL_0_BUFX2_249 ( );
FILL FILL_1_BUFX2_249 ( );
FILL FILL_0_BUFX4_208 ( );
FILL FILL_1_BUFX4_208 ( );
FILL FILL_0_DFFPOSX1_115 ( );
FILL FILL_1_DFFPOSX1_115 ( );
FILL FILL_2_DFFPOSX1_115 ( );
FILL FILL_3_DFFPOSX1_115 ( );
FILL FILL_4_DFFPOSX1_115 ( );
FILL FILL_5_DFFPOSX1_115 ( );
FILL FILL_6_DFFPOSX1_115 ( );
FILL FILL_0_BUFX2_185 ( );
FILL FILL_1_BUFX2_185 ( );
FILL FILL_0_DFFPOSX1_1032 ( );
FILL FILL_1_DFFPOSX1_1032 ( );
FILL FILL_2_DFFPOSX1_1032 ( );
FILL FILL_3_DFFPOSX1_1032 ( );
FILL FILL_4_DFFPOSX1_1032 ( );
FILL FILL_5_DFFPOSX1_1032 ( );
FILL FILL_6_DFFPOSX1_1032 ( );
FILL FILL_0_DFFPOSX1_876 ( );
FILL FILL_1_DFFPOSX1_876 ( );
FILL FILL_2_DFFPOSX1_876 ( );
FILL FILL_3_DFFPOSX1_876 ( );
FILL FILL_4_DFFPOSX1_876 ( );
FILL FILL_5_DFFPOSX1_876 ( );
FILL FILL_6_DFFPOSX1_876 ( );
FILL FILL_0_OAI21X1_909 ( );
FILL FILL_1_OAI21X1_909 ( );
FILL FILL_0_DFFPOSX1_680 ( );
FILL FILL_1_DFFPOSX1_680 ( );
FILL FILL_2_DFFPOSX1_680 ( );
FILL FILL_3_DFFPOSX1_680 ( );
FILL FILL_4_DFFPOSX1_680 ( );
FILL FILL_5_DFFPOSX1_680 ( );
FILL FILL_0_BUFX2_152 ( );
FILL FILL_0_OAI21X1_1215 ( );
FILL FILL_1_OAI21X1_1215 ( );
FILL FILL_0_DFFPOSX1_875 ( );
FILL FILL_1_DFFPOSX1_875 ( );
FILL FILL_2_DFFPOSX1_875 ( );
FILL FILL_3_DFFPOSX1_875 ( );
FILL FILL_4_DFFPOSX1_875 ( );
FILL FILL_5_DFFPOSX1_875 ( );
FILL FILL_0_OAI21X1_1214 ( );
FILL FILL_1_OAI21X1_1214 ( );
FILL FILL_0_OAI21X1_1043 ( );
FILL FILL_1_OAI21X1_1043 ( );
FILL FILL_0_OAI21X1_1111 ( );
FILL FILL_1_OAI21X1_1111 ( );
FILL FILL_0_BUFX2_980 ( );
FILL FILL_1_BUFX2_980 ( );
FILL FILL_0_DFFPOSX1_752 ( );
FILL FILL_1_DFFPOSX1_752 ( );
FILL FILL_2_DFFPOSX1_752 ( );
FILL FILL_3_DFFPOSX1_752 ( );
FILL FILL_4_DFFPOSX1_752 ( );
FILL FILL_5_DFFPOSX1_752 ( );
FILL FILL_6_DFFPOSX1_752 ( );
FILL FILL_0_XNOR2X1_74 ( );
FILL FILL_1_XNOR2X1_74 ( );
FILL FILL_2_XNOR2X1_74 ( );
FILL FILL_3_XNOR2X1_74 ( );
FILL FILL_0_DFFPOSX1_881 ( );
FILL FILL_1_DFFPOSX1_881 ( );
FILL FILL_2_DFFPOSX1_881 ( );
FILL FILL_3_DFFPOSX1_881 ( );
FILL FILL_4_DFFPOSX1_881 ( );
FILL FILL_5_DFFPOSX1_881 ( );
FILL FILL_0_OAI21X1_1233 ( );
FILL FILL_1_OAI21X1_1233 ( );
FILL FILL_0_OAI21X1_1232 ( );
FILL FILL_1_OAI21X1_1232 ( );
FILL FILL_0_BUFX2_132 ( );
FILL FILL_1_BUFX2_132 ( );
FILL FILL_0_OAI21X1_1712 ( );
FILL FILL_1_OAI21X1_1712 ( );
FILL FILL_0_DFFPOSX1_69 ( );
FILL FILL_1_DFFPOSX1_69 ( );
FILL FILL_2_DFFPOSX1_69 ( );
FILL FILL_3_DFFPOSX1_69 ( );
FILL FILL_4_DFFPOSX1_69 ( );
FILL FILL_5_DFFPOSX1_69 ( );
FILL FILL_0_BUFX2_446 ( );
FILL FILL_0_NAND2X1_130 ( );
FILL FILL_1_NAND2X1_130 ( );
FILL FILL_0_OAI21X1_386 ( );
FILL FILL_1_OAI21X1_386 ( );
FILL FILL_0_BUFX2_133 ( );
FILL FILL_1_BUFX2_133 ( );
FILL FILL_0_BUFX2_67 ( );
FILL FILL_1_BUFX2_67 ( );
FILL FILL_0_BUFX2_68 ( );
FILL FILL_1_BUFX2_68 ( );
FILL FILL_0_BUFX2_644 ( );
FILL FILL_0_BUFX2_581 ( );
FILL FILL_0_OAI21X1_141 ( );
FILL FILL_1_OAI21X1_141 ( );
FILL FILL_0_OAI21X1_140 ( );
FILL FILL_1_OAI21X1_140 ( );
FILL FILL_0_BUFX4_316 ( );
FILL FILL_1_BUFX4_316 ( );
FILL FILL_0_DFFPOSX1_756 ( );
FILL FILL_1_DFFPOSX1_756 ( );
FILL FILL_2_DFFPOSX1_756 ( );
FILL FILL_3_DFFPOSX1_756 ( );
FILL FILL_4_DFFPOSX1_756 ( );
FILL FILL_5_DFFPOSX1_756 ( );
FILL FILL_0_DFFPOSX1_483 ( );
FILL FILL_1_DFFPOSX1_483 ( );
FILL FILL_2_DFFPOSX1_483 ( );
FILL FILL_3_DFFPOSX1_483 ( );
FILL FILL_4_DFFPOSX1_483 ( );
FILL FILL_5_DFFPOSX1_483 ( );
FILL FILL_0_DFFPOSX1_755 ( );
FILL FILL_1_DFFPOSX1_755 ( );
FILL FILL_2_DFFPOSX1_755 ( );
FILL FILL_3_DFFPOSX1_755 ( );
FILL FILL_4_DFFPOSX1_755 ( );
FILL FILL_5_DFFPOSX1_755 ( );
FILL FILL_0_OAI21X1_91 ( );
FILL FILL_1_OAI21X1_91 ( );
FILL FILL_0_OAI21X1_90 ( );
FILL FILL_1_OAI21X1_90 ( );
FILL FILL_2_OAI21X1_90 ( );
FILL FILL_0_BUFX4_94 ( );
FILL FILL_1_BUFX4_94 ( );
FILL FILL_0_BUFX2_488 ( );
FILL FILL_0_OAI21X1_234 ( );
FILL FILL_1_OAI21X1_234 ( );
FILL FILL_0_DFFPOSX1_887 ( );
FILL FILL_1_DFFPOSX1_887 ( );
FILL FILL_2_DFFPOSX1_887 ( );
FILL FILL_3_DFFPOSX1_887 ( );
FILL FILL_4_DFFPOSX1_887 ( );
FILL FILL_5_DFFPOSX1_887 ( );
FILL FILL_6_DFFPOSX1_887 ( );
FILL FILL_0_BUFX2_7 ( );
FILL FILL_0_OAI21X1_172 ( );
FILL FILL_1_OAI21X1_172 ( );
FILL FILL_0_OAI21X1_173 ( );
FILL FILL_1_OAI21X1_173 ( );
FILL FILL_0_DFFPOSX1_740 ( );
FILL FILL_1_DFFPOSX1_740 ( );
FILL FILL_2_DFFPOSX1_740 ( );
FILL FILL_3_DFFPOSX1_740 ( );
FILL FILL_4_DFFPOSX1_740 ( );
FILL FILL_5_DFFPOSX1_740 ( );
FILL FILL_0_BUFX2_841 ( );
FILL FILL_0_NAND2X1_38 ( );
FILL FILL_1_NAND2X1_38 ( );
FILL FILL_0_OAI21X1_38 ( );
FILL FILL_1_OAI21X1_38 ( );
FILL FILL_0_OAI21X1_1824 ( );
FILL FILL_1_OAI21X1_1824 ( );
FILL FILL_0_NAND2X1_765 ( );
FILL FILL_0_BUFX2_823 ( );
FILL FILL_0_BUFX2_916 ( );
FILL FILL_1_BUFX2_916 ( );
FILL FILL_0_DFFPOSX1_348 ( );
FILL FILL_1_DFFPOSX1_348 ( );
FILL FILL_2_DFFPOSX1_348 ( );
FILL FILL_3_DFFPOSX1_348 ( );
FILL FILL_4_DFFPOSX1_348 ( );
FILL FILL_5_DFFPOSX1_348 ( );
FILL FILL_0_OAI21X1_313 ( );
FILL FILL_1_OAI21X1_313 ( );
FILL FILL_0_OAI21X1_312 ( );
FILL FILL_1_OAI21X1_312 ( );
FILL FILL_0_OAI21X1_121 ( );
FILL FILL_1_OAI21X1_121 ( );
FILL FILL_0_OAI21X1_120 ( );
FILL FILL_1_OAI21X1_120 ( );
FILL FILL_0_OAI21X1_186 ( );
FILL FILL_1_OAI21X1_186 ( );
FILL FILL_0_OAI21X1_187 ( );
FILL FILL_1_OAI21X1_187 ( );
FILL FILL_0_BUFX2_203 ( );
FILL FILL_1_BUFX2_203 ( );
FILL FILL_0_OAI21X1_1660 ( );
FILL FILL_1_OAI21X1_1660 ( );
FILL FILL_2_OAI21X1_1660 ( );
FILL FILL_0_OAI21X1_1661 ( );
FILL FILL_1_OAI21X1_1661 ( );
FILL FILL_0_BUFX2_728 ( );
FILL FILL_1_BUFX2_728 ( );
FILL FILL_0_OAI21X1_1798 ( );
FILL FILL_1_OAI21X1_1798 ( );
FILL FILL_0_NAND2X1_739 ( );
FILL FILL_0_DFFPOSX1_124 ( );
FILL FILL_1_DFFPOSX1_124 ( );
FILL FILL_2_DFFPOSX1_124 ( );
FILL FILL_3_DFFPOSX1_124 ( );
FILL FILL_4_DFFPOSX1_124 ( );
FILL FILL_5_DFFPOSX1_124 ( );
FILL FILL_6_DFFPOSX1_124 ( );
FILL FILL_0_OAI21X1_1588 ( );
FILL FILL_1_OAI21X1_1588 ( );
FILL FILL_0_NAND2X1_657 ( );
FILL FILL_1_NAND2X1_657 ( );
FILL FILL_0_BUFX4_336 ( );
FILL FILL_1_BUFX4_336 ( );
FILL FILL_0_BUFX2_774 ( );
FILL FILL_0_BUFX2_129 ( );
FILL FILL_0_DFFPOSX1_189 ( );
FILL FILL_1_DFFPOSX1_189 ( );
FILL FILL_2_DFFPOSX1_189 ( );
FILL FILL_3_DFFPOSX1_189 ( );
FILL FILL_4_DFFPOSX1_189 ( );
FILL FILL_5_DFFPOSX1_189 ( );
FILL FILL_6_DFFPOSX1_189 ( );
FILL FILL_0_DFFPOSX1_272 ( );
FILL FILL_1_DFFPOSX1_272 ( );
FILL FILL_2_DFFPOSX1_272 ( );
FILL FILL_3_DFFPOSX1_272 ( );
FILL FILL_4_DFFPOSX1_272 ( );
FILL FILL_5_DFFPOSX1_272 ( );
FILL FILL_0_NAND2X1_663 ( );
FILL FILL_0_OAI21X1_1594 ( );
FILL FILL_1_OAI21X1_1594 ( );
FILL FILL_2_OAI21X1_1594 ( );
FILL FILL_0_DFFPOSX1_126 ( );
FILL FILL_1_DFFPOSX1_126 ( );
FILL FILL_2_DFFPOSX1_126 ( );
FILL FILL_3_DFFPOSX1_126 ( );
FILL FILL_4_DFFPOSX1_126 ( );
FILL FILL_5_DFFPOSX1_126 ( );
FILL FILL_6_DFFPOSX1_126 ( );
FILL FILL_0_DFFPOSX1_111 ( );
FILL FILL_1_DFFPOSX1_111 ( );
FILL FILL_2_DFFPOSX1_111 ( );
FILL FILL_3_DFFPOSX1_111 ( );
FILL FILL_4_DFFPOSX1_111 ( );
FILL FILL_5_DFFPOSX1_111 ( );
FILL FILL_6_DFFPOSX1_111 ( );
FILL FILL_0_DFFPOSX1_175 ( );
FILL FILL_1_DFFPOSX1_175 ( );
FILL FILL_2_DFFPOSX1_175 ( );
FILL FILL_3_DFFPOSX1_175 ( );
FILL FILL_4_DFFPOSX1_175 ( );
FILL FILL_5_DFFPOSX1_175 ( );
FILL FILL_0_DFFPOSX1_217 ( );
FILL FILL_1_DFFPOSX1_217 ( );
FILL FILL_2_DFFPOSX1_217 ( );
FILL FILL_3_DFFPOSX1_217 ( );
FILL FILL_4_DFFPOSX1_217 ( );
FILL FILL_5_DFFPOSX1_217 ( );
FILL FILL_6_DFFPOSX1_217 ( );
FILL FILL_0_NAND2X1_61 ( );
FILL FILL_1_NAND2X1_61 ( );
FILL FILL_0_OAI21X1_61 ( );
FILL FILL_1_OAI21X1_61 ( );
FILL FILL_0_BUFX4_380 ( );
FILL FILL_1_BUFX4_380 ( );
FILL FILL_0_NAND2X1_667 ( );
FILL FILL_0_DFFPOSX1_1013 ( );
FILL FILL_1_DFFPOSX1_1013 ( );
FILL FILL_2_DFFPOSX1_1013 ( );
FILL FILL_3_DFFPOSX1_1013 ( );
FILL FILL_4_DFFPOSX1_1013 ( );
FILL FILL_5_DFFPOSX1_1013 ( );
FILL FILL_0_OAI21X1_158 ( );
FILL FILL_1_OAI21X1_158 ( );
FILL FILL_0_BUFX2_350 ( );
FILL FILL_0_OAI21X1_159 ( );
FILL FILL_1_OAI21X1_159 ( );
FILL FILL_0_OAI21X1_58 ( );
FILL FILL_1_OAI21X1_58 ( );
FILL FILL_2_OAI21X1_58 ( );
FILL FILL_0_NAND2X1_58 ( );
FILL FILL_0_DFFPOSX1_742 ( );
FILL FILL_1_DFFPOSX1_742 ( );
FILL FILL_2_DFFPOSX1_742 ( );
FILL FILL_3_DFFPOSX1_742 ( );
FILL FILL_4_DFFPOSX1_742 ( );
FILL FILL_5_DFFPOSX1_742 ( );
FILL FILL_0_OAI21X1_1032 ( );
FILL FILL_1_OAI21X1_1032 ( );
FILL FILL_2_OAI21X1_1032 ( );
FILL FILL_0_OAI21X1_1033 ( );
FILL FILL_1_OAI21X1_1033 ( );
FILL FILL_0_BUFX2_381 ( );
FILL FILL_0_OAI21X1_269 ( );
FILL FILL_1_OAI21X1_269 ( );
FILL FILL_0_OAI21X1_268 ( );
FILL FILL_1_OAI21X1_268 ( );
FILL FILL_0_DFFPOSX1_50 ( );
FILL FILL_1_DFFPOSX1_50 ( );
FILL FILL_2_DFFPOSX1_50 ( );
FILL FILL_3_DFFPOSX1_50 ( );
FILL FILL_4_DFFPOSX1_50 ( );
FILL FILL_5_DFFPOSX1_50 ( );
FILL FILL_6_DFFPOSX1_50 ( );
FILL FILL_0_OAI21X1_1675 ( );
FILL FILL_1_OAI21X1_1675 ( );
FILL FILL_0_OAI21X1_1711 ( );
FILL FILL_1_OAI21X1_1711 ( );
FILL FILL_0_OAI21X1_1710 ( );
FILL FILL_1_OAI21X1_1710 ( );
FILL FILL_2_OAI21X1_1710 ( );
FILL FILL_0_BUFX4_34 ( );
FILL FILL_1_BUFX4_34 ( );
FILL FILL_0_OAI21X1_97 ( );
FILL FILL_1_OAI21X1_97 ( );
FILL FILL_2_OAI21X1_97 ( );
FILL FILL_0_OAI21X1_96 ( );
FILL FILL_1_OAI21X1_96 ( );
FILL FILL_0_DFFPOSX1_112 ( );
FILL FILL_1_DFFPOSX1_112 ( );
FILL FILL_2_DFFPOSX1_112 ( );
FILL FILL_3_DFFPOSX1_112 ( );
FILL FILL_4_DFFPOSX1_112 ( );
FILL FILL_5_DFFPOSX1_112 ( );
FILL FILL_0_OAI21X1_1786 ( );
FILL FILL_1_OAI21X1_1786 ( );
FILL FILL_0_NAND2X1_727 ( );
FILL FILL_0_BUFX2_649 ( );
FILL FILL_0_BUFX2_781 ( );
FILL FILL_0_BUFX2_809 ( );
FILL FILL_1_BUFX2_809 ( );
FILL FILL_0_NAND2X1_466 ( );
FILL FILL_1_NAND2X1_466 ( );
FILL FILL_0_DFFPOSX1_330 ( );
FILL FILL_1_DFFPOSX1_330 ( );
FILL FILL_2_DFFPOSX1_330 ( );
FILL FILL_3_DFFPOSX1_330 ( );
FILL FILL_4_DFFPOSX1_330 ( );
FILL FILL_5_DFFPOSX1_330 ( );
FILL FILL_6_DFFPOSX1_330 ( );
FILL FILL_0_OAI21X1_277 ( );
FILL FILL_1_OAI21X1_277 ( );
FILL FILL_0_OAI21X1_276 ( );
FILL FILL_1_OAI21X1_276 ( );
FILL FILL_0_BUFX2_65 ( );
FILL FILL_1_BUFX2_65 ( );
FILL FILL_0_BUFX2_937 ( );
FILL FILL_0_INVX2_117 ( );
FILL FILL_0_OAI21X1_1763 ( );
FILL FILL_1_OAI21X1_1763 ( );
FILL FILL_0_OAI21X1_1762 ( );
FILL FILL_1_OAI21X1_1762 ( );
FILL FILL_2_OAI21X1_1762 ( );
FILL FILL_0_DFFPOSX1_94 ( );
FILL FILL_1_DFFPOSX1_94 ( );
FILL FILL_2_DFFPOSX1_94 ( );
FILL FILL_3_DFFPOSX1_94 ( );
FILL FILL_4_DFFPOSX1_94 ( );
FILL FILL_5_DFFPOSX1_94 ( );
FILL FILL_6_DFFPOSX1_94 ( );
FILL FILL_0_BUFX2_1 ( );
FILL FILL_0_BUFX2_651 ( );
FILL FILL_0_BUFX2_764 ( );
FILL FILL_1_BUFX2_764 ( );
FILL FILL_0_OAI21X1_968 ( );
FILL FILL_1_OAI21X1_968 ( );
FILL FILL_0_OAI21X1_969 ( );
FILL FILL_1_OAI21X1_969 ( );
FILL FILL_0_DFFPOSX1_710 ( );
FILL FILL_1_DFFPOSX1_710 ( );
FILL FILL_2_DFFPOSX1_710 ( );
FILL FILL_3_DFFPOSX1_710 ( );
FILL FILL_4_DFFPOSX1_710 ( );
FILL FILL_5_DFFPOSX1_710 ( );
FILL FILL_0_BUFX2_700 ( );
FILL FILL_1_BUFX2_700 ( );
FILL FILL_0_NAND2X1_383 ( );
FILL FILL_0_BUFX2_845 ( );
FILL FILL_1_BUFX2_845 ( );
FILL FILL_0_INVX1_68 ( );
FILL FILL_0_OAI21X1_867 ( );
FILL FILL_1_OAI21X1_867 ( );
FILL FILL_0_DFFPOSX1_639 ( );
FILL FILL_1_DFFPOSX1_639 ( );
FILL FILL_2_DFFPOSX1_639 ( );
FILL FILL_3_DFFPOSX1_639 ( );
FILL FILL_4_DFFPOSX1_639 ( );
FILL FILL_5_DFFPOSX1_639 ( );
FILL FILL_0_INVX1_127 ( );
FILL FILL_1_INVX1_127 ( );
FILL FILL_0_DFFPOSX1_645 ( );
FILL FILL_1_DFFPOSX1_645 ( );
FILL FILL_2_DFFPOSX1_645 ( );
FILL FILL_3_DFFPOSX1_645 ( );
FILL FILL_4_DFFPOSX1_645 ( );
FILL FILL_5_DFFPOSX1_645 ( );
FILL FILL_0_INVX1_74 ( );
FILL FILL_0_OAI21X1_873 ( );
FILL FILL_1_OAI21X1_873 ( );
FILL FILL_0_INVX1_85 ( );
FILL FILL_0_DFFPOSX1_694 ( );
FILL FILL_1_DFFPOSX1_694 ( );
FILL FILL_2_DFFPOSX1_694 ( );
FILL FILL_3_DFFPOSX1_694 ( );
FILL FILL_4_DFFPOSX1_694 ( );
FILL FILL_5_DFFPOSX1_694 ( );
FILL FILL_6_DFFPOSX1_694 ( );
FILL FILL_0_OAI21X1_937 ( );
FILL FILL_1_OAI21X1_937 ( );
FILL FILL_0_INVX2_200 ( );
FILL FILL_0_BUFX2_868 ( );
FILL FILL_1_BUFX2_868 ( );
FILL FILL_0_OAI21X1_936 ( );
FILL FILL_1_OAI21X1_936 ( );
FILL FILL_0_BUFX2_996 ( );
FILL FILL_1_BUFX2_996 ( );
FILL FILL_0_BUFX2_955 ( );
FILL FILL_1_BUFX2_955 ( );
FILL FILL_0_INVX2_167 ( );
FILL FILL_0_OAI21X1_1807 ( );
FILL FILL_1_OAI21X1_1807 ( );
FILL FILL_0_NAND2X1_748 ( );
FILL FILL_1_NAND2X1_748 ( );
FILL FILL_0_DFFPOSX1_133 ( );
FILL FILL_1_DFFPOSX1_133 ( );
FILL FILL_2_DFFPOSX1_133 ( );
FILL FILL_3_DFFPOSX1_133 ( );
FILL FILL_4_DFFPOSX1_133 ( );
FILL FILL_5_DFFPOSX1_133 ( );
FILL FILL_6_DFFPOSX1_133 ( );
FILL FILL_0_OAI21X1_890 ( );
FILL FILL_1_OAI21X1_890 ( );
FILL FILL_0_DFFPOSX1_662 ( );
FILL FILL_1_DFFPOSX1_662 ( );
FILL FILL_2_DFFPOSX1_662 ( );
FILL FILL_3_DFFPOSX1_662 ( );
FILL FILL_4_DFFPOSX1_662 ( );
FILL FILL_5_DFFPOSX1_662 ( );
FILL FILL_0_INVX1_109 ( );
FILL FILL_0_BUFX4_197 ( );
FILL FILL_1_BUFX4_197 ( );
FILL FILL_0_BUFX2_753 ( );
FILL FILL_0_DFFPOSX1_168 ( );
FILL FILL_1_DFFPOSX1_168 ( );
FILL FILL_2_DFFPOSX1_168 ( );
FILL FILL_3_DFFPOSX1_168 ( );
FILL FILL_4_DFFPOSX1_168 ( );
FILL FILL_5_DFFPOSX1_168 ( );
FILL FILL_0_BUFX4_216 ( );
FILL FILL_1_BUFX4_216 ( );
FILL FILL_0_DFFPOSX1_32 ( );
FILL FILL_1_DFFPOSX1_32 ( );
FILL FILL_2_DFFPOSX1_32 ( );
FILL FILL_3_DFFPOSX1_32 ( );
FILL FILL_4_DFFPOSX1_32 ( );
FILL FILL_5_DFFPOSX1_32 ( );
FILL FILL_0_DFFPOSX1_812 ( );
FILL FILL_1_DFFPOSX1_812 ( );
FILL FILL_2_DFFPOSX1_812 ( );
FILL FILL_3_DFFPOSX1_812 ( );
FILL FILL_4_DFFPOSX1_812 ( );
FILL FILL_5_DFFPOSX1_812 ( );
FILL FILL_0_OAI21X1_1106 ( );
FILL FILL_1_OAI21X1_1106 ( );
FILL FILL_0_BUFX2_191 ( );
FILL FILL_0_DFFPOSX1_746 ( );
FILL FILL_1_DFFPOSX1_746 ( );
FILL FILL_2_DFFPOSX1_746 ( );
FILL FILL_3_DFFPOSX1_746 ( );
FILL FILL_4_DFFPOSX1_746 ( );
FILL FILL_5_DFFPOSX1_746 ( );
FILL FILL_6_DFFPOSX1_746 ( );
FILL FILL_0_NAND2X1_404 ( );
FILL FILL_1_NAND2X1_404 ( );
FILL FILL_0_OAI21X1_1038 ( );
FILL FILL_1_OAI21X1_1038 ( );
FILL FILL_0_BUFX2_127 ( );
FILL FILL_1_BUFX2_127 ( );
FILL FILL_0_NAND2X1_409 ( );
FILL FILL_0_DFFPOSX1_814 ( );
FILL FILL_1_DFFPOSX1_814 ( );
FILL FILL_2_DFFPOSX1_814 ( );
FILL FILL_3_DFFPOSX1_814 ( );
FILL FILL_4_DFFPOSX1_814 ( );
FILL FILL_5_DFFPOSX1_814 ( );
FILL FILL_0_BUFX2_575 ( );
FILL FILL_1_BUFX2_575 ( );
FILL FILL_0_DFFPOSX1_119 ( );
FILL FILL_1_DFFPOSX1_119 ( );
FILL FILL_2_DFFPOSX1_119 ( );
FILL FILL_3_DFFPOSX1_119 ( );
FILL FILL_4_DFFPOSX1_119 ( );
FILL FILL_5_DFFPOSX1_119 ( );
FILL FILL_0_OAI21X1_1793 ( );
FILL FILL_1_OAI21X1_1793 ( );
FILL FILL_0_BUFX2_576 ( );
FILL FILL_0_OAI21X1_1213 ( );
FILL FILL_1_OAI21X1_1213 ( );
FILL FILL_0_OAI21X1_1212 ( );
FILL FILL_1_OAI21X1_1212 ( );
FILL FILL_0_BUFX2_746 ( );
FILL FILL_1_BUFX2_746 ( );
FILL FILL_0_DFFPOSX1_232 ( );
FILL FILL_1_DFFPOSX1_232 ( );
FILL FILL_2_DFFPOSX1_232 ( );
FILL FILL_3_DFFPOSX1_232 ( );
FILL FILL_4_DFFPOSX1_232 ( );
FILL FILL_5_DFFPOSX1_232 ( );
FILL FILL_6_DFFPOSX1_232 ( );
FILL FILL_0_OAI21X1_1713 ( );
FILL FILL_1_OAI21X1_1713 ( );
FILL FILL_0_INVX2_155 ( );
FILL FILL_0_BUFX2_579 ( );
FILL FILL_0_DFFPOSX1_414 ( );
FILL FILL_1_DFFPOSX1_414 ( );
FILL FILL_2_DFFPOSX1_414 ( );
FILL FILL_3_DFFPOSX1_414 ( );
FILL FILL_4_DFFPOSX1_414 ( );
FILL FILL_5_DFFPOSX1_414 ( );
FILL FILL_6_DFFPOSX1_414 ( );
FILL FILL_0_DFFPOSX1_262 ( );
FILL FILL_1_DFFPOSX1_262 ( );
FILL FILL_2_DFFPOSX1_262 ( );
FILL FILL_3_DFFPOSX1_262 ( );
FILL FILL_4_DFFPOSX1_262 ( );
FILL FILL_5_DFFPOSX1_262 ( );
FILL FILL_0_DFFPOSX1_145 ( );
FILL FILL_1_DFFPOSX1_145 ( );
FILL FILL_2_DFFPOSX1_145 ( );
FILL FILL_3_DFFPOSX1_145 ( );
FILL FILL_4_DFFPOSX1_145 ( );
FILL FILL_5_DFFPOSX1_145 ( );
FILL FILL_0_OAI21X1_387 ( );
FILL FILL_1_OAI21X1_387 ( );
FILL FILL_0_NAND2X1_131 ( );
FILL FILL_1_NAND2X1_131 ( );
FILL FILL_0_BUFX2_580 ( );
FILL FILL_1_BUFX2_580 ( );
FILL FILL_0_BUFX2_516 ( );
FILL FILL_0_DFFPOSX1_37 ( );
FILL FILL_1_DFFPOSX1_37 ( );
FILL FILL_2_DFFPOSX1_37 ( );
FILL FILL_3_DFFPOSX1_37 ( );
FILL FILL_4_DFFPOSX1_37 ( );
FILL FILL_5_DFFPOSX1_37 ( );
FILL FILL_6_DFFPOSX1_37 ( );
FILL FILL_0_BUFX2_138 ( );
FILL FILL_1_BUFX2_138 ( );
FILL FILL_0_DFFPOSX1_237 ( );
FILL FILL_1_DFFPOSX1_237 ( );
FILL FILL_2_DFFPOSX1_237 ( );
FILL FILL_3_DFFPOSX1_237 ( );
FILL FILL_4_DFFPOSX1_237 ( );
FILL FILL_5_DFFPOSX1_237 ( );
FILL FILL_6_DFFPOSX1_237 ( );
FILL FILL_0_DFFPOSX1_309 ( );
FILL FILL_1_DFFPOSX1_309 ( );
FILL FILL_2_DFFPOSX1_309 ( );
FILL FILL_3_DFFPOSX1_309 ( );
FILL FILL_4_DFFPOSX1_309 ( );
FILL FILL_5_DFFPOSX1_309 ( );
FILL FILL_0_OAI21X1_235 ( );
FILL FILL_1_OAI21X1_235 ( );
FILL FILL_0_OAI21X1_1791 ( );
FILL FILL_1_OAI21X1_1791 ( );
FILL FILL_2_OAI21X1_1791 ( );
FILL FILL_0_NAND2X1_732 ( );
FILL FILL_0_NAND2X1_719 ( );
FILL FILL_0_DFFPOSX1_104 ( );
FILL FILL_1_DFFPOSX1_104 ( );
FILL FILL_2_DFFPOSX1_104 ( );
FILL FILL_3_DFFPOSX1_104 ( );
FILL FILL_4_DFFPOSX1_104 ( );
FILL FILL_5_DFFPOSX1_104 ( );
FILL FILL_6_DFFPOSX1_104 ( );
FILL FILL_0_BUFX2_951 ( );
FILL FILL_1_BUFX2_951 ( );
FILL FILL_0_OAI21X1_1029 ( );
FILL FILL_1_OAI21X1_1029 ( );
FILL FILL_0_OAI21X1_209 ( );
FILL FILL_1_OAI21X1_209 ( );
FILL FILL_0_OAI21X1_208 ( );
FILL FILL_1_OAI21X1_208 ( );
FILL FILL_0_OAI21X1_1028 ( );
FILL FILL_1_OAI21X1_1028 ( );
FILL FILL_0_BUFX2_865 ( );
FILL FILL_0_INVX2_146 ( );
FILL FILL_0_DFFPOSX1_337 ( );
FILL FILL_1_DFFPOSX1_337 ( );
FILL FILL_2_DFFPOSX1_337 ( );
FILL FILL_3_DFFPOSX1_337 ( );
FILL FILL_4_DFFPOSX1_337 ( );
FILL FILL_5_DFFPOSX1_337 ( );
FILL FILL_0_OAI21X1_290 ( );
FILL FILL_1_OAI21X1_290 ( );
FILL FILL_0_DFFPOSX1_322 ( );
FILL FILL_1_DFFPOSX1_322 ( );
FILL FILL_2_DFFPOSX1_322 ( );
FILL FILL_3_DFFPOSX1_322 ( );
FILL FILL_4_DFFPOSX1_322 ( );
FILL FILL_5_DFFPOSX1_322 ( );
FILL FILL_0_OAI21X1_261 ( );
FILL FILL_1_OAI21X1_261 ( );
FILL FILL_0_OAI21X1_260 ( );
FILL FILL_1_OAI21X1_260 ( );
FILL FILL_0_DFFPOSX1_316 ( );
FILL FILL_1_DFFPOSX1_316 ( );
FILL FILL_2_DFFPOSX1_316 ( );
FILL FILL_3_DFFPOSX1_316 ( );
FILL FILL_4_DFFPOSX1_316 ( );
FILL FILL_5_DFFPOSX1_316 ( );
FILL FILL_0_NAND2X1_1 ( );
FILL FILL_0_DFFPOSX1_285 ( );
FILL FILL_1_DFFPOSX1_285 ( );
FILL FILL_2_DFFPOSX1_285 ( );
FILL FILL_3_DFFPOSX1_285 ( );
FILL FILL_4_DFFPOSX1_285 ( );
FILL FILL_5_DFFPOSX1_285 ( );
FILL FILL_0_BUFX2_362 ( );
FILL FILL_1_BUFX2_362 ( );
FILL FILL_0_INVX2_162 ( );
FILL FILL_0_OAI21X1_1830 ( );
FILL FILL_1_OAI21X1_1830 ( );
FILL FILL_2_OAI21X1_1830 ( );
FILL FILL_0_NAND2X1_771 ( );
FILL FILL_0_DFFPOSX1_188 ( );
FILL FILL_1_DFFPOSX1_188 ( );
FILL FILL_2_DFFPOSX1_188 ( );
FILL FILL_3_DFFPOSX1_188 ( );
FILL FILL_4_DFFPOSX1_188 ( );
FILL FILL_5_DFFPOSX1_188 ( );
FILL FILL_0_BUFX2_947 ( );
FILL FILL_1_BUFX2_947 ( );
FILL FILL_0_BUFX2_922 ( );
FILL FILL_0_BUFX4_207 ( );
FILL FILL_1_BUFX4_207 ( );
FILL FILL_0_DFFPOSX1_1011 ( );
FILL FILL_1_DFFPOSX1_1011 ( );
FILL FILL_2_DFFPOSX1_1011 ( );
FILL FILL_3_DFFPOSX1_1011 ( );
FILL FILL_4_DFFPOSX1_1011 ( );
FILL FILL_5_DFFPOSX1_1011 ( );
FILL FILL_0_BUFX2_742 ( );
FILL FILL_0_DFFPOSX1_211 ( );
FILL FILL_1_DFFPOSX1_211 ( );
FILL FILL_2_DFFPOSX1_211 ( );
FILL FILL_3_DFFPOSX1_211 ( );
FILL FILL_4_DFFPOSX1_211 ( );
FILL FILL_5_DFFPOSX1_211 ( );
FILL FILL_6_DFFPOSX1_211 ( );
FILL FILL_0_INVX1_154 ( );
FILL FILL_0_DFFPOSX1_208 ( );
FILL FILL_1_DFFPOSX1_208 ( );
FILL FILL_2_DFFPOSX1_208 ( );
FILL FILL_3_DFFPOSX1_208 ( );
FILL FILL_4_DFFPOSX1_208 ( );
FILL FILL_5_DFFPOSX1_208 ( );
FILL FILL_6_DFFPOSX1_208 ( );
FILL FILL_0_INVX2_176 ( );
FILL FILL_0_NAND2X1_740 ( );
FILL FILL_0_OAI21X1_1799 ( );
FILL FILL_1_OAI21X1_1799 ( );
FILL FILL_0_OAI21X1_1800 ( );
FILL FILL_1_OAI21X1_1800 ( );
FILL FILL_0_NAND2X1_741 ( );
FILL FILL_1_NAND2X1_741 ( );
FILL FILL_0_BUFX2_816 ( );
FILL FILL_1_BUFX2_816 ( );
FILL FILL_0_OAI21X1_1785 ( );
FILL FILL_1_OAI21X1_1785 ( );
FILL FILL_0_NAND2X1_726 ( );
FILL FILL_0_OAI21X1_19 ( );
FILL FILL_1_OAI21X1_19 ( );
FILL FILL_2_OAI21X1_19 ( );
FILL FILL_0_NAND2X1_19 ( );
FILL FILL_0_DFFPOSX1_670 ( );
FILL FILL_1_DFFPOSX1_670 ( );
FILL FILL_2_DFFPOSX1_670 ( );
FILL FILL_3_DFFPOSX1_670 ( );
FILL FILL_4_DFFPOSX1_670 ( );
FILL FILL_5_DFFPOSX1_670 ( );
FILL FILL_6_DFFPOSX1_670 ( );
FILL FILL_0_NAND2X1_699 ( );
FILL FILL_1_NAND2X1_699 ( );
FILL FILL_0_INVX2_171 ( );
FILL FILL_1_INVX2_171 ( );
FILL FILL_0_OAI21X1_1631 ( );
FILL FILL_1_OAI21X1_1631 ( );
FILL FILL_0_NAND2X1_768 ( );
FILL FILL_1_NAND2X1_768 ( );
FILL FILL_0_OAI21X1_1827 ( );
FILL FILL_1_OAI21X1_1827 ( );
FILL FILL_0_OAI21X1_1590 ( );
FILL FILL_1_OAI21X1_1590 ( );
FILL FILL_0_NAND2X1_659 ( );
FILL FILL_0_BUFX2_1018 ( );
FILL FILL_0_BUFX2_658 ( );
FILL FILL_1_BUFX2_658 ( );
FILL FILL_0_BUFX2_217 ( );
FILL FILL_0_OAI21X1_1629 ( );
FILL FILL_1_OAI21X1_1629 ( );
FILL FILL_0_BUFX2_92 ( );
FILL FILL_0_OAI21X1_1596 ( );
FILL FILL_1_OAI21X1_1596 ( );
FILL FILL_0_NAND2X1_665 ( );
FILL FILL_1_NAND2X1_665 ( );
FILL FILL_0_BUFX4_11 ( );
FILL FILL_1_BUFX4_11 ( );
FILL FILL_0_DFFPOSX1_198 ( );
FILL FILL_1_DFFPOSX1_198 ( );
FILL FILL_2_DFFPOSX1_198 ( );
FILL FILL_3_DFFPOSX1_198 ( );
FILL FILL_4_DFFPOSX1_198 ( );
FILL FILL_5_DFFPOSX1_198 ( );
FILL FILL_6_DFFPOSX1_198 ( );
FILL FILL_0_OAI21X1_42 ( );
FILL FILL_1_OAI21X1_42 ( );
FILL FILL_0_NAND2X1_42 ( );
FILL FILL_0_INVX2_132 ( );
FILL FILL_0_DFFPOSX1_242 ( );
FILL FILL_1_DFFPOSX1_242 ( );
FILL FILL_2_DFFPOSX1_242 ( );
FILL FILL_3_DFFPOSX1_242 ( );
FILL FILL_4_DFFPOSX1_242 ( );
FILL FILL_5_DFFPOSX1_242 ( );
FILL FILL_0_OAI21X1_1674 ( );
FILL FILL_1_OAI21X1_1674 ( );
FILL FILL_0_BUFX2_997 ( );
FILL FILL_0_INVX1_171 ( );
FILL FILL_0_BUFX2_719 ( );
FILL FILL_0_DFFPOSX1_304 ( );
FILL FILL_1_DFFPOSX1_304 ( );
FILL FILL_2_DFFPOSX1_304 ( );
FILL FILL_3_DFFPOSX1_304 ( );
FILL FILL_4_DFFPOSX1_304 ( );
FILL FILL_5_DFFPOSX1_304 ( );
FILL FILL_6_DFFPOSX1_304 ( );
FILL FILL_0_OAI21X1_225 ( );
FILL FILL_1_OAI21X1_225 ( );
FILL FILL_0_OAI21X1_224 ( );
FILL FILL_1_OAI21X1_224 ( );
FILL FILL_0_DFFPOSX1_319 ( );
FILL FILL_1_DFFPOSX1_319 ( );
FILL FILL_2_DFFPOSX1_319 ( );
FILL FILL_3_DFFPOSX1_319 ( );
FILL FILL_4_DFFPOSX1_319 ( );
FILL FILL_5_DFFPOSX1_319 ( );
FILL FILL_6_DFFPOSX1_319 ( );
FILL FILL_0_BUFX2_973 ( );
FILL FILL_1_BUFX2_973 ( );
FILL FILL_0_OAI21X1_35 ( );
FILL FILL_1_OAI21X1_35 ( );
FILL FILL_0_NAND2X1_35 ( );
FILL FILL_1_NAND2X1_35 ( );
FILL FILL_0_INVX2_131 ( );
FILL FILL_0_DFFPOSX1_718 ( );
FILL FILL_1_DFFPOSX1_718 ( );
FILL FILL_2_DFFPOSX1_718 ( );
FILL FILL_3_DFFPOSX1_718 ( );
FILL FILL_4_DFFPOSX1_718 ( );
FILL FILL_5_DFFPOSX1_718 ( );
FILL FILL_6_DFFPOSX1_718 ( );
FILL FILL_0_OAI21X1_1727 ( );
FILL FILL_1_OAI21X1_1727 ( );
FILL FILL_0_DFFPOSX1_76 ( );
FILL FILL_1_DFFPOSX1_76 ( );
FILL FILL_2_DFFPOSX1_76 ( );
FILL FILL_3_DFFPOSX1_76 ( );
FILL FILL_4_DFFPOSX1_76 ( );
FILL FILL_5_DFFPOSX1_76 ( );
FILL FILL_6_DFFPOSX1_76 ( );
FILL FILL_0_BUFX2_1001 ( );
FILL FILL_1_BUFX2_1001 ( );
FILL FILL_0_DFFPOSX1_59 ( );
FILL FILL_1_DFFPOSX1_59 ( );
FILL FILL_2_DFFPOSX1_59 ( );
FILL FILL_3_DFFPOSX1_59 ( );
FILL FILL_4_DFFPOSX1_59 ( );
FILL FILL_5_DFFPOSX1_59 ( );
FILL FILL_6_DFFPOSX1_59 ( );
FILL FILL_0_OAI21X1_1693 ( );
FILL FILL_1_OAI21X1_1693 ( );
FILL FILL_0_OAI21X1_1692 ( );
FILL FILL_1_OAI21X1_1692 ( );
FILL FILL_2_OAI21X1_1692 ( );
FILL FILL_0_INVX2_143 ( );
FILL FILL_1_INVX2_143 ( );
FILL FILL_0_OAI21X1_126 ( );
FILL FILL_1_OAI21X1_126 ( );
FILL FILL_0_OAI21X1_127 ( );
FILL FILL_1_OAI21X1_127 ( );
FILL FILL_0_DFFPOSX1_255 ( );
FILL FILL_1_DFFPOSX1_255 ( );
FILL FILL_2_DFFPOSX1_255 ( );
FILL FILL_3_DFFPOSX1_255 ( );
FILL FILL_4_DFFPOSX1_255 ( );
FILL FILL_5_DFFPOSX1_255 ( );
FILL FILL_0_BUFX2_278 ( );
FILL FILL_1_BUFX2_278 ( );
FILL FILL_0_NAND2X1_373 ( );
FILL FILL_1_NAND2X1_373 ( );
FILL FILL_0_NAND2X1_375 ( );
FILL FILL_0_INVX1_139 ( );
FILL FILL_0_BUFX2_277 ( );
FILL FILL_0_NAND2X1_361 ( );
FILL FILL_1_NAND2X1_361 ( );
FILL FILL_0_NAND2X1_358 ( );
FILL FILL_1_NAND2X1_358 ( );
FILL FILL_0_BUFX2_301 ( );
FILL FILL_1_BUFX2_301 ( );
FILL FILL_0_DFFPOSX1_664 ( );
FILL FILL_1_DFFPOSX1_664 ( );
FILL FILL_2_DFFPOSX1_664 ( );
FILL FILL_3_DFFPOSX1_664 ( );
FILL FILL_4_DFFPOSX1_664 ( );
FILL FILL_5_DFFPOSX1_664 ( );
FILL FILL_0_OAI21X1_892 ( );
FILL FILL_1_OAI21X1_892 ( );
FILL FILL_0_NAND2X1_386 ( );
FILL FILL_1_NAND2X1_386 ( );
FILL FILL_0_BUFX2_283 ( );
FILL FILL_1_BUFX2_283 ( );
FILL FILL_0_NAND2X1_367 ( );
FILL FILL_1_NAND2X1_367 ( );
FILL FILL_0_BUFX2_348 ( );
FILL FILL_1_BUFX2_348 ( );
FILL FILL_0_BUFX2_331 ( );
FILL FILL_1_BUFX2_331 ( );
FILL FILL_0_DFFPOSX1_683 ( );
FILL FILL_1_DFFPOSX1_683 ( );
FILL FILL_2_DFFPOSX1_683 ( );
FILL FILL_3_DFFPOSX1_683 ( );
FILL FILL_4_DFFPOSX1_683 ( );
FILL FILL_5_DFFPOSX1_683 ( );
FILL FILL_6_DFFPOSX1_683 ( );
FILL FILL_0_OAI21X1_915 ( );
FILL FILL_1_OAI21X1_915 ( );
FILL FILL_0_OAI21X1_914 ( );
FILL FILL_1_OAI21X1_914 ( );
FILL FILL_0_OAI21X1_929 ( );
FILL FILL_1_OAI21X1_929 ( );
FILL FILL_0_OAI21X1_928 ( );
FILL FILL_1_OAI21X1_928 ( );
FILL FILL_2_OAI21X1_928 ( );
FILL FILL_0_OAI21X1_956 ( );
FILL FILL_1_OAI21X1_956 ( );
FILL FILL_0_BUFX2_804 ( );
FILL FILL_1_BUFX2_804 ( );
FILL FILL_0_DFFPOSX1_690 ( );
FILL FILL_1_DFFPOSX1_690 ( );
FILL FILL_2_DFFPOSX1_690 ( );
FILL FILL_3_DFFPOSX1_690 ( );
FILL FILL_4_DFFPOSX1_690 ( );
FILL FILL_5_DFFPOSX1_690 ( );
FILL FILL_0_OAI21X1_139 ( );
FILL FILL_1_OAI21X1_139 ( );
FILL FILL_0_OAI21X1_138 ( );
FILL FILL_1_OAI21X1_138 ( );
FILL FILL_0_NAND2X1_384 ( );
FILL FILL_1_NAND2X1_384 ( );
FILL FILL_0_BUFX2_299 ( );
FILL FILL_1_BUFX2_299 ( );
FILL FILL_0_BUFX2_670 ( );
FILL FILL_0_DFFPOSX1_261 ( );
FILL FILL_1_DFFPOSX1_261 ( );
FILL FILL_2_DFFPOSX1_261 ( );
FILL FILL_3_DFFPOSX1_261 ( );
FILL FILL_4_DFFPOSX1_261 ( );
FILL FILL_5_DFFPOSX1_261 ( );
FILL FILL_0_DFFPOSX1_672 ( );
FILL FILL_1_DFFPOSX1_672 ( );
FILL FILL_2_DFFPOSX1_672 ( );
FILL FILL_3_DFFPOSX1_672 ( );
FILL FILL_4_DFFPOSX1_672 ( );
FILL FILL_5_DFFPOSX1_672 ( );
FILL FILL_6_DFFPOSX1_672 ( );
FILL FILL_0_BUFX2_238 ( );
FILL FILL_0_BUFX2_163 ( );
FILL FILL_0_NAND2X1_12 ( );
FILL FILL_1_NAND2X1_12 ( );
FILL FILL_0_OAI21X1_12 ( );
FILL FILL_1_OAI21X1_12 ( );
FILL FILL_0_OAI21X1_1642 ( );
FILL FILL_1_OAI21X1_1642 ( );
FILL FILL_0_NAND2X1_710 ( );
FILL FILL_1_NAND2X1_710 ( );
FILL FILL_0_NAND2X1_471 ( );
FILL FILL_1_NAND2X1_471 ( );
FILL FILL_0_DFFPOSX1_815 ( );
FILL FILL_1_DFFPOSX1_815 ( );
FILL FILL_2_DFFPOSX1_815 ( );
FILL FILL_3_DFFPOSX1_815 ( );
FILL FILL_4_DFFPOSX1_815 ( );
FILL FILL_5_DFFPOSX1_815 ( );
FILL FILL_6_DFFPOSX1_815 ( );
FILL FILL_0_OAI21X1_1114 ( );
FILL FILL_1_OAI21X1_1114 ( );
FILL FILL_0_NAND2X1_478 ( );
FILL FILL_1_NAND2X1_478 ( );
FILL FILL_0_OAI21X1_23 ( );
FILL FILL_1_OAI21X1_23 ( );
FILL FILL_0_BUFX2_64 ( );
FILL FILL_0_DFFPOSX1_179 ( );
FILL FILL_1_DFFPOSX1_179 ( );
FILL FILL_2_DFFPOSX1_179 ( );
FILL FILL_3_DFFPOSX1_179 ( );
FILL FILL_4_DFFPOSX1_179 ( );
FILL FILL_5_DFFPOSX1_179 ( );
FILL FILL_0_BUFX2_121 ( );
FILL FILL_0_NAND2X1_475 ( );
FILL FILL_0_BUFX2_912 ( );
FILL FILL_1_BUFX2_912 ( );
FILL FILL_0_DFFPOSX1_751 ( );
FILL FILL_1_DFFPOSX1_751 ( );
FILL FILL_2_DFFPOSX1_751 ( );
FILL FILL_3_DFFPOSX1_751 ( );
FILL FILL_4_DFFPOSX1_751 ( );
FILL FILL_5_DFFPOSX1_751 ( );
FILL FILL_0_BUFX2_788 ( );
FILL FILL_1_BUFX2_788 ( );
FILL FILL_0_NAND2X1_734 ( );
FILL FILL_1_NAND2X1_734 ( );
FILL FILL_0_BUFX2_192 ( );
FILL FILL_1_BUFX2_192 ( );
FILL FILL_0_DFFPOSX1_874 ( );
FILL FILL_1_DFFPOSX1_874 ( );
FILL FILL_2_DFFPOSX1_874 ( );
FILL FILL_3_DFFPOSX1_874 ( );
FILL FILL_4_DFFPOSX1_874 ( );
FILL FILL_5_DFFPOSX1_874 ( );
FILL FILL_6_DFFPOSX1_874 ( );
FILL FILL_0_OAI21X1_106 ( );
FILL FILL_1_OAI21X1_106 ( );
FILL FILL_0_OAI21X1_107 ( );
FILL FILL_1_OAI21X1_107 ( );
FILL FILL_0_BUFX2_489 ( );
FILL FILL_1_BUFX2_489 ( );
FILL FILL_0_OAI21X1_81 ( );
FILL FILL_1_OAI21X1_81 ( );
FILL FILL_0_BUFX2_197 ( );
FILL FILL_1_BUFX2_197 ( );
FILL FILL_0_OAI21X1_80 ( );
FILL FILL_1_OAI21X1_80 ( );
FILL FILL_0_BUFX2_447 ( );
FILL FILL_1_BUFX2_447 ( );
FILL FILL_0_BUFX2_689 ( );
FILL FILL_1_BUFX2_689 ( );
FILL FILL_0_BUFX2_657 ( );
FILL FILL_0_NAND2X1_666 ( );
FILL FILL_1_NAND2X1_666 ( );
FILL FILL_0_OAI21X1_1597 ( );
FILL FILL_1_OAI21X1_1597 ( );
FILL FILL_0_BUFX2_933 ( );
FILL FILL_1_BUFX2_933 ( );
FILL FILL_0_BUFX2_817 ( );
FILL FILL_1_BUFX2_817 ( );
FILL FILL_0_BUFX2_5 ( );
FILL FILL_1_BUFX2_5 ( );
FILL FILL_0_DFFPOSX1_1020 ( );
FILL FILL_1_DFFPOSX1_1020 ( );
FILL FILL_2_DFFPOSX1_1020 ( );
FILL FILL_3_DFFPOSX1_1020 ( );
FILL FILL_4_DFFPOSX1_1020 ( );
FILL FILL_5_DFFPOSX1_1020 ( );
FILL FILL_0_NAND2X1_760 ( );
FILL FILL_1_NAND2X1_760 ( );
FILL FILL_0_OAI21X1_1819 ( );
FILL FILL_1_OAI21X1_1819 ( );
FILL FILL_0_DFFPOSX1_415 ( );
FILL FILL_1_DFFPOSX1_415 ( );
FILL FILL_2_DFFPOSX1_415 ( );
FILL FILL_3_DFFPOSX1_415 ( );
FILL FILL_4_DFFPOSX1_415 ( );
FILL FILL_5_DFFPOSX1_415 ( );
FILL FILL_0_BUFX2_714 ( );
FILL FILL_0_BUFX2_196 ( );
FILL FILL_0_OAI21X1_1648 ( );
FILL FILL_1_OAI21X1_1648 ( );
FILL FILL_0_BUFX2_4 ( );
FILL FILL_0_OAI21X1_1649 ( );
FILL FILL_1_OAI21X1_1649 ( );
FILL FILL_0_BUFX2_71 ( );
FILL FILL_1_BUFX2_71 ( );
FILL FILL_0_BUFX2_968 ( );
FILL FILL_1_BUFX2_968 ( );
FILL FILL_0_BUFX2_136 ( );
FILL FILL_1_BUFX2_136 ( );
FILL FILL_0_OAI21X1_1126 ( );
FILL FILL_1_OAI21X1_1126 ( );
FILL FILL_0_DFFPOSX1_5 ( );
FILL FILL_1_DFFPOSX1_5 ( );
FILL FILL_2_DFFPOSX1_5 ( );
FILL FILL_3_DFFPOSX1_5 ( );
FILL FILL_4_DFFPOSX1_5 ( );
FILL FILL_5_DFFPOSX1_5 ( );
FILL FILL_6_DFFPOSX1_5 ( );
FILL FILL_0_OAI21X1_1778 ( );
FILL FILL_1_OAI21X1_1778 ( );
FILL FILL_2_OAI21X1_1778 ( );
FILL FILL_0_DFFPOSX1_117 ( );
FILL FILL_1_DFFPOSX1_117 ( );
FILL FILL_2_DFFPOSX1_117 ( );
FILL FILL_3_DFFPOSX1_117 ( );
FILL FILL_4_DFFPOSX1_117 ( );
FILL FILL_5_DFFPOSX1_117 ( );
FILL FILL_6_DFFPOSX1_117 ( );
FILL FILL_0_DFFPOSX1_296 ( );
FILL FILL_1_DFFPOSX1_296 ( );
FILL FILL_2_DFFPOSX1_296 ( );
FILL FILL_3_DFFPOSX1_296 ( );
FILL FILL_4_DFFPOSX1_296 ( );
FILL FILL_5_DFFPOSX1_296 ( );
FILL FILL_0_BUFX2_202 ( );
FILL FILL_0_OAI21X1_979 ( );
FILL FILL_1_OAI21X1_979 ( );
FILL FILL_0_BUFX2_8 ( );
FILL FILL_1_BUFX2_8 ( );
FILL FILL_0_OAI21X1_978 ( );
FILL FILL_1_OAI21X1_978 ( );
FILL FILL_0_BUFX2_378 ( );
FILL FILL_0_OAI21X1_291 ( );
FILL FILL_1_OAI21X1_291 ( );
FILL FILL_0_OAI21X1_163 ( );
FILL FILL_1_OAI21X1_163 ( );
FILL FILL_0_OAI21X1_162 ( );
FILL FILL_1_OAI21X1_162 ( );
FILL FILL_2_OAI21X1_162 ( );
FILL FILL_0_BUFX2_1009 ( );
FILL FILL_1_BUFX2_1009 ( );
FILL FILL_0_BUFX2_201 ( );
FILL FILL_1_BUFX2_201 ( );
FILL FILL_0_BUFX2_929 ( );
FILL FILL_1_BUFX2_929 ( );
FILL FILL_0_OAI21X1_248 ( );
FILL FILL_1_OAI21X1_248 ( );
FILL FILL_0_BUFX2_137 ( );
FILL FILL_0_OAI21X1_249 ( );
FILL FILL_1_OAI21X1_249 ( );
FILL FILL_0_BUFX2_993 ( );
FILL FILL_1_BUFX2_993 ( );
FILL FILL_0_OAI21X1_1 ( );
FILL FILL_1_OAI21X1_1 ( );
FILL FILL_0_DFFPOSX1_157 ( );
FILL FILL_1_DFFPOSX1_157 ( );
FILL FILL_2_DFFPOSX1_157 ( );
FILL FILL_3_DFFPOSX1_157 ( );
FILL FILL_4_DFFPOSX1_157 ( );
FILL FILL_5_DFFPOSX1_157 ( );
FILL FILL_0_DFFPOSX1_156 ( );
FILL FILL_1_DFFPOSX1_156 ( );
FILL FILL_2_DFFPOSX1_156 ( );
FILL FILL_3_DFFPOSX1_156 ( );
FILL FILL_4_DFFPOSX1_156 ( );
FILL FILL_5_DFFPOSX1_156 ( );
FILL FILL_6_DFFPOSX1_156 ( );
FILL FILL_0_OAI21X1_32 ( );
FILL FILL_1_OAI21X1_32 ( );
FILL FILL_2_OAI21X1_32 ( );
FILL FILL_0_NAND2X1_32 ( );
FILL FILL_0_BUFX2_794 ( );
FILL FILL_0_BUFX2_858 ( );
FILL FILL_1_BUFX2_858 ( );
FILL FILL_0_OAI21X1_55 ( );
FILL FILL_1_OAI21X1_55 ( );
FILL FILL_0_NAND2X1_55 ( );
FILL FILL_0_BUFX2_678 ( );
FILL FILL_1_BUFX2_678 ( );
FILL FILL_0_BUFX2_883 ( );
FILL FILL_0_BUFX2_859 ( );
FILL FILL_0_BUFX2_88 ( );
FILL FILL_1_BUFX2_88 ( );
FILL FILL_0_NAND2X1_52 ( );
FILL FILL_1_NAND2X1_52 ( );
FILL FILL_0_OAI21X1_52 ( );
FILL FILL_1_OAI21X1_52 ( );
FILL FILL_0_BUFX2_944 ( );
FILL FILL_1_BUFX2_944 ( );
FILL FILL_0_DFFPOSX1_190 ( );
FILL FILL_1_DFFPOSX1_190 ( );
FILL FILL_2_DFFPOSX1_190 ( );
FILL FILL_3_DFFPOSX1_190 ( );
FILL FILL_4_DFFPOSX1_190 ( );
FILL FILL_5_DFFPOSX1_190 ( );
FILL FILL_0_NAND2X1_34 ( );
FILL FILL_1_NAND2X1_34 ( );
FILL FILL_0_OAI21X1_34 ( );
FILL FILL_1_OAI21X1_34 ( );
FILL FILL_0_DFFPOSX1_125 ( );
FILL FILL_1_DFFPOSX1_125 ( );
FILL FILL_2_DFFPOSX1_125 ( );
FILL FILL_3_DFFPOSX1_125 ( );
FILL FILL_4_DFFPOSX1_125 ( );
FILL FILL_5_DFFPOSX1_125 ( );
FILL FILL_0_BUFX2_820 ( );
FILL FILL_0_BUFX2_780 ( );
FILL FILL_1_BUFX2_780 ( );
FILL FILL_0_BUFX2_884 ( );
FILL FILL_1_BUFX2_884 ( );
FILL FILL_0_BUFX2_844 ( );
FILL FILL_0_OAI21X1_898 ( );
FILL FILL_1_OAI21X1_898 ( );
FILL FILL_0_NAND2X1_392 ( );
FILL FILL_1_NAND2X1_392 ( );
FILL FILL_0_DFFPOSX1_21 ( );
FILL FILL_1_DFFPOSX1_21 ( );
FILL FILL_2_DFFPOSX1_21 ( );
FILL FILL_3_DFFPOSX1_21 ( );
FILL FILL_4_DFFPOSX1_21 ( );
FILL FILL_5_DFFPOSX1_21 ( );
FILL FILL_0_DFFPOSX1_153 ( );
FILL FILL_1_DFFPOSX1_153 ( );
FILL FILL_2_DFFPOSX1_153 ( );
FILL FILL_3_DFFPOSX1_153 ( );
FILL FILL_4_DFFPOSX1_153 ( );
FILL FILL_5_DFFPOSX1_153 ( );
FILL FILL_0_DFFPOSX1_178 ( );
FILL FILL_1_DFFPOSX1_178 ( );
FILL FILL_2_DFFPOSX1_178 ( );
FILL FILL_3_DFFPOSX1_178 ( );
FILL FILL_4_DFFPOSX1_178 ( );
FILL FILL_5_DFFPOSX1_178 ( );
FILL FILL_6_DFFPOSX1_178 ( );
FILL FILL_0_DFFPOSX1_19 ( );
FILL FILL_1_DFFPOSX1_19 ( );
FILL FILL_2_DFFPOSX1_19 ( );
FILL FILL_3_DFFPOSX1_19 ( );
FILL FILL_4_DFFPOSX1_19 ( );
FILL FILL_5_DFFPOSX1_19 ( );
FILL FILL_0_NAND2X1_697 ( );
FILL FILL_1_NAND2X1_697 ( );
FILL FILL_0_DFFPOSX1_1019 ( );
FILL FILL_1_DFFPOSX1_1019 ( );
FILL FILL_2_DFFPOSX1_1019 ( );
FILL FILL_3_DFFPOSX1_1019 ( );
FILL FILL_4_DFFPOSX1_1019 ( );
FILL FILL_5_DFFPOSX1_1019 ( );
FILL FILL_6_DFFPOSX1_1019 ( );
FILL FILL_0_OAI21X1_948 ( );
FILL FILL_1_OAI21X1_948 ( );
FILL FILL_0_BUFX2_680 ( );
FILL FILL_0_OAI21X1_1788 ( );
FILL FILL_1_OAI21X1_1788 ( );
FILL FILL_0_NAND2X1_729 ( );
FILL FILL_1_NAND2X1_729 ( );
FILL FILL_0_DFFPOSX1_114 ( );
FILL FILL_1_DFFPOSX1_114 ( );
FILL FILL_2_DFFPOSX1_114 ( );
FILL FILL_3_DFFPOSX1_114 ( );
FILL FILL_4_DFFPOSX1_114 ( );
FILL FILL_5_DFFPOSX1_114 ( );
FILL FILL_0_OAI21X1_100 ( );
FILL FILL_1_OAI21X1_100 ( );
FILL FILL_0_OAI21X1_101 ( );
FILL FILL_1_OAI21X1_101 ( );
FILL FILL_0_OAI21X1_229 ( );
FILL FILL_1_OAI21X1_229 ( );
FILL FILL_0_DFFPOSX1_306 ( );
FILL FILL_1_DFFPOSX1_306 ( );
FILL FILL_2_DFFPOSX1_306 ( );
FILL FILL_3_DFFPOSX1_306 ( );
FILL FILL_4_DFFPOSX1_306 ( );
FILL FILL_5_DFFPOSX1_306 ( );
FILL FILL_6_DFFPOSX1_306 ( );
FILL FILL_0_OAI21X1_228 ( );
FILL FILL_1_OAI21X1_228 ( );
FILL FILL_0_BUFX4_60 ( );
FILL FILL_1_BUFX4_60 ( );
FILL FILL_0_BUFX2_745 ( );
FILL FILL_0_OAI21X1_974 ( );
FILL FILL_1_OAI21X1_974 ( );
FILL FILL_0_OAI21X1_254 ( );
FILL FILL_1_OAI21X1_254 ( );
FILL FILL_0_BUFX2_921 ( );
FILL FILL_1_BUFX2_921 ( );
FILL FILL_0_BUFX2_909 ( );
FILL FILL_0_OAI21X1_255 ( );
FILL FILL_1_OAI21X1_255 ( );
FILL FILL_0_DFFPOSX1_191 ( );
FILL FILL_1_DFFPOSX1_191 ( );
FILL FILL_2_DFFPOSX1_191 ( );
FILL FILL_3_DFFPOSX1_191 ( );
FILL FILL_4_DFFPOSX1_191 ( );
FILL FILL_5_DFFPOSX1_191 ( );
FILL FILL_6_DFFPOSX1_191 ( );
FILL FILL_0_OAI21X1_984 ( );
FILL FILL_1_OAI21X1_984 ( );
FILL FILL_0_OAI21X1_985 ( );
FILL FILL_1_OAI21X1_985 ( );
FILL FILL_2_OAI21X1_985 ( );
FILL FILL_0_OAI21X1_1030 ( );
FILL FILL_1_OAI21X1_1030 ( );
FILL FILL_0_BUFX2_385 ( );
FILL FILL_1_BUFX2_385 ( );
FILL FILL_0_OAI21X1_1726 ( );
FILL FILL_1_OAI21X1_1726 ( );
FILL FILL_0_OAI21X1_1756 ( );
FILL FILL_1_OAI21X1_1756 ( );
FILL FILL_0_OAI21X1_1757 ( );
FILL FILL_1_OAI21X1_1757 ( );
FILL FILL_0_DFFPOSX1_91 ( );
FILL FILL_1_DFFPOSX1_91 ( );
FILL FILL_2_DFFPOSX1_91 ( );
FILL FILL_3_DFFPOSX1_91 ( );
FILL FILL_4_DFFPOSX1_91 ( );
FILL FILL_5_DFFPOSX1_91 ( );
FILL FILL_6_DFFPOSX1_91 ( );
FILL FILL_0_BUFX2_761 ( );
FILL FILL_0_OAI21X1_1637 ( );
FILL FILL_1_OAI21X1_1637 ( );
FILL FILL_0_NAND2X1_705 ( );
FILL FILL_1_NAND2X1_705 ( );
FILL FILL_0_DFFPOSX1_27 ( );
FILL FILL_1_DFFPOSX1_27 ( );
FILL FILL_2_DFFPOSX1_27 ( );
FILL FILL_3_DFFPOSX1_27 ( );
FILL FILL_4_DFFPOSX1_27 ( );
FILL FILL_5_DFFPOSX1_27 ( );
FILL FILL_0_OAI21X1_930 ( );
FILL FILL_1_OAI21X1_930 ( );
FILL FILL_0_OAI21X1_931 ( );
FILL FILL_1_OAI21X1_931 ( );
FILL FILL_0_DFFPOSX1_691 ( );
FILL FILL_1_DFFPOSX1_691 ( );
FILL FILL_2_DFFPOSX1_691 ( );
FILL FILL_3_DFFPOSX1_691 ( );
FILL FILL_4_DFFPOSX1_691 ( );
FILL FILL_5_DFFPOSX1_691 ( );
FILL FILL_0_BUFX2_729 ( );
FILL FILL_0_OAI21X1_879 ( );
FILL FILL_1_OAI21X1_879 ( );
FILL FILL_0_INVX1_93 ( );
FILL FILL_0_BUFX2_318 ( );
FILL FILL_1_BUFX2_318 ( );
FILL FILL_0_INVX1_108 ( );
FILL FILL_0_OAI21X1_907 ( );
FILL FILL_1_OAI21X1_907 ( );
FILL FILL_2_OAI21X1_907 ( );
FILL FILL_0_NAND2X1_401 ( );
FILL FILL_0_DFFPOSX1_679 ( );
FILL FILL_1_DFFPOSX1_679 ( );
FILL FILL_2_DFFPOSX1_679 ( );
FILL FILL_3_DFFPOSX1_679 ( );
FILL FILL_4_DFFPOSX1_679 ( );
FILL FILL_5_DFFPOSX1_679 ( );
FILL FILL_6_DFFPOSX1_679 ( );
FILL FILL_0_INVX1_84 ( );
FILL FILL_0_INVX1_123 ( );
FILL FILL_0_BUFX2_322 ( );
FILL FILL_1_BUFX2_322 ( );
FILL FILL_0_NAND2X1_377 ( );
FILL FILL_1_NAND2X1_377 ( );
FILL FILL_0_OAI21X1_883 ( );
FILL FILL_1_OAI21X1_883 ( );
FILL FILL_0_DFFPOSX1_655 ( );
FILL FILL_1_DFFPOSX1_655 ( );
FILL FILL_2_DFFPOSX1_655 ( );
FILL FILL_3_DFFPOSX1_655 ( );
FILL FILL_4_DFFPOSX1_655 ( );
FILL FILL_5_DFFPOSX1_655 ( );
FILL FILL_6_DFFPOSX1_655 ( );
FILL FILL_0_INVX2_179 ( );
FILL FILL_0_INVX1_112 ( );
FILL FILL_0_INVX1_119 ( );
FILL FILL_0_BUFX2_327 ( );
FILL FILL_1_BUFX2_327 ( );
FILL FILL_0_INVX1_133 ( );
FILL FILL_0_BUFX2_342 ( );
FILL FILL_0_BUFX2_932 ( );
FILL FILL_0_OAI21X1_957 ( );
FILL FILL_1_OAI21X1_957 ( );
FILL FILL_0_DFFPOSX1_704 ( );
FILL FILL_1_DFFPOSX1_704 ( );
FILL FILL_2_DFFPOSX1_704 ( );
FILL FILL_3_DFFPOSX1_704 ( );
FILL FILL_4_DFFPOSX1_704 ( );
FILL FILL_5_DFFPOSX1_704 ( );
FILL FILL_0_INVX2_145 ( );
FILL FILL_0_INVX2_165 ( );
FILL FILL_0_INVX2_161 ( );
FILL FILL_0_INVX1_91 ( );
FILL FILL_0_INVX1_101 ( );
FILL FILL_0_BUFX2_310 ( );
FILL FILL_1_BUFX2_310 ( );
FILL FILL_0_OAI21X1_900 ( );
FILL FILL_1_OAI21X1_900 ( );
FILL FILL_2_OAI21X1_900 ( );
FILL FILL_0_NAND2X1_394 ( );
FILL FILL_0_BUFX2_99 ( );
FILL FILL_1_BUFX2_99 ( );
FILL FILL_0_BUFX2_77 ( );
FILL FILL_0_BUFX2_875 ( );
FILL FILL_0_BUFX2_721 ( );
FILL FILL_1_BUFX2_721 ( );
FILL FILL_0_BUFX2_325 ( );
FILL FILL_1_BUFX2_325 ( );
FILL FILL_0_BUFX2_702 ( );
FILL FILL_1_BUFX2_702 ( );
FILL FILL_0_INVX2_133 ( );
FILL FILL_0_INVX2_150 ( );
FILL FILL_0_BUFX2_126 ( );
FILL FILL_0_NAND2X1_468 ( );
FILL FILL_0_OAI21X1_1102 ( );
FILL FILL_1_OAI21X1_1102 ( );
FILL FILL_0_DFFPOSX1_810 ( );
FILL FILL_1_DFFPOSX1_810 ( );
FILL FILL_2_DFFPOSX1_810 ( );
FILL FILL_3_DFFPOSX1_810 ( );
FILL FILL_4_DFFPOSX1_810 ( );
FILL FILL_5_DFFPOSX1_810 ( );
FILL FILL_0_BUFX2_558 ( );
FILL FILL_0_BUFX2_13 ( );
FILL FILL_1_BUFX2_13 ( );
FILL FILL_0_BUFX2_110 ( );
FILL FILL_1_BUFX2_110 ( );
FILL FILL_0_BUFX2_62 ( );
FILL FILL_1_BUFX2_62 ( );
FILL FILL_0_BUFX2_850 ( );
FILL FILL_1_BUFX2_850 ( );
FILL FILL_0_BUFX2_848 ( );
FILL FILL_1_BUFX2_848 ( );
FILL FILL_0_BUFX2_63 ( );
FILL FILL_1_BUFX2_63 ( );
FILL FILL_0_INVX2_163 ( );
FILL FILL_0_NAND2X1_23 ( );
FILL FILL_1_NAND2X1_23 ( );
FILL FILL_0_NAND2X1_25 ( );
FILL FILL_1_NAND2X1_25 ( );
FILL FILL_0_OAI21X1_25 ( );
FILL FILL_1_OAI21X1_25 ( );
FILL FILL_0_DFFPOSX1_181 ( );
FILL FILL_1_DFFPOSX1_181 ( );
FILL FILL_2_DFFPOSX1_181 ( );
FILL FILL_3_DFFPOSX1_181 ( );
FILL FILL_4_DFFPOSX1_181 ( );
FILL FILL_5_DFFPOSX1_181 ( );
FILL FILL_0_BUFX2_976 ( );
FILL FILL_0_BUFX2_914 ( );
FILL FILL_0_BUFX2_24 ( );
FILL FILL_1_BUFX2_24 ( );
FILL FILL_0_BUFX2_511 ( );
FILL FILL_0_BUFX2_881 ( );
FILL FILL_1_BUFX2_881 ( );
FILL FILL_0_BUFX2_195 ( );
FILL FILL_1_BUFX2_195 ( );
FILL FILL_0_BUFX2_141 ( );
FILL FILL_1_BUFX2_141 ( );
FILL FILL_0_BUFX2_198 ( );
FILL FILL_1_BUFX2_198 ( );
FILL FILL_0_BUFX2_939 ( );
FILL FILL_1_BUFX2_939 ( );
FILL FILL_0_INVX2_118 ( );
FILL FILL_0_BUFX2_490 ( );
FILL FILL_0_DFFPOSX1_245 ( );
FILL FILL_1_DFFPOSX1_245 ( );
FILL FILL_2_DFFPOSX1_245 ( );
FILL FILL_3_DFFPOSX1_245 ( );
FILL FILL_4_DFFPOSX1_245 ( );
FILL FILL_5_DFFPOSX1_245 ( );
FILL FILL_6_DFFPOSX1_245 ( );
FILL FILL_0_DFFPOSX1_209 ( );
FILL FILL_1_DFFPOSX1_209 ( );
FILL FILL_2_DFFPOSX1_209 ( );
FILL FILL_3_DFFPOSX1_209 ( );
FILL FILL_4_DFFPOSX1_209 ( );
FILL FILL_5_DFFPOSX1_209 ( );
FILL FILL_0_NAND2X1_53 ( );
FILL FILL_1_NAND2X1_53 ( );
FILL FILL_0_OAI21X1_53 ( );
FILL FILL_1_OAI21X1_53 ( );
FILL FILL_0_INVX2_191 ( );
FILL FILL_0_BUFX2_805 ( );
FILL FILL_0_DFFPOSX1_134 ( );
FILL FILL_1_DFFPOSX1_134 ( );
FILL FILL_2_DFFPOSX1_134 ( );
FILL FILL_3_DFFPOSX1_134 ( );
FILL FILL_4_DFFPOSX1_134 ( );
FILL FILL_5_DFFPOSX1_134 ( );
FILL FILL_0_NAND2X1_749 ( );
FILL FILL_1_NAND2X1_749 ( );
FILL FILL_0_OAI21X1_1808 ( );
FILL FILL_1_OAI21X1_1808 ( );
FILL FILL_0_BUFX2_578 ( );
FILL FILL_1_BUFX2_578 ( );
FILL FILL_0_BUFX2_448 ( );
FILL FILL_1_BUFX2_448 ( );
FILL FILL_0_BUFX2_517 ( );
FILL FILL_1_BUFX2_517 ( );
FILL FILL_0_BUFX2_650 ( );
FILL FILL_1_BUFX2_650 ( );
FILL FILL_0_NAND2X1_651 ( );
FILL FILL_0_OAI21X1_1582 ( );
FILL FILL_1_OAI21X1_1582 ( );
FILL FILL_0_DFFPOSX1_1005 ( );
FILL FILL_1_DFFPOSX1_1005 ( );
FILL FILL_2_DFFPOSX1_1005 ( );
FILL FILL_3_DFFPOSX1_1005 ( );
FILL FILL_4_DFFPOSX1_1005 ( );
FILL FILL_5_DFFPOSX1_1005 ( );
FILL FILL_0_BUFX2_978 ( );
FILL FILL_1_BUFX2_978 ( );
FILL FILL_0_BUFX2_682 ( );
FILL FILL_1_BUFX2_682 ( );
FILL FILL_0_BUFX2_403 ( );
FILL FILL_1_BUFX2_403 ( );
FILL FILL_0_NAND2X1_683 ( );
FILL FILL_1_NAND2X1_683 ( );
FILL FILL_0_OAI21X1_1615 ( );
FILL FILL_1_OAI21X1_1615 ( );
FILL FILL_0_BUFX2_70 ( );
FILL FILL_1_BUFX2_70 ( );
FILL FILL_0_NAND2X1_491 ( );
FILL FILL_1_NAND2X1_491 ( );
FILL FILL_0_DFFPOSX1_821 ( );
FILL FILL_1_DFFPOSX1_821 ( );
FILL FILL_2_DFFPOSX1_821 ( );
FILL FILL_3_DFFPOSX1_821 ( );
FILL FILL_4_DFFPOSX1_821 ( );
FILL FILL_5_DFFPOSX1_821 ( );
FILL FILL_0_BUFX2_786 ( );
FILL FILL_1_BUFX2_786 ( );
FILL FILL_0_BUFX2_811 ( );
FILL FILL_1_BUFX2_811 ( );
FILL FILL_0_BUFX2_139 ( );
FILL FILL_0_BUFX2_1003 ( );
FILL FILL_1_BUFX2_1003 ( );
FILL FILL_0_INVX1_169 ( );
FILL FILL_0_BUFX2_380 ( );
FILL FILL_1_BUFX2_380 ( );
FILL FILL_0_INVX1_144 ( );
FILL FILL_0_DFFPOSX1_715 ( );
FILL FILL_1_DFFPOSX1_715 ( );
FILL FILL_2_DFFPOSX1_715 ( );
FILL FILL_3_DFFPOSX1_715 ( );
FILL FILL_4_DFFPOSX1_715 ( );
FILL FILL_5_DFFPOSX1_715 ( );
FILL FILL_6_DFFPOSX1_715 ( );
FILL FILL_0_BUFX2_969 ( );
FILL FILL_0_DFFPOSX1_273 ( );
FILL FILL_1_DFFPOSX1_273 ( );
FILL FILL_2_DFFPOSX1_273 ( );
FILL FILL_3_DFFPOSX1_273 ( );
FILL FILL_4_DFFPOSX1_273 ( );
FILL FILL_5_DFFPOSX1_273 ( );
FILL FILL_6_DFFPOSX1_273 ( );
FILL FILL_0_BUFX2_945 ( );
FILL FILL_0_BUFX2_957 ( );
FILL FILL_1_BUFX2_957 ( );
FILL FILL_0_BUFX2_986 ( );
FILL FILL_1_BUFX2_986 ( );
FILL FILL_0_BUFX2_1021 ( );
FILL FILL_0_BUFX2_830 ( );
FILL FILL_1_BUFX2_830 ( );
FILL FILL_0_BUFX2_664 ( );
FILL FILL_0_DFFPOSX1_220 ( );
FILL FILL_1_DFFPOSX1_220 ( );
FILL FILL_2_DFFPOSX1_220 ( );
FILL FILL_3_DFFPOSX1_220 ( );
FILL FILL_4_DFFPOSX1_220 ( );
FILL FILL_5_DFFPOSX1_220 ( );
FILL FILL_0_OAI21X1_64 ( );
FILL FILL_1_OAI21X1_64 ( );
FILL FILL_0_BUFX2_958 ( );
FILL FILL_0_NAND2X1_64 ( );
FILL FILL_1_NAND2X1_64 ( );
FILL FILL_0_BUFX2_849 ( );
FILL FILL_0_BUFX2_893 ( );
FILL FILL_0_INVX2_1 ( );
FILL FILL_1_INVX2_1 ( );
FILL FILL_0_INVX2_202 ( );
FILL FILL_0_INVX2_139 ( );
FILL FILL_0_OAI21X1_1621 ( );
FILL FILL_1_OAI21X1_1621 ( );
FILL FILL_0_NAND2X1_689 ( );
FILL FILL_1_NAND2X1_689 ( );
FILL FILL_0_INVX2_124 ( );
FILL FILL_0_BUFX2_829 ( );
FILL FILL_1_BUFX2_829 ( );
FILL FILL_0_DFFPOSX1_11 ( );
FILL FILL_1_DFFPOSX1_11 ( );
FILL FILL_2_DFFPOSX1_11 ( );
FILL FILL_3_DFFPOSX1_11 ( );
FILL FILL_4_DFFPOSX1_11 ( );
FILL FILL_5_DFFPOSX1_11 ( );
FILL FILL_6_DFFPOSX1_11 ( );
FILL FILL_0_INVX2_170 ( );
FILL FILL_0_BUFX2_801 ( );
FILL FILL_1_BUFX2_801 ( );
FILL FILL_0_BUFX2_1011 ( );
FILL FILL_1_BUFX2_1011 ( );
FILL FILL_0_BUFX2_710 ( );
FILL FILL_1_BUFX2_710 ( );
FILL FILL_0_INVX2_193 ( );
FILL FILL_0_BUFX2_988 ( );
FILL FILL_1_BUFX2_988 ( );
FILL FILL_0_BUFX2_999 ( );
FILL FILL_1_BUFX2_999 ( );
FILL FILL_0_BUFX2_736 ( );
FILL FILL_1_BUFX2_736 ( );
FILL FILL_0_INVX2_130 ( );
FILL FILL_1_INVX2_130 ( );
FILL FILL_0_BUFX2_880 ( );
FILL FILL_0_BUFX2_654 ( );
FILL FILL_0_INVX2_190 ( );
FILL FILL_0_BUFX2_796 ( );
FILL FILL_1_BUFX2_796 ( );
FILL FILL_0_BUFX2_860 ( );
FILL FILL_1_BUFX2_860 ( );
FILL FILL_0_BUFX2_795 ( );
FILL FILL_1_BUFX2_795 ( );
FILL FILL_0_BUFX2_271 ( );
FILL FILL_1_BUFX2_271 ( );
FILL FILL_0_BUFX2_915 ( );
FILL FILL_1_BUFX2_915 ( );
FILL FILL_0_BUFX2_924 ( );
FILL FILL_0_INVX2_194 ( );
FILL FILL_0_INVX2_172 ( );
FILL FILL_0_BUFX2_987 ( );
FILL FILL_0_BUFX2_908 ( );
FILL FILL_1_BUFX2_908 ( );
FILL FILL_0_BUFX2_890 ( );
FILL FILL_1_BUFX2_890 ( );
FILL FILL_0_BUFX2_826 ( );
FILL FILL_0_BUFX2_308 ( );
FILL FILL_0_BUFX2_690 ( );
FILL FILL_0_BUFX2_82 ( );
FILL FILL_0_INVX2_157 ( );
FILL FILL_0_INVX1_99 ( );
FILL FILL_0_DFFPOSX1_13 ( );
FILL FILL_1_DFFPOSX1_13 ( );
FILL FILL_2_DFFPOSX1_13 ( );
FILL FILL_3_DFFPOSX1_13 ( );
FILL FILL_4_DFFPOSX1_13 ( );
FILL FILL_5_DFFPOSX1_13 ( );
FILL FILL_6_DFFPOSX1_13 ( );
FILL FILL_0_INVX1_140 ( );
FILL FILL_1_INVX1_140 ( );
FILL FILL_0_OAI21X1_1623 ( );
FILL FILL_1_OAI21X1_1623 ( );
FILL FILL_0_INVX2_199 ( );
FILL FILL_0_NAND2X1_691 ( );
FILL FILL_1_NAND2X1_691 ( );
FILL FILL_0_BUFX2_712 ( );
FILL FILL_1_BUFX2_712 ( );
FILL FILL_0_INVX2_134 ( );
FILL FILL_0_BUFX2_656 ( );
FILL FILL_1_BUFX2_656 ( );
FILL FILL_0_OAI21X1_22 ( );
FILL FILL_1_OAI21X1_22 ( );
FILL FILL_0_NAND2X1_22 ( );
FILL FILL_1_NAND2X1_22 ( );
FILL FILL_0_BUFX2_847 ( );
FILL FILL_1_BUFX2_847 ( );
FILL FILL_0_BUFX2_688 ( );
FILL FILL_0_BUFX2_943 ( );
FILL FILL_0_DFFPOSX1_700 ( );
FILL FILL_1_DFFPOSX1_700 ( );
FILL FILL_2_DFFPOSX1_700 ( );
FILL FILL_3_DFFPOSX1_700 ( );
FILL FILL_4_DFFPOSX1_700 ( );
FILL FILL_5_DFFPOSX1_700 ( );
FILL FILL_6_DFFPOSX1_700 ( );
FILL FILL_0_BUFX2_887 ( );
FILL FILL_1_BUFX2_887 ( );
FILL FILL_0_BUFX2_338 ( );
FILL FILL_1_BUFX2_338 ( );
FILL FILL_0_OAI21X1_949 ( );
FILL FILL_1_OAI21X1_949 ( );
FILL FILL_2_OAI21X1_949 ( );
FILL FILL_0_INVX1_129 ( );
FILL FILL_0_INVX2_160 ( );
FILL FILL_0_INVX2_180 ( );
FILL FILL_0_BUFX2_869 ( );
FILL FILL_1_BUFX2_869 ( );
FILL FILL_0_BUFX2_783 ( );
FILL FILL_1_BUFX2_783 ( );
FILL FILL_0_DFFPOSX1_342 ( );
FILL FILL_1_DFFPOSX1_342 ( );
FILL FILL_2_DFFPOSX1_342 ( );
FILL FILL_3_DFFPOSX1_342 ( );
FILL FILL_4_DFFPOSX1_342 ( );
FILL FILL_5_DFFPOSX1_342 ( );
FILL FILL_0_OAI21X1_301 ( );
FILL FILL_1_OAI21X1_301 ( );
FILL FILL_0_BUFX2_911 ( );
FILL FILL_0_OAI21X1_300 ( );
FILL FILL_1_OAI21X1_300 ( );
FILL FILL_0_BUFX2_1015 ( );
FILL FILL_0_INVX2_196 ( );
FILL FILL_0_DFFPOSX1_713 ( );
FILL FILL_1_DFFPOSX1_713 ( );
FILL FILL_2_DFFPOSX1_713 ( );
FILL FILL_3_DFFPOSX1_713 ( );
FILL FILL_4_DFFPOSX1_713 ( );
FILL FILL_5_DFFPOSX1_713 ( );
FILL FILL_6_DFFPOSX1_713 ( );
FILL FILL_0_BUFX2_975 ( );
FILL FILL_1_BUFX2_975 ( );
FILL FILL_0_OAI21X1_975 ( );
FILL FILL_1_OAI21X1_975 ( );
FILL FILL_2_OAI21X1_975 ( );
FILL FILL_0_INVX1_142 ( );
FILL FILL_0_BUFX2_358 ( );
FILL FILL_0_BUFX2_989 ( );
FILL FILL_0_DFFPOSX1_741 ( );
FILL FILL_1_DFFPOSX1_741 ( );
FILL FILL_2_DFFPOSX1_741 ( );
FILL FILL_3_DFFPOSX1_741 ( );
FILL FILL_4_DFFPOSX1_741 ( );
FILL FILL_5_DFFPOSX1_741 ( );
FILL FILL_6_DFFPOSX1_741 ( );
FILL FILL_0_OAI21X1_1031 ( );
FILL FILL_1_OAI21X1_1031 ( );
FILL FILL_0_INVX1_170 ( );
FILL FILL_0_BUFX2_861 ( );
FILL FILL_1_BUFX2_861 ( );
FILL FILL_0_BUFX2_379 ( );
FILL FILL_1_BUFX2_379 ( );
FILL FILL_0_INVX1_147 ( );
FILL FILL_0_DFFPOSX1_127 ( );
FILL FILL_1_DFFPOSX1_127 ( );
FILL FILL_2_DFFPOSX1_127 ( );
FILL FILL_3_DFFPOSX1_127 ( );
FILL FILL_4_DFFPOSX1_127 ( );
FILL FILL_5_DFFPOSX1_127 ( );
FILL FILL_0_OAI21X1_1801 ( );
FILL FILL_1_OAI21X1_1801 ( );
FILL FILL_0_NAND2X1_742 ( );
FILL FILL_1_NAND2X1_742 ( );
FILL FILL_0_BUFX2_797 ( );
FILL FILL_0_BUFX2_775 ( );
FILL FILL_1_BUFX2_775 ( );
FILL FILL_0_DFFPOSX1_1027 ( );
FILL FILL_1_DFFPOSX1_1027 ( );
FILL FILL_2_DFFPOSX1_1027 ( );
FILL FILL_3_DFFPOSX1_1027 ( );
FILL FILL_4_DFFPOSX1_1027 ( );
FILL FILL_5_DFFPOSX1_1027 ( );
FILL FILL_6_DFFPOSX1_1027 ( );
FILL FILL_0_OAI21X1_1604 ( );
FILL FILL_1_OAI21X1_1604 ( );
FILL FILL_0_NAND2X1_673 ( );
FILL FILL_1_NAND2X1_673 ( );
FILL FILL_0_INVX2_126 ( );
FILL FILL_0_INVX2_140 ( );
FILL FILL_0_INVX2_189 ( );
FILL FILL_0_INVX2_125 ( );
FILL FILL_0_BUFX2_697 ( );
FILL FILL_1_BUFX2_697 ( );
FILL FILL_0_INVX2_158 ( );
FILL FILL_1_INVX2_158 ( );
FILL FILL_0_BUFX2_665 ( );
FILL FILL_1_BUFX2_665 ( );
FILL FILL_0_INVX2_173 ( );
FILL FILL_0_INVX1_120 ( );
FILL FILL_0_OAI21X1_882 ( );
FILL FILL_1_OAI21X1_882 ( );
FILL FILL_0_DFFPOSX1_654 ( );
FILL FILL_1_DFFPOSX1_654 ( );
FILL FILL_2_DFFPOSX1_654 ( );
FILL FILL_3_DFFPOSX1_654 ( );
FILL FILL_4_DFFPOSX1_654 ( );
FILL FILL_5_DFFPOSX1_654 ( );
FILL FILL_0_0_0 ( );
FILL FILL_0_0_1 ( );
FILL FILL_0_1_0 ( );
FILL FILL_0_1_1 ( );
FILL FILL_0_2_0 ( );
FILL FILL_0_2_1 ( );
FILL FILL_0_3_0 ( );
FILL FILL_0_3_1 ( );
FILL FILL_0_4_0 ( );
FILL FILL_0_4_1 ( );
FILL FILL_0_5_0 ( );
FILL FILL_0_5_1 ( );
FILL FILL_0_6_0 ( );
FILL FILL_0_6_1 ( );
FILL FILL_0_7_0 ( );
FILL FILL_0_7_1 ( );
FILL FILL_0_8_0 ( );
FILL FILL_0_8_1 ( );
FILL FILL_0_9_0 ( );
FILL FILL_0_9_1 ( );
FILL FILL_0_10_0 ( );
FILL FILL_0_10_1 ( );
FILL FILL_0_11_0 ( );
FILL FILL_0_11_1 ( );
FILL FILL_0_12_0 ( );
FILL FILL_0_12_1 ( );
FILL FILL_0_13_0 ( );
FILL FILL_0_13_1 ( );
FILL FILL_0_14_0 ( );
FILL FILL_0_14_1 ( );
FILL FILL_0_15_0 ( );
FILL FILL_0_15_1 ( );
FILL FILL_0_16_0 ( );
FILL FILL_0_16_1 ( );
FILL FILL_0_17_0 ( );
FILL FILL_0_17_1 ( );
FILL FILL_0_18_0 ( );
FILL FILL_0_18_1 ( );
FILL FILL_1_1 ( );
FILL FILL_1_0_0 ( );
FILL FILL_1_0_1 ( );
FILL FILL_1_1_0 ( );
FILL FILL_1_1_1 ( );
FILL FILL_1_2_0 ( );
FILL FILL_1_2_1 ( );
FILL FILL_1_3_0 ( );
FILL FILL_1_3_1 ( );
FILL FILL_1_4_0 ( );
FILL FILL_1_4_1 ( );
FILL FILL_1_5_0 ( );
FILL FILL_1_5_1 ( );
FILL FILL_1_6_0 ( );
FILL FILL_1_6_1 ( );
FILL FILL_1_7_0 ( );
FILL FILL_1_7_1 ( );
FILL FILL_1_8_0 ( );
FILL FILL_1_8_1 ( );
FILL FILL_1_9_0 ( );
FILL FILL_1_9_1 ( );
FILL FILL_1_10_0 ( );
FILL FILL_1_10_1 ( );
FILL FILL_1_11_0 ( );
FILL FILL_1_11_1 ( );
FILL FILL_1_12_0 ( );
FILL FILL_1_12_1 ( );
FILL FILL_1_13_0 ( );
FILL FILL_1_13_1 ( );
FILL FILL_1_14_0 ( );
FILL FILL_1_14_1 ( );
FILL FILL_1_15_0 ( );
FILL FILL_1_15_1 ( );
FILL FILL_1_16_0 ( );
FILL FILL_1_16_1 ( );
FILL FILL_1_17_0 ( );
FILL FILL_1_17_1 ( );
FILL FILL_1_18_0 ( );
FILL FILL_1_18_1 ( );
FILL FILL_2_1 ( );
FILL FILL_2_0_0 ( );
FILL FILL_2_0_1 ( );
FILL FILL_2_1_0 ( );
FILL FILL_2_1_1 ( );
FILL FILL_2_2_0 ( );
FILL FILL_2_2_1 ( );
FILL FILL_2_3_0 ( );
FILL FILL_2_3_1 ( );
FILL FILL_2_4_0 ( );
FILL FILL_2_4_1 ( );
FILL FILL_2_5_0 ( );
FILL FILL_2_5_1 ( );
FILL FILL_2_6_0 ( );
FILL FILL_2_6_1 ( );
FILL FILL_2_7_0 ( );
FILL FILL_2_7_1 ( );
FILL FILL_2_8_0 ( );
FILL FILL_2_8_1 ( );
FILL FILL_2_9_0 ( );
FILL FILL_2_9_1 ( );
FILL FILL_2_10_0 ( );
FILL FILL_2_10_1 ( );
FILL FILL_2_11_0 ( );
FILL FILL_2_11_1 ( );
FILL FILL_2_12_0 ( );
FILL FILL_2_12_1 ( );
FILL FILL_2_13_0 ( );
FILL FILL_2_13_1 ( );
FILL FILL_2_14_0 ( );
FILL FILL_2_14_1 ( );
FILL FILL_2_15_0 ( );
FILL FILL_2_15_1 ( );
FILL FILL_2_16_0 ( );
FILL FILL_2_16_1 ( );
FILL FILL_2_17_0 ( );
FILL FILL_2_17_1 ( );
FILL FILL_2_18_0 ( );
FILL FILL_2_18_1 ( );
FILL FILL_3_1 ( );
FILL FILL_3_0_0 ( );
FILL FILL_3_0_1 ( );
FILL FILL_3_1_0 ( );
FILL FILL_3_1_1 ( );
FILL FILL_3_2_0 ( );
FILL FILL_3_2_1 ( );
FILL FILL_3_3_0 ( );
FILL FILL_3_3_1 ( );
FILL FILL_3_4_0 ( );
FILL FILL_3_4_1 ( );
FILL FILL_3_5_0 ( );
FILL FILL_3_5_1 ( );
FILL FILL_3_6_0 ( );
FILL FILL_3_6_1 ( );
FILL FILL_3_7_0 ( );
FILL FILL_3_7_1 ( );
FILL FILL_3_8_0 ( );
FILL FILL_3_8_1 ( );
FILL FILL_3_9_0 ( );
FILL FILL_3_9_1 ( );
FILL FILL_3_10_0 ( );
FILL FILL_3_10_1 ( );
FILL FILL_3_11_0 ( );
FILL FILL_3_11_1 ( );
FILL FILL_3_12_0 ( );
FILL FILL_3_12_1 ( );
FILL FILL_3_13_0 ( );
FILL FILL_3_13_1 ( );
FILL FILL_3_14_0 ( );
FILL FILL_3_14_1 ( );
FILL FILL_3_15_0 ( );
FILL FILL_3_15_1 ( );
FILL FILL_3_16_0 ( );
FILL FILL_3_16_1 ( );
FILL FILL_3_17_0 ( );
FILL FILL_3_17_1 ( );
FILL FILL_3_18_0 ( );
FILL FILL_3_18_1 ( );
FILL FILL_4_1 ( );
FILL FILL_4_2 ( );
FILL FILL_4_3 ( );
FILL FILL_4_0_0 ( );
FILL FILL_4_0_1 ( );
FILL FILL_4_1_0 ( );
FILL FILL_4_1_1 ( );
FILL FILL_4_2_0 ( );
FILL FILL_4_2_1 ( );
FILL FILL_4_3_0 ( );
FILL FILL_4_3_1 ( );
FILL FILL_4_4_0 ( );
FILL FILL_4_4_1 ( );
FILL FILL_4_5_0 ( );
FILL FILL_4_5_1 ( );
FILL FILL_4_6_0 ( );
FILL FILL_4_6_1 ( );
FILL FILL_4_7_0 ( );
FILL FILL_4_7_1 ( );
FILL FILL_4_8_0 ( );
FILL FILL_4_8_1 ( );
FILL FILL_4_9_0 ( );
FILL FILL_4_9_1 ( );
FILL FILL_4_10_0 ( );
FILL FILL_4_10_1 ( );
FILL FILL_4_11_0 ( );
FILL FILL_4_11_1 ( );
FILL FILL_4_12_0 ( );
FILL FILL_4_12_1 ( );
FILL FILL_4_13_0 ( );
FILL FILL_4_13_1 ( );
FILL FILL_4_14_0 ( );
FILL FILL_4_14_1 ( );
FILL FILL_4_15_0 ( );
FILL FILL_4_15_1 ( );
FILL FILL_4_16_0 ( );
FILL FILL_4_16_1 ( );
FILL FILL_4_17_0 ( );
FILL FILL_4_17_1 ( );
FILL FILL_4_18_0 ( );
FILL FILL_4_18_1 ( );
FILL FILL_5_1 ( );
FILL FILL_5_2 ( );
FILL FILL_5_3 ( );
FILL FILL_5_0_0 ( );
FILL FILL_5_0_1 ( );
FILL FILL_5_1_0 ( );
FILL FILL_5_1_1 ( );
FILL FILL_5_2_0 ( );
FILL FILL_5_2_1 ( );
FILL FILL_5_3_0 ( );
FILL FILL_5_3_1 ( );
FILL FILL_5_4_0 ( );
FILL FILL_5_4_1 ( );
FILL FILL_5_5_0 ( );
FILL FILL_5_5_1 ( );
FILL FILL_5_6_0 ( );
FILL FILL_5_6_1 ( );
FILL FILL_5_7_0 ( );
FILL FILL_5_7_1 ( );
FILL FILL_5_8_0 ( );
FILL FILL_5_8_1 ( );
FILL FILL_5_9_0 ( );
FILL FILL_5_9_1 ( );
FILL FILL_5_10_0 ( );
FILL FILL_5_10_1 ( );
FILL FILL_5_11_0 ( );
FILL FILL_5_11_1 ( );
FILL FILL_5_12_0 ( );
FILL FILL_5_12_1 ( );
FILL FILL_5_13_0 ( );
FILL FILL_5_13_1 ( );
FILL FILL_5_14_0 ( );
FILL FILL_5_14_1 ( );
FILL FILL_5_15_0 ( );
FILL FILL_5_15_1 ( );
FILL FILL_5_16_0 ( );
FILL FILL_5_16_1 ( );
FILL FILL_5_17_0 ( );
FILL FILL_5_17_1 ( );
FILL FILL_5_18_0 ( );
FILL FILL_5_18_1 ( );
FILL FILL_6_1 ( );
FILL FILL_6_2 ( );
FILL FILL_6_3 ( );
FILL FILL_6_0_0 ( );
FILL FILL_6_0_1 ( );
FILL FILL_6_1_0 ( );
FILL FILL_6_1_1 ( );
FILL FILL_6_2_0 ( );
FILL FILL_6_2_1 ( );
FILL FILL_6_3_0 ( );
FILL FILL_6_3_1 ( );
FILL FILL_6_4_0 ( );
FILL FILL_6_4_1 ( );
FILL FILL_6_5_0 ( );
FILL FILL_6_5_1 ( );
FILL FILL_6_6_0 ( );
FILL FILL_6_6_1 ( );
FILL FILL_6_7_0 ( );
FILL FILL_6_7_1 ( );
FILL FILL_6_8_0 ( );
FILL FILL_6_8_1 ( );
FILL FILL_6_9_0 ( );
FILL FILL_6_9_1 ( );
FILL FILL_6_10_0 ( );
FILL FILL_6_10_1 ( );
FILL FILL_6_11_0 ( );
FILL FILL_6_11_1 ( );
FILL FILL_6_12_0 ( );
FILL FILL_6_12_1 ( );
FILL FILL_6_13_0 ( );
FILL FILL_6_13_1 ( );
FILL FILL_6_14_0 ( );
FILL FILL_6_14_1 ( );
FILL FILL_6_15_0 ( );
FILL FILL_6_15_1 ( );
FILL FILL_6_16_0 ( );
FILL FILL_6_16_1 ( );
FILL FILL_6_17_0 ( );
FILL FILL_6_17_1 ( );
FILL FILL_6_18_0 ( );
FILL FILL_6_18_1 ( );
FILL FILL_7_1 ( );
FILL FILL_7_2 ( );
FILL FILL_7_3 ( );
FILL FILL_7_0_0 ( );
FILL FILL_7_0_1 ( );
FILL FILL_7_1_0 ( );
FILL FILL_7_1_1 ( );
FILL FILL_7_2_0 ( );
FILL FILL_7_2_1 ( );
FILL FILL_7_3_0 ( );
FILL FILL_7_3_1 ( );
FILL FILL_7_4_0 ( );
FILL FILL_7_4_1 ( );
FILL FILL_7_5_0 ( );
FILL FILL_7_5_1 ( );
FILL FILL_7_6_0 ( );
FILL FILL_7_6_1 ( );
FILL FILL_7_7_0 ( );
FILL FILL_7_7_1 ( );
FILL FILL_7_8_0 ( );
FILL FILL_7_8_1 ( );
FILL FILL_7_9_0 ( );
FILL FILL_7_9_1 ( );
FILL FILL_7_10_0 ( );
FILL FILL_7_10_1 ( );
FILL FILL_7_11_0 ( );
FILL FILL_7_11_1 ( );
FILL FILL_7_12_0 ( );
FILL FILL_7_12_1 ( );
FILL FILL_7_13_0 ( );
FILL FILL_7_13_1 ( );
FILL FILL_7_14_0 ( );
FILL FILL_7_14_1 ( );
FILL FILL_7_15_0 ( );
FILL FILL_7_15_1 ( );
FILL FILL_7_16_0 ( );
FILL FILL_7_16_1 ( );
FILL FILL_7_17_0 ( );
FILL FILL_7_17_1 ( );
FILL FILL_7_18_0 ( );
FILL FILL_7_18_1 ( );
FILL FILL_8_1 ( );
FILL FILL_8_0_0 ( );
FILL FILL_8_0_1 ( );
FILL FILL_8_1_0 ( );
FILL FILL_8_1_1 ( );
FILL FILL_8_2_0 ( );
FILL FILL_8_2_1 ( );
FILL FILL_8_3_0 ( );
FILL FILL_8_3_1 ( );
FILL FILL_8_4_0 ( );
FILL FILL_8_4_1 ( );
FILL FILL_8_5_0 ( );
FILL FILL_8_5_1 ( );
FILL FILL_8_6_0 ( );
FILL FILL_8_6_1 ( );
FILL FILL_8_7_0 ( );
FILL FILL_8_7_1 ( );
FILL FILL_8_8_0 ( );
FILL FILL_8_8_1 ( );
FILL FILL_8_9_0 ( );
FILL FILL_8_9_1 ( );
FILL FILL_8_10_0 ( );
FILL FILL_8_10_1 ( );
FILL FILL_8_11_0 ( );
FILL FILL_8_11_1 ( );
FILL FILL_8_12_0 ( );
FILL FILL_8_12_1 ( );
FILL FILL_8_13_0 ( );
FILL FILL_8_13_1 ( );
FILL FILL_8_14_0 ( );
FILL FILL_8_14_1 ( );
FILL FILL_8_15_0 ( );
FILL FILL_8_15_1 ( );
FILL FILL_8_16_0 ( );
FILL FILL_8_16_1 ( );
FILL FILL_8_17_0 ( );
FILL FILL_8_17_1 ( );
FILL FILL_8_18_0 ( );
FILL FILL_8_18_1 ( );
FILL FILL_9_0_0 ( );
FILL FILL_9_0_1 ( );
FILL FILL_9_1_0 ( );
FILL FILL_9_1_1 ( );
FILL FILL_9_2_0 ( );
FILL FILL_9_2_1 ( );
FILL FILL_9_3_0 ( );
FILL FILL_9_3_1 ( );
FILL FILL_9_4_0 ( );
FILL FILL_9_4_1 ( );
FILL FILL_9_5_0 ( );
FILL FILL_9_5_1 ( );
FILL FILL_9_6_0 ( );
FILL FILL_9_6_1 ( );
FILL FILL_9_7_0 ( );
FILL FILL_9_7_1 ( );
FILL FILL_9_8_0 ( );
FILL FILL_9_8_1 ( );
FILL FILL_9_9_0 ( );
FILL FILL_9_9_1 ( );
FILL FILL_9_10_0 ( );
FILL FILL_9_10_1 ( );
FILL FILL_9_11_0 ( );
FILL FILL_9_11_1 ( );
FILL FILL_9_12_0 ( );
FILL FILL_9_12_1 ( );
FILL FILL_9_13_0 ( );
FILL FILL_9_13_1 ( );
FILL FILL_9_14_0 ( );
FILL FILL_9_14_1 ( );
FILL FILL_9_15_0 ( );
FILL FILL_9_15_1 ( );
FILL FILL_9_16_0 ( );
FILL FILL_9_16_1 ( );
FILL FILL_9_17_0 ( );
FILL FILL_9_17_1 ( );
FILL FILL_9_18_0 ( );
FILL FILL_9_18_1 ( );
FILL FILL_10_1 ( );
FILL FILL_10_0_0 ( );
FILL FILL_10_0_1 ( );
FILL FILL_10_1_0 ( );
FILL FILL_10_1_1 ( );
FILL FILL_10_2_0 ( );
FILL FILL_10_2_1 ( );
FILL FILL_10_3_0 ( );
FILL FILL_10_3_1 ( );
FILL FILL_10_4_0 ( );
FILL FILL_10_4_1 ( );
FILL FILL_10_5_0 ( );
FILL FILL_10_5_1 ( );
FILL FILL_10_6_0 ( );
FILL FILL_10_6_1 ( );
FILL FILL_10_7_0 ( );
FILL FILL_10_7_1 ( );
FILL FILL_10_8_0 ( );
FILL FILL_10_8_1 ( );
FILL FILL_10_9_0 ( );
FILL FILL_10_9_1 ( );
FILL FILL_10_10_0 ( );
FILL FILL_10_10_1 ( );
FILL FILL_10_11_0 ( );
FILL FILL_10_11_1 ( );
FILL FILL_10_12_0 ( );
FILL FILL_10_12_1 ( );
FILL FILL_10_13_0 ( );
FILL FILL_10_13_1 ( );
FILL FILL_10_14_0 ( );
FILL FILL_10_14_1 ( );
FILL FILL_10_15_0 ( );
FILL FILL_10_15_1 ( );
FILL FILL_10_16_0 ( );
FILL FILL_10_16_1 ( );
FILL FILL_10_17_0 ( );
FILL FILL_10_17_1 ( );
FILL FILL_10_18_0 ( );
FILL FILL_10_18_1 ( );
FILL FILL_11_1 ( );
FILL FILL_11_0_0 ( );
FILL FILL_11_0_1 ( );
FILL FILL_11_1_0 ( );
FILL FILL_11_1_1 ( );
FILL FILL_11_2_0 ( );
FILL FILL_11_2_1 ( );
FILL FILL_11_3_0 ( );
FILL FILL_11_3_1 ( );
FILL FILL_11_4_0 ( );
FILL FILL_11_4_1 ( );
FILL FILL_11_5_0 ( );
FILL FILL_11_5_1 ( );
FILL FILL_11_6_0 ( );
FILL FILL_11_6_1 ( );
FILL FILL_11_7_0 ( );
FILL FILL_11_7_1 ( );
FILL FILL_11_8_0 ( );
FILL FILL_11_8_1 ( );
FILL FILL_11_9_0 ( );
FILL FILL_11_9_1 ( );
FILL FILL_11_10_0 ( );
FILL FILL_11_10_1 ( );
FILL FILL_11_11_0 ( );
FILL FILL_11_11_1 ( );
FILL FILL_11_12_0 ( );
FILL FILL_11_12_1 ( );
FILL FILL_11_13_0 ( );
FILL FILL_11_13_1 ( );
FILL FILL_11_14_0 ( );
FILL FILL_11_14_1 ( );
FILL FILL_11_15_0 ( );
FILL FILL_11_15_1 ( );
FILL FILL_11_16_0 ( );
FILL FILL_11_16_1 ( );
FILL FILL_11_17_0 ( );
FILL FILL_11_17_1 ( );
FILL FILL_11_18_0 ( );
FILL FILL_11_18_1 ( );
FILL FILL_12_1 ( );
FILL FILL_12_2 ( );
FILL FILL_12_3 ( );
FILL FILL_12_4 ( );
FILL FILL_12_0_0 ( );
FILL FILL_12_0_1 ( );
FILL FILL_12_1_0 ( );
FILL FILL_12_1_1 ( );
FILL FILL_12_2_0 ( );
FILL FILL_12_2_1 ( );
FILL FILL_12_3_0 ( );
FILL FILL_12_3_1 ( );
FILL FILL_12_4_0 ( );
FILL FILL_12_4_1 ( );
FILL FILL_12_5_0 ( );
FILL FILL_12_5_1 ( );
FILL FILL_12_6_0 ( );
FILL FILL_12_6_1 ( );
FILL FILL_12_7_0 ( );
FILL FILL_12_7_1 ( );
FILL FILL_12_8_0 ( );
FILL FILL_12_8_1 ( );
FILL FILL_12_9_0 ( );
FILL FILL_12_9_1 ( );
FILL FILL_12_10_0 ( );
FILL FILL_12_10_1 ( );
FILL FILL_12_11_0 ( );
FILL FILL_12_11_1 ( );
FILL FILL_12_12_0 ( );
FILL FILL_12_12_1 ( );
FILL FILL_12_13_0 ( );
FILL FILL_12_13_1 ( );
FILL FILL_12_14_0 ( );
FILL FILL_12_14_1 ( );
FILL FILL_12_15_0 ( );
FILL FILL_12_15_1 ( );
FILL FILL_12_16_0 ( );
FILL FILL_12_16_1 ( );
FILL FILL_12_17_0 ( );
FILL FILL_12_17_1 ( );
FILL FILL_12_18_0 ( );
FILL FILL_12_18_1 ( );
FILL FILL_13_0_0 ( );
FILL FILL_13_0_1 ( );
FILL FILL_13_1_0 ( );
FILL FILL_13_1_1 ( );
FILL FILL_13_2_0 ( );
FILL FILL_13_2_1 ( );
FILL FILL_13_3_0 ( );
FILL FILL_13_3_1 ( );
FILL FILL_13_4_0 ( );
FILL FILL_13_4_1 ( );
FILL FILL_13_5_0 ( );
FILL FILL_13_5_1 ( );
FILL FILL_13_6_0 ( );
FILL FILL_13_6_1 ( );
FILL FILL_13_7_0 ( );
FILL FILL_13_7_1 ( );
FILL FILL_13_8_0 ( );
FILL FILL_13_8_1 ( );
FILL FILL_13_9_0 ( );
FILL FILL_13_9_1 ( );
FILL FILL_13_10_0 ( );
FILL FILL_13_10_1 ( );
FILL FILL_13_11_0 ( );
FILL FILL_13_11_1 ( );
FILL FILL_13_12_0 ( );
FILL FILL_13_12_1 ( );
FILL FILL_13_13_0 ( );
FILL FILL_13_13_1 ( );
FILL FILL_13_14_0 ( );
FILL FILL_13_14_1 ( );
FILL FILL_13_15_0 ( );
FILL FILL_13_15_1 ( );
FILL FILL_13_16_0 ( );
FILL FILL_13_16_1 ( );
FILL FILL_13_17_0 ( );
FILL FILL_13_17_1 ( );
FILL FILL_13_18_0 ( );
FILL FILL_13_18_1 ( );
FILL FILL_14_0_0 ( );
FILL FILL_14_0_1 ( );
FILL FILL_14_1_0 ( );
FILL FILL_14_1_1 ( );
FILL FILL_14_2_0 ( );
FILL FILL_14_2_1 ( );
FILL FILL_14_3_0 ( );
FILL FILL_14_3_1 ( );
FILL FILL_14_4_0 ( );
FILL FILL_14_4_1 ( );
FILL FILL_14_5_0 ( );
FILL FILL_14_5_1 ( );
FILL FILL_14_6_0 ( );
FILL FILL_14_6_1 ( );
FILL FILL_14_7_0 ( );
FILL FILL_14_7_1 ( );
FILL FILL_14_8_0 ( );
FILL FILL_14_8_1 ( );
FILL FILL_14_9_0 ( );
FILL FILL_14_9_1 ( );
FILL FILL_14_10_0 ( );
FILL FILL_14_10_1 ( );
FILL FILL_14_11_0 ( );
FILL FILL_14_11_1 ( );
FILL FILL_14_12_0 ( );
FILL FILL_14_12_1 ( );
FILL FILL_14_13_0 ( );
FILL FILL_14_13_1 ( );
FILL FILL_14_14_0 ( );
FILL FILL_14_14_1 ( );
FILL FILL_14_15_0 ( );
FILL FILL_14_15_1 ( );
FILL FILL_14_16_0 ( );
FILL FILL_14_16_1 ( );
FILL FILL_14_17_0 ( );
FILL FILL_14_17_1 ( );
FILL FILL_14_18_0 ( );
FILL FILL_14_18_1 ( );
FILL FILL_15_0_0 ( );
FILL FILL_15_0_1 ( );
FILL FILL_15_1_0 ( );
FILL FILL_15_1_1 ( );
FILL FILL_15_2_0 ( );
FILL FILL_15_2_1 ( );
FILL FILL_15_3_0 ( );
FILL FILL_15_3_1 ( );
FILL FILL_15_4_0 ( );
FILL FILL_15_4_1 ( );
FILL FILL_15_5_0 ( );
FILL FILL_15_5_1 ( );
FILL FILL_15_6_0 ( );
FILL FILL_15_6_1 ( );
FILL FILL_15_7_0 ( );
FILL FILL_15_7_1 ( );
FILL FILL_15_8_0 ( );
FILL FILL_15_8_1 ( );
FILL FILL_15_9_0 ( );
FILL FILL_15_9_1 ( );
FILL FILL_15_10_0 ( );
FILL FILL_15_10_1 ( );
FILL FILL_15_11_0 ( );
FILL FILL_15_11_1 ( );
FILL FILL_15_12_0 ( );
FILL FILL_15_12_1 ( );
FILL FILL_15_13_0 ( );
FILL FILL_15_13_1 ( );
FILL FILL_15_14_0 ( );
FILL FILL_15_14_1 ( );
FILL FILL_15_15_0 ( );
FILL FILL_15_15_1 ( );
FILL FILL_15_16_0 ( );
FILL FILL_15_16_1 ( );
FILL FILL_15_17_0 ( );
FILL FILL_15_17_1 ( );
FILL FILL_15_18_0 ( );
FILL FILL_15_18_1 ( );
FILL FILL_16_1 ( );
FILL FILL_16_2 ( );
FILL FILL_16_3 ( );
FILL FILL_16_0_0 ( );
FILL FILL_16_0_1 ( );
FILL FILL_16_1_0 ( );
FILL FILL_16_1_1 ( );
FILL FILL_16_2_0 ( );
FILL FILL_16_2_1 ( );
FILL FILL_16_3_0 ( );
FILL FILL_16_3_1 ( );
FILL FILL_16_4_0 ( );
FILL FILL_16_4_1 ( );
FILL FILL_16_5_0 ( );
FILL FILL_16_5_1 ( );
FILL FILL_16_6_0 ( );
FILL FILL_16_6_1 ( );
FILL FILL_16_7_0 ( );
FILL FILL_16_7_1 ( );
FILL FILL_16_8_0 ( );
FILL FILL_16_8_1 ( );
FILL FILL_16_9_0 ( );
FILL FILL_16_9_1 ( );
FILL FILL_16_10_0 ( );
FILL FILL_16_10_1 ( );
FILL FILL_16_11_0 ( );
FILL FILL_16_11_1 ( );
FILL FILL_16_12_0 ( );
FILL FILL_16_12_1 ( );
FILL FILL_16_13_0 ( );
FILL FILL_16_13_1 ( );
FILL FILL_16_14_0 ( );
FILL FILL_16_14_1 ( );
FILL FILL_16_15_0 ( );
FILL FILL_16_15_1 ( );
FILL FILL_16_16_0 ( );
FILL FILL_16_16_1 ( );
FILL FILL_16_17_0 ( );
FILL FILL_16_17_1 ( );
FILL FILL_16_18_0 ( );
FILL FILL_16_18_1 ( );
FILL FILL_17_1 ( );
FILL FILL_17_2 ( );
FILL FILL_17_0_0 ( );
FILL FILL_17_0_1 ( );
FILL FILL_17_1_0 ( );
FILL FILL_17_1_1 ( );
FILL FILL_17_2_0 ( );
FILL FILL_17_2_1 ( );
FILL FILL_17_3_0 ( );
FILL FILL_17_3_1 ( );
FILL FILL_17_4_0 ( );
FILL FILL_17_4_1 ( );
FILL FILL_17_5_0 ( );
FILL FILL_17_5_1 ( );
FILL FILL_17_6_0 ( );
FILL FILL_17_6_1 ( );
FILL FILL_17_7_0 ( );
FILL FILL_17_7_1 ( );
FILL FILL_17_8_0 ( );
FILL FILL_17_8_1 ( );
FILL FILL_17_9_0 ( );
FILL FILL_17_9_1 ( );
FILL FILL_17_10_0 ( );
FILL FILL_17_10_1 ( );
FILL FILL_17_11_0 ( );
FILL FILL_17_11_1 ( );
FILL FILL_17_12_0 ( );
FILL FILL_17_12_1 ( );
FILL FILL_17_13_0 ( );
FILL FILL_17_13_1 ( );
FILL FILL_17_14_0 ( );
FILL FILL_17_14_1 ( );
FILL FILL_17_15_0 ( );
FILL FILL_17_15_1 ( );
FILL FILL_17_16_0 ( );
FILL FILL_17_16_1 ( );
FILL FILL_17_17_0 ( );
FILL FILL_17_17_1 ( );
FILL FILL_17_18_0 ( );
FILL FILL_17_18_1 ( );
FILL FILL_18_1 ( );
FILL FILL_18_2 ( );
FILL FILL_18_3 ( );
FILL FILL_18_4 ( );
FILL FILL_18_0_0 ( );
FILL FILL_18_0_1 ( );
FILL FILL_18_1_0 ( );
FILL FILL_18_1_1 ( );
FILL FILL_18_2_0 ( );
FILL FILL_18_2_1 ( );
FILL FILL_18_3_0 ( );
FILL FILL_18_3_1 ( );
FILL FILL_18_4_0 ( );
FILL FILL_18_4_1 ( );
FILL FILL_18_5_0 ( );
FILL FILL_18_5_1 ( );
FILL FILL_18_6_0 ( );
FILL FILL_18_6_1 ( );
FILL FILL_18_7_0 ( );
FILL FILL_18_7_1 ( );
FILL FILL_18_8_0 ( );
FILL FILL_18_8_1 ( );
FILL FILL_18_9_0 ( );
FILL FILL_18_9_1 ( );
FILL FILL_18_10_0 ( );
FILL FILL_18_10_1 ( );
FILL FILL_18_11_0 ( );
FILL FILL_18_11_1 ( );
FILL FILL_18_12_0 ( );
FILL FILL_18_12_1 ( );
FILL FILL_18_13_0 ( );
FILL FILL_18_13_1 ( );
FILL FILL_18_14_0 ( );
FILL FILL_18_14_1 ( );
FILL FILL_18_15_0 ( );
FILL FILL_18_15_1 ( );
FILL FILL_18_16_0 ( );
FILL FILL_18_16_1 ( );
FILL FILL_18_17_0 ( );
FILL FILL_18_17_1 ( );
FILL FILL_18_18_0 ( );
FILL FILL_18_18_1 ( );
FILL FILL_19_1 ( );
FILL FILL_19_2 ( );
FILL FILL_19_3 ( );
FILL FILL_19_4 ( );
FILL FILL_19_0_0 ( );
FILL FILL_19_0_1 ( );
FILL FILL_19_1_0 ( );
FILL FILL_19_1_1 ( );
FILL FILL_19_2_0 ( );
FILL FILL_19_2_1 ( );
FILL FILL_19_3_0 ( );
FILL FILL_19_3_1 ( );
FILL FILL_19_4_0 ( );
FILL FILL_19_4_1 ( );
FILL FILL_19_5_0 ( );
FILL FILL_19_5_1 ( );
FILL FILL_19_6_0 ( );
FILL FILL_19_6_1 ( );
FILL FILL_19_7_0 ( );
FILL FILL_19_7_1 ( );
FILL FILL_19_8_0 ( );
FILL FILL_19_8_1 ( );
FILL FILL_19_9_0 ( );
FILL FILL_19_9_1 ( );
FILL FILL_19_10_0 ( );
FILL FILL_19_10_1 ( );
FILL FILL_19_11_0 ( );
FILL FILL_19_11_1 ( );
FILL FILL_19_12_0 ( );
FILL FILL_19_12_1 ( );
FILL FILL_19_13_0 ( );
FILL FILL_19_13_1 ( );
FILL FILL_19_14_0 ( );
FILL FILL_19_14_1 ( );
FILL FILL_19_15_0 ( );
FILL FILL_19_15_1 ( );
FILL FILL_19_16_0 ( );
FILL FILL_19_16_1 ( );
FILL FILL_19_17_0 ( );
FILL FILL_19_17_1 ( );
FILL FILL_19_18_0 ( );
FILL FILL_19_18_1 ( );
FILL FILL_20_0_0 ( );
FILL FILL_20_0_1 ( );
FILL FILL_20_1_0 ( );
FILL FILL_20_1_1 ( );
FILL FILL_20_2_0 ( );
FILL FILL_20_2_1 ( );
FILL FILL_20_3_0 ( );
FILL FILL_20_3_1 ( );
FILL FILL_20_4_0 ( );
FILL FILL_20_4_1 ( );
FILL FILL_20_5_0 ( );
FILL FILL_20_5_1 ( );
FILL FILL_20_6_0 ( );
FILL FILL_20_6_1 ( );
FILL FILL_20_7_0 ( );
FILL FILL_20_7_1 ( );
FILL FILL_20_8_0 ( );
FILL FILL_20_8_1 ( );
FILL FILL_20_9_0 ( );
FILL FILL_20_9_1 ( );
FILL FILL_20_10_0 ( );
FILL FILL_20_10_1 ( );
FILL FILL_20_11_0 ( );
FILL FILL_20_11_1 ( );
FILL FILL_20_12_0 ( );
FILL FILL_20_12_1 ( );
FILL FILL_20_13_0 ( );
FILL FILL_20_13_1 ( );
FILL FILL_20_14_0 ( );
FILL FILL_20_14_1 ( );
FILL FILL_20_15_0 ( );
FILL FILL_20_15_1 ( );
FILL FILL_20_16_0 ( );
FILL FILL_20_16_1 ( );
FILL FILL_20_17_0 ( );
FILL FILL_20_17_1 ( );
FILL FILL_20_18_0 ( );
FILL FILL_20_18_1 ( );
FILL FILL_21_1 ( );
FILL FILL_21_2 ( );
FILL FILL_21_3 ( );
FILL FILL_21_0_0 ( );
FILL FILL_21_0_1 ( );
FILL FILL_21_1_0 ( );
FILL FILL_21_1_1 ( );
FILL FILL_21_2_0 ( );
FILL FILL_21_2_1 ( );
FILL FILL_21_3_0 ( );
FILL FILL_21_3_1 ( );
FILL FILL_21_4_0 ( );
FILL FILL_21_4_1 ( );
FILL FILL_21_5_0 ( );
FILL FILL_21_5_1 ( );
FILL FILL_21_6_0 ( );
FILL FILL_21_6_1 ( );
FILL FILL_21_7_0 ( );
FILL FILL_21_7_1 ( );
FILL FILL_21_8_0 ( );
FILL FILL_21_8_1 ( );
FILL FILL_21_9_0 ( );
FILL FILL_21_9_1 ( );
FILL FILL_21_10_0 ( );
FILL FILL_21_10_1 ( );
FILL FILL_21_11_0 ( );
FILL FILL_21_11_1 ( );
FILL FILL_21_12_0 ( );
FILL FILL_21_12_1 ( );
FILL FILL_21_13_0 ( );
FILL FILL_21_13_1 ( );
FILL FILL_21_14_0 ( );
FILL FILL_21_14_1 ( );
FILL FILL_21_15_0 ( );
FILL FILL_21_15_1 ( );
FILL FILL_21_16_0 ( );
FILL FILL_21_16_1 ( );
FILL FILL_21_17_0 ( );
FILL FILL_21_17_1 ( );
FILL FILL_21_18_0 ( );
FILL FILL_21_18_1 ( );
FILL FILL_22_1 ( );
FILL FILL_22_2 ( );
FILL FILL_22_3 ( );
FILL FILL_22_0_0 ( );
FILL FILL_22_0_1 ( );
FILL FILL_22_1_0 ( );
FILL FILL_22_1_1 ( );
FILL FILL_22_2_0 ( );
FILL FILL_22_2_1 ( );
FILL FILL_22_3_0 ( );
FILL FILL_22_3_1 ( );
FILL FILL_22_4_0 ( );
FILL FILL_22_4_1 ( );
FILL FILL_22_5_0 ( );
FILL FILL_22_5_1 ( );
FILL FILL_22_6_0 ( );
FILL FILL_22_6_1 ( );
FILL FILL_22_7_0 ( );
FILL FILL_22_7_1 ( );
FILL FILL_22_8_0 ( );
FILL FILL_22_8_1 ( );
FILL FILL_22_9_0 ( );
FILL FILL_22_9_1 ( );
FILL FILL_22_10_0 ( );
FILL FILL_22_10_1 ( );
FILL FILL_22_11_0 ( );
FILL FILL_22_11_1 ( );
FILL FILL_22_12_0 ( );
FILL FILL_22_12_1 ( );
FILL FILL_22_13_0 ( );
FILL FILL_22_13_1 ( );
FILL FILL_22_14_0 ( );
FILL FILL_22_14_1 ( );
FILL FILL_22_15_0 ( );
FILL FILL_22_15_1 ( );
FILL FILL_22_16_0 ( );
FILL FILL_22_16_1 ( );
FILL FILL_22_17_0 ( );
FILL FILL_22_17_1 ( );
FILL FILL_22_18_0 ( );
FILL FILL_22_18_1 ( );
FILL FILL_23_1 ( );
FILL FILL_23_0_0 ( );
FILL FILL_23_0_1 ( );
FILL FILL_23_1_0 ( );
FILL FILL_23_1_1 ( );
FILL FILL_23_2_0 ( );
FILL FILL_23_2_1 ( );
FILL FILL_23_3_0 ( );
FILL FILL_23_3_1 ( );
FILL FILL_23_4_0 ( );
FILL FILL_23_4_1 ( );
FILL FILL_23_5_0 ( );
FILL FILL_23_5_1 ( );
FILL FILL_23_6_0 ( );
FILL FILL_23_6_1 ( );
FILL FILL_23_7_0 ( );
FILL FILL_23_7_1 ( );
FILL FILL_23_8_0 ( );
FILL FILL_23_8_1 ( );
FILL FILL_23_9_0 ( );
FILL FILL_23_9_1 ( );
FILL FILL_23_10_0 ( );
FILL FILL_23_10_1 ( );
FILL FILL_23_11_0 ( );
FILL FILL_23_11_1 ( );
FILL FILL_23_12_0 ( );
FILL FILL_23_12_1 ( );
FILL FILL_23_13_0 ( );
FILL FILL_23_13_1 ( );
FILL FILL_23_14_0 ( );
FILL FILL_23_14_1 ( );
FILL FILL_23_15_0 ( );
FILL FILL_23_15_1 ( );
FILL FILL_23_16_0 ( );
FILL FILL_23_16_1 ( );
FILL FILL_23_17_0 ( );
FILL FILL_23_17_1 ( );
FILL FILL_23_18_0 ( );
FILL FILL_23_18_1 ( );
FILL FILL_24_1 ( );
FILL FILL_24_2 ( );
FILL FILL_24_3 ( );
FILL FILL_24_4 ( );
FILL FILL_24_0_0 ( );
FILL FILL_24_0_1 ( );
FILL FILL_24_1_0 ( );
FILL FILL_24_1_1 ( );
FILL FILL_24_2_0 ( );
FILL FILL_24_2_1 ( );
FILL FILL_24_3_0 ( );
FILL FILL_24_3_1 ( );
FILL FILL_24_4_0 ( );
FILL FILL_24_4_1 ( );
FILL FILL_24_5_0 ( );
FILL FILL_24_5_1 ( );
FILL FILL_24_6_0 ( );
FILL FILL_24_6_1 ( );
FILL FILL_24_7_0 ( );
FILL FILL_24_7_1 ( );
FILL FILL_24_8_0 ( );
FILL FILL_24_8_1 ( );
FILL FILL_24_9_0 ( );
FILL FILL_24_9_1 ( );
FILL FILL_24_10_0 ( );
FILL FILL_24_10_1 ( );
FILL FILL_24_11_0 ( );
FILL FILL_24_11_1 ( );
FILL FILL_24_12_0 ( );
FILL FILL_24_12_1 ( );
FILL FILL_24_13_0 ( );
FILL FILL_24_13_1 ( );
FILL FILL_24_14_0 ( );
FILL FILL_24_14_1 ( );
FILL FILL_24_15_0 ( );
FILL FILL_24_15_1 ( );
FILL FILL_24_16_0 ( );
FILL FILL_24_16_1 ( );
FILL FILL_24_17_0 ( );
FILL FILL_24_17_1 ( );
FILL FILL_24_18_0 ( );
FILL FILL_24_18_1 ( );
FILL FILL_25_1 ( );
FILL FILL_25_2 ( );
FILL FILL_25_0_0 ( );
FILL FILL_25_0_1 ( );
FILL FILL_25_1_0 ( );
FILL FILL_25_1_1 ( );
FILL FILL_25_2_0 ( );
FILL FILL_25_2_1 ( );
FILL FILL_25_3_0 ( );
FILL FILL_25_3_1 ( );
FILL FILL_25_4_0 ( );
FILL FILL_25_4_1 ( );
FILL FILL_25_5_0 ( );
FILL FILL_25_5_1 ( );
FILL FILL_25_6_0 ( );
FILL FILL_25_6_1 ( );
FILL FILL_25_7_0 ( );
FILL FILL_25_7_1 ( );
FILL FILL_25_8_0 ( );
FILL FILL_25_8_1 ( );
FILL FILL_25_9_0 ( );
FILL FILL_25_9_1 ( );
FILL FILL_25_10_0 ( );
FILL FILL_25_10_1 ( );
FILL FILL_25_11_0 ( );
FILL FILL_25_11_1 ( );
FILL FILL_25_12_0 ( );
FILL FILL_25_12_1 ( );
FILL FILL_25_13_0 ( );
FILL FILL_25_13_1 ( );
FILL FILL_25_14_0 ( );
FILL FILL_25_14_1 ( );
FILL FILL_25_15_0 ( );
FILL FILL_25_15_1 ( );
FILL FILL_25_16_0 ( );
FILL FILL_25_16_1 ( );
FILL FILL_25_17_0 ( );
FILL FILL_25_17_1 ( );
FILL FILL_25_18_0 ( );
FILL FILL_25_18_1 ( );
FILL FILL_26_1 ( );
FILL FILL_26_2 ( );
FILL FILL_26_0_0 ( );
FILL FILL_26_0_1 ( );
FILL FILL_26_1_0 ( );
FILL FILL_26_1_1 ( );
FILL FILL_26_2_0 ( );
FILL FILL_26_2_1 ( );
FILL FILL_26_3_0 ( );
FILL FILL_26_3_1 ( );
FILL FILL_26_4_0 ( );
FILL FILL_26_4_1 ( );
FILL FILL_26_5_0 ( );
FILL FILL_26_5_1 ( );
FILL FILL_26_6_0 ( );
FILL FILL_26_6_1 ( );
FILL FILL_26_7_0 ( );
FILL FILL_26_7_1 ( );
FILL FILL_26_8_0 ( );
FILL FILL_26_8_1 ( );
FILL FILL_26_9_0 ( );
FILL FILL_26_9_1 ( );
FILL FILL_26_10_0 ( );
FILL FILL_26_10_1 ( );
FILL FILL_26_11_0 ( );
FILL FILL_26_11_1 ( );
FILL FILL_26_12_0 ( );
FILL FILL_26_12_1 ( );
FILL FILL_26_13_0 ( );
FILL FILL_26_13_1 ( );
FILL FILL_26_14_0 ( );
FILL FILL_26_14_1 ( );
FILL FILL_26_15_0 ( );
FILL FILL_26_15_1 ( );
FILL FILL_26_16_0 ( );
FILL FILL_26_16_1 ( );
FILL FILL_26_17_0 ( );
FILL FILL_26_17_1 ( );
FILL FILL_26_18_0 ( );
FILL FILL_26_18_1 ( );
FILL FILL_27_1 ( );
FILL FILL_27_2 ( );
FILL FILL_27_0_0 ( );
FILL FILL_27_0_1 ( );
FILL FILL_27_1_0 ( );
FILL FILL_27_1_1 ( );
FILL FILL_27_2_0 ( );
FILL FILL_27_2_1 ( );
FILL FILL_27_3_0 ( );
FILL FILL_27_3_1 ( );
FILL FILL_27_4_0 ( );
FILL FILL_27_4_1 ( );
FILL FILL_27_5_0 ( );
FILL FILL_27_5_1 ( );
FILL FILL_27_6_0 ( );
FILL FILL_27_6_1 ( );
FILL FILL_27_7_0 ( );
FILL FILL_27_7_1 ( );
FILL FILL_27_8_0 ( );
FILL FILL_27_8_1 ( );
FILL FILL_27_9_0 ( );
FILL FILL_27_9_1 ( );
FILL FILL_27_10_0 ( );
FILL FILL_27_10_1 ( );
FILL FILL_27_11_0 ( );
FILL FILL_27_11_1 ( );
FILL FILL_27_12_0 ( );
FILL FILL_27_12_1 ( );
FILL FILL_27_13_0 ( );
FILL FILL_27_13_1 ( );
FILL FILL_27_14_0 ( );
FILL FILL_27_14_1 ( );
FILL FILL_27_15_0 ( );
FILL FILL_27_15_1 ( );
FILL FILL_27_16_0 ( );
FILL FILL_27_16_1 ( );
FILL FILL_27_17_0 ( );
FILL FILL_27_17_1 ( );
FILL FILL_27_18_0 ( );
FILL FILL_27_18_1 ( );
FILL FILL_28_1 ( );
FILL FILL_28_0_0 ( );
FILL FILL_28_0_1 ( );
FILL FILL_28_1_0 ( );
FILL FILL_28_1_1 ( );
FILL FILL_28_2_0 ( );
FILL FILL_28_2_1 ( );
FILL FILL_28_3_0 ( );
FILL FILL_28_3_1 ( );
FILL FILL_28_4_0 ( );
FILL FILL_28_4_1 ( );
FILL FILL_28_5_0 ( );
FILL FILL_28_5_1 ( );
FILL FILL_28_6_0 ( );
FILL FILL_28_6_1 ( );
FILL FILL_28_7_0 ( );
FILL FILL_28_7_1 ( );
FILL FILL_28_8_0 ( );
FILL FILL_28_8_1 ( );
FILL FILL_28_9_0 ( );
FILL FILL_28_9_1 ( );
FILL FILL_28_10_0 ( );
FILL FILL_28_10_1 ( );
FILL FILL_28_11_0 ( );
FILL FILL_28_11_1 ( );
FILL FILL_28_12_0 ( );
FILL FILL_28_12_1 ( );
FILL FILL_28_13_0 ( );
FILL FILL_28_13_1 ( );
FILL FILL_28_14_0 ( );
FILL FILL_28_14_1 ( );
FILL FILL_28_15_0 ( );
FILL FILL_28_15_1 ( );
FILL FILL_28_16_0 ( );
FILL FILL_28_16_1 ( );
FILL FILL_28_17_0 ( );
FILL FILL_28_17_1 ( );
FILL FILL_28_18_0 ( );
FILL FILL_28_18_1 ( );
FILL FILL_29_1 ( );
FILL FILL_29_2 ( );
FILL FILL_29_3 ( );
FILL FILL_29_4 ( );
FILL FILL_29_0_0 ( );
FILL FILL_29_0_1 ( );
FILL FILL_29_1_0 ( );
FILL FILL_29_1_1 ( );
FILL FILL_29_2_0 ( );
FILL FILL_29_2_1 ( );
FILL FILL_29_3_0 ( );
FILL FILL_29_3_1 ( );
FILL FILL_29_4_0 ( );
FILL FILL_29_4_1 ( );
FILL FILL_29_5_0 ( );
FILL FILL_29_5_1 ( );
FILL FILL_29_6_0 ( );
FILL FILL_29_6_1 ( );
FILL FILL_29_7_0 ( );
FILL FILL_29_7_1 ( );
FILL FILL_29_8_0 ( );
FILL FILL_29_8_1 ( );
FILL FILL_29_9_0 ( );
FILL FILL_29_9_1 ( );
FILL FILL_29_10_0 ( );
FILL FILL_29_10_1 ( );
FILL FILL_29_11_0 ( );
FILL FILL_29_11_1 ( );
FILL FILL_29_12_0 ( );
FILL FILL_29_12_1 ( );
FILL FILL_29_13_0 ( );
FILL FILL_29_13_1 ( );
FILL FILL_29_14_0 ( );
FILL FILL_29_14_1 ( );
FILL FILL_29_15_0 ( );
FILL FILL_29_15_1 ( );
FILL FILL_29_16_0 ( );
FILL FILL_29_16_1 ( );
FILL FILL_29_17_0 ( );
FILL FILL_29_17_1 ( );
FILL FILL_29_18_0 ( );
FILL FILL_29_18_1 ( );
FILL FILL_30_1 ( );
FILL FILL_30_0_0 ( );
FILL FILL_30_0_1 ( );
FILL FILL_30_1_0 ( );
FILL FILL_30_1_1 ( );
FILL FILL_30_2_0 ( );
FILL FILL_30_2_1 ( );
FILL FILL_30_3_0 ( );
FILL FILL_30_3_1 ( );
FILL FILL_30_4_0 ( );
FILL FILL_30_4_1 ( );
FILL FILL_30_5_0 ( );
FILL FILL_30_5_1 ( );
FILL FILL_30_6_0 ( );
FILL FILL_30_6_1 ( );
FILL FILL_30_7_0 ( );
FILL FILL_30_7_1 ( );
FILL FILL_30_8_0 ( );
FILL FILL_30_8_1 ( );
FILL FILL_30_9_0 ( );
FILL FILL_30_9_1 ( );
FILL FILL_30_10_0 ( );
FILL FILL_30_10_1 ( );
FILL FILL_30_11_0 ( );
FILL FILL_30_11_1 ( );
FILL FILL_30_12_0 ( );
FILL FILL_30_12_1 ( );
FILL FILL_30_13_0 ( );
FILL FILL_30_13_1 ( );
FILL FILL_30_14_0 ( );
FILL FILL_30_14_1 ( );
FILL FILL_30_15_0 ( );
FILL FILL_30_15_1 ( );
FILL FILL_30_16_0 ( );
FILL FILL_30_16_1 ( );
FILL FILL_30_17_0 ( );
FILL FILL_30_17_1 ( );
FILL FILL_30_18_0 ( );
FILL FILL_30_18_1 ( );
FILL FILL_31_1 ( );
FILL FILL_31_2 ( );
FILL FILL_31_0_0 ( );
FILL FILL_31_0_1 ( );
FILL FILL_31_1_0 ( );
FILL FILL_31_1_1 ( );
FILL FILL_31_2_0 ( );
FILL FILL_31_2_1 ( );
FILL FILL_31_3_0 ( );
FILL FILL_31_3_1 ( );
FILL FILL_31_4_0 ( );
FILL FILL_31_4_1 ( );
FILL FILL_31_5_0 ( );
FILL FILL_31_5_1 ( );
FILL FILL_31_6_0 ( );
FILL FILL_31_6_1 ( );
FILL FILL_31_7_0 ( );
FILL FILL_31_7_1 ( );
FILL FILL_31_8_0 ( );
FILL FILL_31_8_1 ( );
FILL FILL_31_9_0 ( );
FILL FILL_31_9_1 ( );
FILL FILL_31_10_0 ( );
FILL FILL_31_10_1 ( );
FILL FILL_31_11_0 ( );
FILL FILL_31_11_1 ( );
FILL FILL_31_12_0 ( );
FILL FILL_31_12_1 ( );
FILL FILL_31_13_0 ( );
FILL FILL_31_13_1 ( );
FILL FILL_31_14_0 ( );
FILL FILL_31_14_1 ( );
FILL FILL_31_15_0 ( );
FILL FILL_31_15_1 ( );
FILL FILL_31_16_0 ( );
FILL FILL_31_16_1 ( );
FILL FILL_31_17_0 ( );
FILL FILL_31_17_1 ( );
FILL FILL_31_18_0 ( );
FILL FILL_31_18_1 ( );
FILL FILL_32_1 ( );
FILL FILL_32_0_0 ( );
FILL FILL_32_0_1 ( );
FILL FILL_32_1_0 ( );
FILL FILL_32_1_1 ( );
FILL FILL_32_2_0 ( );
FILL FILL_32_2_1 ( );
FILL FILL_32_3_0 ( );
FILL FILL_32_3_1 ( );
FILL FILL_32_4_0 ( );
FILL FILL_32_4_1 ( );
FILL FILL_32_5_0 ( );
FILL FILL_32_5_1 ( );
FILL FILL_32_6_0 ( );
FILL FILL_32_6_1 ( );
FILL FILL_32_7_0 ( );
FILL FILL_32_7_1 ( );
FILL FILL_32_8_0 ( );
FILL FILL_32_8_1 ( );
FILL FILL_32_9_0 ( );
FILL FILL_32_9_1 ( );
FILL FILL_32_10_0 ( );
FILL FILL_32_10_1 ( );
FILL FILL_32_11_0 ( );
FILL FILL_32_11_1 ( );
FILL FILL_32_12_0 ( );
FILL FILL_32_12_1 ( );
FILL FILL_32_13_0 ( );
FILL FILL_32_13_1 ( );
FILL FILL_32_14_0 ( );
FILL FILL_32_14_1 ( );
FILL FILL_32_15_0 ( );
FILL FILL_32_15_1 ( );
FILL FILL_32_16_0 ( );
FILL FILL_32_16_1 ( );
FILL FILL_32_17_0 ( );
FILL FILL_32_17_1 ( );
FILL FILL_32_18_0 ( );
FILL FILL_32_18_1 ( );
FILL FILL_33_1 ( );
FILL FILL_33_0_0 ( );
FILL FILL_33_0_1 ( );
FILL FILL_33_1_0 ( );
FILL FILL_33_1_1 ( );
FILL FILL_33_2_0 ( );
FILL FILL_33_2_1 ( );
FILL FILL_33_3_0 ( );
FILL FILL_33_3_1 ( );
FILL FILL_33_4_0 ( );
FILL FILL_33_4_1 ( );
FILL FILL_33_5_0 ( );
FILL FILL_33_5_1 ( );
FILL FILL_33_6_0 ( );
FILL FILL_33_6_1 ( );
FILL FILL_33_7_0 ( );
FILL FILL_33_7_1 ( );
FILL FILL_33_8_0 ( );
FILL FILL_33_8_1 ( );
FILL FILL_33_9_0 ( );
FILL FILL_33_9_1 ( );
FILL FILL_33_10_0 ( );
FILL FILL_33_10_1 ( );
FILL FILL_33_11_0 ( );
FILL FILL_33_11_1 ( );
FILL FILL_33_12_0 ( );
FILL FILL_33_12_1 ( );
FILL FILL_33_13_0 ( );
FILL FILL_33_13_1 ( );
FILL FILL_33_14_0 ( );
FILL FILL_33_14_1 ( );
FILL FILL_33_15_0 ( );
FILL FILL_33_15_1 ( );
FILL FILL_33_16_0 ( );
FILL FILL_33_16_1 ( );
FILL FILL_33_17_0 ( );
FILL FILL_33_17_1 ( );
FILL FILL_33_18_0 ( );
FILL FILL_33_18_1 ( );
FILL FILL_34_1 ( );
FILL FILL_34_2 ( );
FILL FILL_34_3 ( );
FILL FILL_34_4 ( );
FILL FILL_34_0_0 ( );
FILL FILL_34_0_1 ( );
FILL FILL_34_1_0 ( );
FILL FILL_34_1_1 ( );
FILL FILL_34_2_0 ( );
FILL FILL_34_2_1 ( );
FILL FILL_34_3_0 ( );
FILL FILL_34_3_1 ( );
FILL FILL_34_4_0 ( );
FILL FILL_34_4_1 ( );
FILL FILL_34_5_0 ( );
FILL FILL_34_5_1 ( );
FILL FILL_34_6_0 ( );
FILL FILL_34_6_1 ( );
FILL FILL_34_7_0 ( );
FILL FILL_34_7_1 ( );
FILL FILL_34_8_0 ( );
FILL FILL_34_8_1 ( );
FILL FILL_34_9_0 ( );
FILL FILL_34_9_1 ( );
FILL FILL_34_10_0 ( );
FILL FILL_34_10_1 ( );
FILL FILL_34_11_0 ( );
FILL FILL_34_11_1 ( );
FILL FILL_34_12_0 ( );
FILL FILL_34_12_1 ( );
FILL FILL_34_13_0 ( );
FILL FILL_34_13_1 ( );
FILL FILL_34_14_0 ( );
FILL FILL_34_14_1 ( );
FILL FILL_34_15_0 ( );
FILL FILL_34_15_1 ( );
FILL FILL_34_16_0 ( );
FILL FILL_34_16_1 ( );
FILL FILL_34_17_0 ( );
FILL FILL_34_17_1 ( );
FILL FILL_34_18_0 ( );
FILL FILL_34_18_1 ( );
FILL FILL_35_1 ( );
FILL FILL_35_2 ( );
FILL FILL_35_0_0 ( );
FILL FILL_35_0_1 ( );
FILL FILL_35_1_0 ( );
FILL FILL_35_1_1 ( );
FILL FILL_35_2_0 ( );
FILL FILL_35_2_1 ( );
FILL FILL_35_3_0 ( );
FILL FILL_35_3_1 ( );
FILL FILL_35_4_0 ( );
FILL FILL_35_4_1 ( );
FILL FILL_35_5_0 ( );
FILL FILL_35_5_1 ( );
FILL FILL_35_6_0 ( );
FILL FILL_35_6_1 ( );
FILL FILL_35_7_0 ( );
FILL FILL_35_7_1 ( );
FILL FILL_35_8_0 ( );
FILL FILL_35_8_1 ( );
FILL FILL_35_9_0 ( );
FILL FILL_35_9_1 ( );
FILL FILL_35_10_0 ( );
FILL FILL_35_10_1 ( );
FILL FILL_35_11_0 ( );
FILL FILL_35_11_1 ( );
FILL FILL_35_12_0 ( );
FILL FILL_35_12_1 ( );
FILL FILL_35_13_0 ( );
FILL FILL_35_13_1 ( );
FILL FILL_35_14_0 ( );
FILL FILL_35_14_1 ( );
FILL FILL_35_15_0 ( );
FILL FILL_35_15_1 ( );
FILL FILL_35_16_0 ( );
FILL FILL_35_16_1 ( );
FILL FILL_35_17_0 ( );
FILL FILL_35_17_1 ( );
FILL FILL_35_18_0 ( );
FILL FILL_35_18_1 ( );
FILL FILL_36_1 ( );
FILL FILL_36_2 ( );
FILL FILL_36_3 ( );
FILL FILL_36_4 ( );
FILL FILL_36_0_0 ( );
FILL FILL_36_0_1 ( );
FILL FILL_36_1_0 ( );
FILL FILL_36_1_1 ( );
FILL FILL_36_2_0 ( );
FILL FILL_36_2_1 ( );
FILL FILL_36_3_0 ( );
FILL FILL_36_3_1 ( );
FILL FILL_36_4_0 ( );
FILL FILL_36_4_1 ( );
FILL FILL_36_5_0 ( );
FILL FILL_36_5_1 ( );
FILL FILL_36_6_0 ( );
FILL FILL_36_6_1 ( );
FILL FILL_36_7_0 ( );
FILL FILL_36_7_1 ( );
FILL FILL_36_8_0 ( );
FILL FILL_36_8_1 ( );
FILL FILL_36_9_0 ( );
FILL FILL_36_9_1 ( );
FILL FILL_36_10_0 ( );
FILL FILL_36_10_1 ( );
FILL FILL_36_11_0 ( );
FILL FILL_36_11_1 ( );
FILL FILL_36_12_0 ( );
FILL FILL_36_12_1 ( );
FILL FILL_36_13_0 ( );
FILL FILL_36_13_1 ( );
FILL FILL_36_14_0 ( );
FILL FILL_36_14_1 ( );
FILL FILL_36_15_0 ( );
FILL FILL_36_15_1 ( );
FILL FILL_36_16_0 ( );
FILL FILL_36_16_1 ( );
FILL FILL_36_17_0 ( );
FILL FILL_36_17_1 ( );
FILL FILL_36_18_0 ( );
FILL FILL_36_18_1 ( );
FILL FILL_37_1 ( );
FILL FILL_37_0_0 ( );
FILL FILL_37_0_1 ( );
FILL FILL_37_1_0 ( );
FILL FILL_37_1_1 ( );
FILL FILL_37_2_0 ( );
FILL FILL_37_2_1 ( );
FILL FILL_37_3_0 ( );
FILL FILL_37_3_1 ( );
FILL FILL_37_4_0 ( );
FILL FILL_37_4_1 ( );
FILL FILL_37_5_0 ( );
FILL FILL_37_5_1 ( );
FILL FILL_37_6_0 ( );
FILL FILL_37_6_1 ( );
FILL FILL_37_7_0 ( );
FILL FILL_37_7_1 ( );
FILL FILL_37_8_0 ( );
FILL FILL_37_8_1 ( );
FILL FILL_37_9_0 ( );
FILL FILL_37_9_1 ( );
FILL FILL_37_10_0 ( );
FILL FILL_37_10_1 ( );
FILL FILL_37_11_0 ( );
FILL FILL_37_11_1 ( );
FILL FILL_37_12_0 ( );
FILL FILL_37_12_1 ( );
FILL FILL_37_13_0 ( );
FILL FILL_37_13_1 ( );
FILL FILL_37_14_0 ( );
FILL FILL_37_14_1 ( );
FILL FILL_37_15_0 ( );
FILL FILL_37_15_1 ( );
FILL FILL_37_16_0 ( );
FILL FILL_37_16_1 ( );
FILL FILL_37_17_0 ( );
FILL FILL_37_17_1 ( );
FILL FILL_37_18_0 ( );
FILL FILL_37_18_1 ( );
FILL FILL_38_1 ( );
FILL FILL_38_0_0 ( );
FILL FILL_38_0_1 ( );
FILL FILL_38_1_0 ( );
FILL FILL_38_1_1 ( );
FILL FILL_38_2_0 ( );
FILL FILL_38_2_1 ( );
FILL FILL_38_3_0 ( );
FILL FILL_38_3_1 ( );
FILL FILL_38_4_0 ( );
FILL FILL_38_4_1 ( );
FILL FILL_38_5_0 ( );
FILL FILL_38_5_1 ( );
FILL FILL_38_6_0 ( );
FILL FILL_38_6_1 ( );
FILL FILL_38_7_0 ( );
FILL FILL_38_7_1 ( );
FILL FILL_38_8_0 ( );
FILL FILL_38_8_1 ( );
FILL FILL_38_9_0 ( );
FILL FILL_38_9_1 ( );
FILL FILL_38_10_0 ( );
FILL FILL_38_10_1 ( );
FILL FILL_38_11_0 ( );
FILL FILL_38_11_1 ( );
FILL FILL_38_12_0 ( );
FILL FILL_38_12_1 ( );
FILL FILL_38_13_0 ( );
FILL FILL_38_13_1 ( );
FILL FILL_38_14_0 ( );
FILL FILL_38_14_1 ( );
FILL FILL_38_15_0 ( );
FILL FILL_38_15_1 ( );
FILL FILL_38_16_0 ( );
FILL FILL_38_16_1 ( );
FILL FILL_38_17_0 ( );
FILL FILL_38_17_1 ( );
FILL FILL_38_18_0 ( );
FILL FILL_38_18_1 ( );
FILL FILL_39_1 ( );
FILL FILL_39_2 ( );
FILL FILL_39_3 ( );
endmodule
